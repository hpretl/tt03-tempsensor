magic
tech sky130A
magscale 1 2
timestamp 1703666357
<< viali >>
rect 4721 32385 4755 32419
rect 4813 32385 4847 32419
rect 8585 32385 8619 32419
rect 3893 32317 3927 32351
rect 4261 32317 4295 32351
rect 4353 32317 4387 32351
rect 5181 32317 5215 32351
rect 6377 32317 6411 32351
rect 6745 32317 6779 32351
rect 6837 32317 6871 32351
rect 7205 32317 7239 32351
rect 7757 32317 7791 32351
rect 8125 32317 8159 32351
rect 8217 32317 8251 32351
rect 9321 32317 9355 32351
rect 9689 32317 9723 32351
rect 4261 32181 4295 32215
rect 4353 32181 4387 32215
rect 5181 32181 5215 32215
rect 6377 32181 6411 32215
rect 7205 32181 7239 32215
rect 7757 32181 7791 32215
rect 8217 32181 8251 32215
rect 9321 32181 9355 32215
rect 11069 32181 11103 32215
rect 4261 31909 4295 31943
rect 4721 31909 4755 31943
rect 4353 31841 4387 31875
rect 5549 31841 5583 31875
rect 6009 31841 6043 31875
rect 6469 31841 6503 31875
rect 7849 31841 7883 31875
rect 8769 31841 8803 31875
rect 9781 31841 9815 31875
rect 10241 31841 10275 31875
rect 11161 31841 11195 31875
rect 3893 31773 3927 31807
rect 5089 31773 5123 31807
rect 5457 31773 5491 31807
rect 5917 31773 5951 31807
rect 6377 31773 6411 31807
rect 6837 31773 6871 31807
rect 6929 31773 6963 31807
rect 7297 31773 7331 31807
rect 7389 31773 7423 31807
rect 7757 31773 7791 31807
rect 8217 31773 8251 31807
rect 8401 31773 8435 31807
rect 8953 31773 8987 31807
rect 9321 31773 9355 31807
rect 9689 31773 9723 31807
rect 10149 31773 10183 31807
rect 10609 31773 10643 31807
rect 10793 31773 10827 31807
rect 4261 31637 4295 31671
rect 4721 31637 4755 31671
rect 5457 31637 5491 31671
rect 5917 31637 5951 31671
rect 6377 31637 6411 31671
rect 6837 31637 6871 31671
rect 6929 31637 6963 31671
rect 7757 31637 7791 31671
rect 8217 31637 8251 31671
rect 8401 31637 8435 31671
rect 9137 31637 9171 31671
rect 9689 31637 9723 31671
rect 10149 31637 10183 31671
rect 10609 31637 10643 31671
rect 10793 31637 10827 31671
rect 1961 31433 1995 31467
rect 2421 31433 2455 31467
rect 3249 31433 3283 31467
rect 4261 31433 4295 31467
rect 5181 31433 5215 31467
rect 6193 31433 6227 31467
rect 6745 31433 6779 31467
rect 7573 31433 7607 31467
rect 8033 31433 8067 31467
rect 8493 31433 8527 31467
rect 1961 31297 1995 31331
rect 2329 31297 2363 31331
rect 2789 31297 2823 31331
rect 2881 31297 2915 31331
rect 3893 31297 3927 31331
rect 4261 31297 4295 31331
rect 4445 31297 4479 31331
rect 4537 31297 4571 31331
rect 5181 31297 5215 31331
rect 6193 31297 6227 31331
rect 6745 31297 6779 31331
rect 7205 31297 7239 31331
rect 7665 31297 7699 31331
rect 8125 31297 8159 31331
rect 9689 31297 9723 31331
rect 10333 31297 10367 31331
rect 11069 31297 11103 31331
rect 2421 31229 2455 31263
rect 4721 31229 4755 31263
rect 4813 31229 4847 31263
rect 5825 31229 5859 31263
rect 6377 31229 6411 31263
rect 7573 31229 7607 31263
rect 8033 31229 8067 31263
rect 8493 31229 8527 31263
rect 9321 31229 9355 31263
rect 9781 31229 9815 31263
rect 10149 31229 10183 31263
rect 3249 31161 3283 31195
rect 9689 31093 9723 31127
rect 10149 31093 10183 31127
rect 10425 31093 10459 31127
rect 10885 31093 10919 31127
rect 1961 30889 1995 30923
rect 4169 30889 4203 30923
rect 4997 30889 5031 30923
rect 9229 30889 9263 30923
rect 4353 30821 4387 30855
rect 10057 30821 10091 30855
rect 11989 30821 12023 30855
rect 2421 30753 2455 30787
rect 4721 30753 4755 30787
rect 8493 30753 8527 30787
rect 9597 30753 9631 30787
rect 11161 30753 11195 30787
rect 1685 30685 1719 30719
rect 1869 30685 1903 30719
rect 2145 30685 2179 30719
rect 2789 30685 2823 30719
rect 4077 30685 4111 30719
rect 4813 30685 4847 30719
rect 6837 30685 6871 30719
rect 8677 30685 8711 30719
rect 8953 30685 8987 30719
rect 9137 30685 9171 30719
rect 9229 30685 9263 30719
rect 9689 30685 9723 30719
rect 10241 30685 10275 30719
rect 10609 30685 10643 30719
rect 10701 30685 10735 30719
rect 11069 30685 11103 30719
rect 11529 30685 11563 30719
rect 11621 30685 11655 30719
rect 9045 30617 9079 30651
rect 1777 30549 1811 30583
rect 2789 30549 2823 30583
rect 4353 30549 4387 30583
rect 7021 30549 7055 30583
rect 10057 30549 10091 30583
rect 10609 30549 10643 30583
rect 10701 30549 10735 30583
rect 11161 30549 11195 30583
rect 11989 30549 12023 30583
rect 3617 30345 3651 30379
rect 4445 30345 4479 30379
rect 9505 30345 9539 30379
rect 9965 30345 9999 30379
rect 10425 30345 10459 30379
rect 10885 30345 10919 30379
rect 11345 30345 11379 30379
rect 11989 30345 12023 30379
rect 12081 30345 12115 30379
rect 12541 30345 12575 30379
rect 2697 30277 2731 30311
rect 4077 30277 4111 30311
rect 6837 30277 6871 30311
rect 2789 30209 2823 30243
rect 7021 30209 7055 30243
rect 9505 30209 9539 30243
rect 9965 30209 9999 30243
rect 10425 30209 10459 30243
rect 10885 30209 10919 30243
rect 11345 30209 11379 30243
rect 11989 30209 12023 30243
rect 12541 30209 12575 30243
rect 15853 30209 15887 30243
rect 1961 30141 1995 30175
rect 2237 30141 2271 30175
rect 2881 30141 2915 30175
rect 3249 30141 3283 30175
rect 3801 30141 3835 30175
rect 3985 30141 4019 30175
rect 4537 30141 4571 30175
rect 9137 30141 9171 30175
rect 9597 30141 9631 30175
rect 10057 30141 10091 30175
rect 10517 30141 10551 30175
rect 10977 30141 11011 30175
rect 11621 30141 11655 30175
rect 12081 30141 12115 30175
rect 12449 30141 12483 30175
rect 12909 30141 12943 30175
rect 2329 30073 2363 30107
rect 3617 30073 3651 30107
rect 6653 30005 6687 30039
rect 15669 30005 15703 30039
rect 3433 29801 3467 29835
rect 10149 29801 10183 29835
rect 16129 29801 16163 29835
rect 10609 29733 10643 29767
rect 11069 29733 11103 29767
rect 11897 29733 11931 29767
rect 14289 29733 14323 29767
rect 16221 29733 16255 29767
rect 16865 29733 16899 29767
rect 1409 29665 1443 29699
rect 1869 29665 1903 29699
rect 2329 29665 2363 29699
rect 10977 29665 11011 29699
rect 11437 29665 11471 29699
rect 11529 29665 11563 29699
rect 1777 29597 1811 29631
rect 2237 29597 2271 29631
rect 2697 29597 2731 29631
rect 3525 29597 3559 29631
rect 4445 29597 4479 29631
rect 5917 29597 5951 29631
rect 7389 29597 7423 29631
rect 9505 29597 9539 29631
rect 9781 29597 9815 29631
rect 10057 29597 10091 29631
rect 14657 29597 14691 29631
rect 18245 29597 18279 29631
rect 4712 29529 4746 29563
rect 6184 29529 6218 29563
rect 7656 29529 7690 29563
rect 8953 29529 8987 29563
rect 9965 29529 9999 29563
rect 14565 29529 14599 29563
rect 14902 29529 14936 29563
rect 16589 29529 16623 29563
rect 17978 29529 18012 29563
rect 1777 29461 1811 29495
rect 2237 29461 2271 29495
rect 2697 29461 2731 29495
rect 5825 29461 5859 29495
rect 7297 29461 7331 29495
rect 8769 29461 8803 29495
rect 10609 29461 10643 29495
rect 11069 29461 11103 29495
rect 11897 29461 11931 29495
rect 14105 29461 14139 29495
rect 16037 29461 16071 29495
rect 1869 29257 1903 29291
rect 3249 29257 3283 29291
rect 5089 29257 5123 29291
rect 6101 29257 6135 29291
rect 8049 29257 8083 29291
rect 11161 29257 11195 29291
rect 20821 29257 20855 29291
rect 4261 29189 4295 29223
rect 7849 29189 7883 29223
rect 15200 29189 15234 29223
rect 17693 29189 17727 29223
rect 2237 29121 2271 29155
rect 4169 29121 4203 29155
rect 5181 29121 5215 29155
rect 5365 29121 5399 29155
rect 5641 29121 5675 29155
rect 5825 29121 5859 29155
rect 5917 29121 5951 29155
rect 10158 29121 10192 29155
rect 10425 29121 10459 29155
rect 11345 29121 11379 29155
rect 13277 29121 13311 29155
rect 13544 29121 13578 29155
rect 14933 29121 14967 29155
rect 18052 29121 18086 29155
rect 19708 29121 19742 29155
rect 2881 29053 2915 29087
rect 4077 29053 4111 29087
rect 5457 29053 5491 29087
rect 6929 29053 6963 29087
rect 7205 29053 7239 29087
rect 8401 29053 8435 29087
rect 16681 29053 16715 29087
rect 17785 29053 17819 29087
rect 19441 29053 19475 29087
rect 1869 28985 1903 29019
rect 3249 28985 3283 29019
rect 4629 28985 4663 29019
rect 4905 28985 4939 29019
rect 9045 28985 9079 29019
rect 16313 28985 16347 29019
rect 16957 28985 16991 29019
rect 17417 28985 17451 29019
rect 19165 28985 19199 29019
rect 6377 28917 6411 28951
rect 7757 28917 7791 28951
rect 8033 28917 8067 28951
rect 8217 28917 8251 28951
rect 8953 28917 8987 28951
rect 14657 28917 14691 28951
rect 17141 28917 17175 28951
rect 17233 28917 17267 28951
rect 1593 28713 1627 28747
rect 2329 28713 2363 28747
rect 5273 28713 5307 28747
rect 6377 28713 6411 28747
rect 7757 28713 7791 28747
rect 9137 28713 9171 28747
rect 13645 28713 13679 28747
rect 14933 28713 14967 28747
rect 17601 28713 17635 28747
rect 7389 28645 7423 28679
rect 9505 28645 9539 28679
rect 14565 28645 14599 28679
rect 17233 28645 17267 28679
rect 3249 28577 3283 28611
rect 8677 28577 8711 28611
rect 9413 28577 9447 28611
rect 14197 28577 14231 28611
rect 14657 28577 14691 28611
rect 1777 28509 1811 28543
rect 2053 28509 2087 28543
rect 2237 28509 2271 28543
rect 2513 28509 2547 28543
rect 3433 28509 3467 28543
rect 5273 28509 5307 28543
rect 5457 28509 5491 28543
rect 5641 28509 5675 28543
rect 6561 28509 6595 28543
rect 6837 28509 6871 28543
rect 7113 28509 7147 28543
rect 7481 28509 7515 28543
rect 7757 28509 7791 28543
rect 7941 28509 7975 28543
rect 8585 28509 8619 28543
rect 8769 28509 8803 28543
rect 8953 28509 8987 28543
rect 9137 28509 9171 28543
rect 9689 28509 9723 28543
rect 9781 28509 9815 28543
rect 10333 28509 10367 28543
rect 10609 28509 10643 28543
rect 13829 28509 13863 28543
rect 14749 28509 14783 28543
rect 15393 28509 15427 28543
rect 17049 28509 17083 28543
rect 17417 28509 17451 28543
rect 17877 28509 17911 28543
rect 19257 28509 19291 28543
rect 21465 28509 21499 28543
rect 7389 28441 7423 28475
rect 19502 28441 19536 28475
rect 2145 28373 2179 28407
rect 2605 28373 2639 28407
rect 2973 28373 3007 28407
rect 3065 28373 3099 28407
rect 3525 28373 3559 28407
rect 6285 28373 6319 28407
rect 6745 28373 6779 28407
rect 7205 28373 7239 28407
rect 11713 28373 11747 28407
rect 15209 28373 15243 28407
rect 18061 28373 18095 28407
rect 20637 28373 20671 28407
rect 21649 28373 21683 28407
rect 1767 28169 1801 28203
rect 5733 28169 5767 28203
rect 7389 28169 7423 28203
rect 10057 28169 10091 28203
rect 19165 28169 19199 28203
rect 19717 28169 19751 28203
rect 2237 28101 2271 28135
rect 5917 28101 5951 28135
rect 9137 28101 9171 28135
rect 9597 28101 9631 28135
rect 14924 28101 14958 28135
rect 18622 28101 18656 28135
rect 20536 28101 20570 28135
rect 22078 28101 22112 28135
rect 9367 28067 9401 28101
rect 2053 28033 2087 28067
rect 2881 28033 2915 28067
rect 3249 28033 3283 28067
rect 3490 28033 3524 28067
rect 4169 28033 4203 28067
rect 4436 28033 4470 28067
rect 5641 28033 5675 28067
rect 6745 28033 6779 28067
rect 6837 28033 6871 28067
rect 7021 28033 7055 28067
rect 7297 28033 7331 28067
rect 7481 28033 7515 28067
rect 8953 28033 8987 28067
rect 9873 28033 9907 28067
rect 9965 28033 9999 28067
rect 12817 28033 12851 28067
rect 14105 28033 14139 28067
rect 14289 28033 14323 28067
rect 18981 28033 19015 28067
rect 19901 28033 19935 28067
rect 2329 27965 2363 27999
rect 14657 27965 14691 27999
rect 18889 27965 18923 27999
rect 20269 27965 20303 27999
rect 21833 27965 21867 27999
rect 8769 27897 8803 27931
rect 3249 27829 3283 27863
rect 3387 27829 3421 27863
rect 5549 27829 5583 27863
rect 5917 27829 5951 27863
rect 7205 27829 7239 27863
rect 9229 27829 9263 27863
rect 9413 27829 9447 27863
rect 12633 27829 12667 27863
rect 13921 27829 13955 27863
rect 16037 27829 16071 27863
rect 17509 27829 17543 27863
rect 21649 27829 21683 27863
rect 23213 27829 23247 27863
rect 18153 27625 18187 27659
rect 18889 27625 18923 27659
rect 19993 27625 20027 27659
rect 20729 27625 20763 27659
rect 21465 27625 21499 27659
rect 2881 27557 2915 27591
rect 4905 27557 4939 27591
rect 9137 27557 9171 27591
rect 14657 27557 14691 27591
rect 17509 27557 17543 27591
rect 18061 27557 18095 27591
rect 22017 27557 22051 27591
rect 1777 27489 1811 27523
rect 2329 27489 2363 27523
rect 3341 27489 3375 27523
rect 4445 27489 4479 27523
rect 4629 27489 4663 27523
rect 10425 27489 10459 27523
rect 21741 27489 21775 27523
rect 22201 27489 22235 27523
rect 2145 27421 2179 27455
rect 2237 27421 2271 27455
rect 2421 27421 2455 27455
rect 3433 27421 3467 27455
rect 4905 27421 4939 27455
rect 5089 27421 5123 27455
rect 6837 27421 6871 27455
rect 6929 27421 6963 27455
rect 9321 27421 9355 27455
rect 10701 27421 10735 27455
rect 12357 27421 12391 27455
rect 12624 27421 12658 27455
rect 14105 27421 14139 27455
rect 14473 27421 14507 27455
rect 14749 27421 14783 27455
rect 14933 27421 14967 27455
rect 15025 27421 15059 27455
rect 15117 27421 15151 27455
rect 15393 27421 15427 27455
rect 15541 27421 15575 27455
rect 15669 27421 15703 27455
rect 15761 27421 15795 27455
rect 15899 27421 15933 27455
rect 16129 27421 16163 27455
rect 19625 27421 19659 27455
rect 20269 27421 20303 27455
rect 20637 27421 20671 27455
rect 20913 27421 20947 27455
rect 23673 27421 23707 27455
rect 23949 27421 23983 27455
rect 6592 27353 6626 27387
rect 7196 27353 7230 27387
rect 12081 27353 12115 27387
rect 14289 27353 14323 27387
rect 14381 27353 14415 27387
rect 16396 27353 16430 27387
rect 17693 27353 17727 27387
rect 18521 27353 18555 27387
rect 18705 27353 18739 27387
rect 19809 27353 19843 27387
rect 20453 27353 20487 27387
rect 21097 27353 21131 27387
rect 21281 27353 21315 27387
rect 23428 27353 23462 27387
rect 2145 27285 2179 27319
rect 3341 27285 3375 27319
rect 3801 27285 3835 27319
rect 4169 27285 4203 27319
rect 4261 27285 4295 27319
rect 5457 27285 5491 27319
rect 8309 27285 8343 27319
rect 13737 27285 13771 27319
rect 15301 27285 15335 27319
rect 16037 27285 16071 27319
rect 22293 27285 22327 27319
rect 23765 27285 23799 27319
rect 1777 27081 1811 27115
rect 1869 27081 1903 27115
rect 2697 27081 2731 27115
rect 5181 27081 5215 27115
rect 9781 27081 9815 27115
rect 10701 27081 10735 27115
rect 13461 27081 13495 27115
rect 15393 27081 15427 27115
rect 4169 27013 4203 27047
rect 5349 27013 5383 27047
rect 5549 27013 5583 27047
rect 13798 27013 13832 27047
rect 17049 27013 17083 27047
rect 19349 27013 19383 27047
rect 1409 26945 1443 26979
rect 1869 26945 1903 26979
rect 2973 26945 3007 26979
rect 3065 26945 3099 26979
rect 3341 26945 3375 26979
rect 3525 26945 3559 26979
rect 4077 26945 4111 26979
rect 5825 26945 5859 26979
rect 6009 26945 6043 26979
rect 7757 26945 7791 26979
rect 8033 26945 8067 26979
rect 9321 26945 9355 26979
rect 10425 26945 10459 26979
rect 10609 26945 10643 26979
rect 11713 26945 11747 26979
rect 11980 26945 12014 26979
rect 13277 26945 13311 26979
rect 15577 26945 15611 26979
rect 15761 26945 15795 26979
rect 16681 26945 16715 26979
rect 16829 26945 16863 26979
rect 16957 26945 16991 26979
rect 17146 26945 17180 26979
rect 19165 26945 19199 26979
rect 19708 26945 19742 26979
rect 24234 26945 24268 26979
rect 24501 26945 24535 26979
rect 1777 26877 1811 26911
rect 2237 26877 2271 26911
rect 2329 26877 2363 26911
rect 6469 26877 6503 26911
rect 7941 26877 7975 26911
rect 9689 26877 9723 26911
rect 9873 26877 9907 26911
rect 13553 26877 13587 26911
rect 19441 26877 19475 26911
rect 22569 26877 22603 26911
rect 2697 26809 2731 26843
rect 3249 26809 3283 26843
rect 7573 26809 7607 26843
rect 10241 26809 10275 26843
rect 22937 26809 22971 26843
rect 5365 26741 5399 26775
rect 6193 26741 6227 26775
rect 7021 26741 7055 26775
rect 7757 26741 7791 26775
rect 9413 26741 9447 26775
rect 13093 26741 13127 26775
rect 14933 26741 14967 26775
rect 17325 26741 17359 26775
rect 18981 26741 19015 26775
rect 20821 26741 20855 26775
rect 23029 26741 23063 26775
rect 23121 26741 23155 26775
rect 4721 26537 4755 26571
rect 4905 26537 4939 26571
rect 6837 26537 6871 26571
rect 9965 26537 9999 26571
rect 11989 26537 12023 26571
rect 12725 26537 12759 26571
rect 16589 26537 16623 26571
rect 19717 26537 19751 26571
rect 23581 26537 23615 26571
rect 4077 26469 4111 26503
rect 12633 26469 12667 26503
rect 13185 26469 13219 26503
rect 17417 26469 17451 26503
rect 20729 26469 20763 26503
rect 6009 26401 6043 26435
rect 9505 26401 9539 26435
rect 3985 26333 4019 26367
rect 4353 26333 4387 26367
rect 4537 26333 4571 26367
rect 5549 26333 5583 26367
rect 5917 26333 5951 26367
rect 6193 26333 6227 26367
rect 6377 26333 6411 26367
rect 6653 26333 6687 26367
rect 6929 26333 6963 26367
rect 7113 26333 7147 26367
rect 12173 26333 12207 26367
rect 15761 26333 15795 26367
rect 16773 26333 16807 26367
rect 17233 26333 17267 26367
rect 17509 26333 17543 26367
rect 17765 26333 17799 26367
rect 19533 26333 19567 26367
rect 22109 26333 22143 26367
rect 23397 26333 23431 26367
rect 3433 26265 3467 26299
rect 4905 26265 4939 26299
rect 5089 26265 5123 26299
rect 7021 26265 7055 26299
rect 9413 26265 9447 26299
rect 9505 26265 9539 26299
rect 12265 26265 12299 26299
rect 12817 26265 12851 26299
rect 21842 26265 21876 26299
rect 2145 26197 2179 26231
rect 6469 26197 6503 26231
rect 13277 26197 13311 26231
rect 15577 26197 15611 26231
rect 18889 26197 18923 26231
rect 3985 25993 4019 26027
rect 4353 25993 4387 26027
rect 7665 25993 7699 26027
rect 15761 25993 15795 26027
rect 17417 25993 17451 26027
rect 18705 25993 18739 26027
rect 21465 25993 21499 26027
rect 2651 25925 2685 25959
rect 2973 25925 3007 25959
rect 8861 25925 8895 25959
rect 16957 25925 16991 25959
rect 18061 25925 18095 25959
rect 19042 25925 19076 25959
rect 21833 25925 21867 25959
rect 2145 25857 2179 25891
rect 2329 25857 2363 25891
rect 2421 25857 2455 25891
rect 2513 25857 2547 25891
rect 3249 25857 3283 25891
rect 3525 25857 3559 25891
rect 3893 25857 3927 25891
rect 4813 25857 4847 25891
rect 5089 25857 5123 25891
rect 7205 25857 7239 25891
rect 7389 25857 7423 25891
rect 7481 25857 7515 25891
rect 7849 25857 7883 25891
rect 7941 25857 7975 25891
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 8769 25857 8803 25891
rect 9689 25857 9723 25891
rect 10241 25857 10275 25891
rect 10333 25857 10367 25891
rect 10517 25857 10551 25891
rect 13093 25857 13127 25891
rect 16129 25857 16163 25891
rect 16221 25857 16255 25891
rect 18245 25857 18279 25891
rect 18521 25857 18555 25891
rect 21281 25857 21315 25891
rect 22017 25857 22051 25891
rect 2789 25789 2823 25823
rect 2881 25789 2915 25823
rect 3433 25789 3467 25823
rect 4445 25789 4479 25823
rect 4629 25789 4663 25823
rect 9965 25789 9999 25823
rect 15301 25789 15335 25823
rect 18797 25789 18831 25823
rect 22201 25789 22235 25823
rect 15669 25721 15703 25755
rect 17325 25721 17359 25755
rect 3525 25653 3559 25687
rect 4905 25653 4939 25687
rect 5273 25653 5307 25687
rect 7021 25653 7055 25687
rect 9505 25653 9539 25687
rect 9873 25653 9907 25687
rect 10149 25653 10183 25687
rect 10425 25653 10459 25687
rect 12909 25653 12943 25687
rect 15945 25653 15979 25687
rect 16405 25653 16439 25687
rect 20177 25653 20211 25687
rect 4629 25449 4663 25483
rect 10977 25449 11011 25483
rect 19257 25449 19291 25483
rect 25789 25449 25823 25483
rect 7849 25381 7883 25415
rect 10149 25381 10183 25415
rect 11253 25381 11287 25415
rect 12081 25381 12115 25415
rect 14473 25381 14507 25415
rect 23765 25381 23799 25415
rect 2513 25313 2547 25347
rect 5181 25313 5215 25347
rect 7205 25313 7239 25347
rect 8953 25313 8987 25347
rect 11069 25313 11103 25347
rect 11161 25313 11195 25347
rect 11529 25313 11563 25347
rect 11989 25313 12023 25347
rect 12541 25313 12575 25347
rect 14565 25313 14599 25347
rect 22201 25313 22235 25347
rect 3065 25245 3099 25279
rect 3341 25245 3375 25279
rect 3525 25245 3559 25279
rect 3801 25245 3835 25279
rect 3985 25245 4019 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 4997 25245 5031 25279
rect 5089 25245 5123 25279
rect 5457 25245 5491 25279
rect 5641 25245 5675 25279
rect 6377 25245 6411 25279
rect 6469 25245 6503 25279
rect 6653 25245 6687 25279
rect 6745 25245 6779 25279
rect 7297 25245 7331 25279
rect 7665 25245 7699 25279
rect 7757 25245 7791 25279
rect 8125 25245 8159 25279
rect 8309 25245 8343 25279
rect 8585 25245 8619 25279
rect 8769 25245 8803 25279
rect 9321 25245 9355 25279
rect 9597 25245 9631 25279
rect 9781 25245 9815 25279
rect 10333 25245 10367 25279
rect 10425 25245 10459 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 10793 25245 10827 25279
rect 10885 25245 10919 25279
rect 11437 25245 11471 25279
rect 11713 25245 11747 25279
rect 11897 25245 11931 25279
rect 12081 25245 12115 25279
rect 12265 25245 12299 25279
rect 12808 25245 12842 25279
rect 14841 25245 14875 25279
rect 15393 25245 15427 25279
rect 15660 25245 15694 25279
rect 16865 25245 16899 25279
rect 17325 25245 17359 25279
rect 19625 25245 19659 25279
rect 20729 25245 20763 25279
rect 24409 25245 24443 25279
rect 6193 25177 6227 25211
rect 14105 25177 14139 25211
rect 17049 25177 17083 25211
rect 17592 25177 17626 25211
rect 19441 25177 19475 25211
rect 20996 25177 21030 25211
rect 22468 25177 22502 25211
rect 24133 25177 24167 25211
rect 24654 25177 24688 25211
rect 5549 25109 5583 25143
rect 7021 25109 7055 25143
rect 7389 25109 7423 25143
rect 7573 25109 7607 25143
rect 8953 25109 8987 25143
rect 13921 25109 13955 25143
rect 14657 25109 14691 25143
rect 16773 25109 16807 25143
rect 17233 25109 17267 25143
rect 18705 25109 18739 25143
rect 22109 25109 22143 25143
rect 23581 25109 23615 25143
rect 23673 25109 23707 25143
rect 4537 24905 4571 24939
rect 4905 24905 4939 24939
rect 8217 24905 8251 24939
rect 12173 24905 12207 24939
rect 17785 24905 17819 24939
rect 21281 24905 21315 24939
rect 22477 24905 22511 24939
rect 23949 24905 23983 24939
rect 2237 24837 2271 24871
rect 2421 24837 2455 24871
rect 9321 24837 9355 24871
rect 10609 24837 10643 24871
rect 10809 24837 10843 24871
rect 14280 24837 14314 24871
rect 16957 24837 16991 24871
rect 21833 24837 21867 24871
rect 1685 24769 1719 24803
rect 1961 24769 1995 24803
rect 2697 24769 2731 24803
rect 5641 24769 5675 24803
rect 5733 24769 5767 24803
rect 5917 24769 5951 24803
rect 6009 24769 6043 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 6837 24769 6871 24803
rect 6929 24769 6963 24803
rect 8401 24769 8435 24803
rect 8493 24769 8527 24803
rect 8677 24769 8711 24803
rect 9137 24769 9171 24803
rect 9413 24769 9447 24803
rect 10057 24769 10091 24803
rect 10149 24769 10183 24803
rect 10241 24769 10275 24803
rect 10425 24769 10459 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 11897 24769 11931 24803
rect 12081 24769 12115 24803
rect 14013 24769 14047 24803
rect 16681 24769 16715 24803
rect 16865 24769 16899 24803
rect 17049 24769 17083 24803
rect 17325 24769 17359 24803
rect 17509 24769 17543 24803
rect 17693 24769 17727 24803
rect 17969 24769 18003 24803
rect 18981 24769 19015 24803
rect 19513 24769 19547 24803
rect 20729 24769 20763 24803
rect 21465 24769 21499 24803
rect 22017 24769 22051 24803
rect 22201 24769 22235 24803
rect 22293 24769 22327 24803
rect 23765 24769 23799 24803
rect 4997 24701 5031 24735
rect 5181 24701 5215 24735
rect 6377 24701 6411 24735
rect 7297 24701 7331 24735
rect 7757 24701 7791 24735
rect 8585 24701 8619 24735
rect 9781 24701 9815 24735
rect 15945 24701 15979 24735
rect 19257 24701 19291 24735
rect 21189 24701 21223 24735
rect 25237 24701 25271 24735
rect 1869 24633 1903 24667
rect 7481 24633 7515 24667
rect 8953 24633 8987 24667
rect 10977 24633 11011 24667
rect 15393 24633 15427 24667
rect 15669 24633 15703 24667
rect 19165 24633 19199 24667
rect 21005 24633 21039 24667
rect 24961 24633 24995 24667
rect 2237 24565 2271 24599
rect 3985 24565 4019 24599
rect 5457 24565 5491 24599
rect 10793 24565 10827 24599
rect 15485 24565 15519 24599
rect 17233 24565 17267 24599
rect 20637 24565 20671 24599
rect 24777 24565 24811 24599
rect 2605 24361 2639 24395
rect 3525 24361 3559 24395
rect 4905 24361 4939 24395
rect 10057 24361 10091 24395
rect 15669 24361 15703 24395
rect 19257 24361 19291 24395
rect 6193 24293 6227 24327
rect 6929 24293 6963 24327
rect 13553 24293 13587 24327
rect 23397 24293 23431 24327
rect 1409 24225 1443 24259
rect 3157 24225 3191 24259
rect 3617 24225 3651 24259
rect 4445 24225 4479 24259
rect 10977 24225 11011 24259
rect 11805 24225 11839 24259
rect 13645 24225 13679 24259
rect 23581 24225 23615 24259
rect 1869 24157 1903 24191
rect 2237 24157 2271 24191
rect 2329 24157 2363 24191
rect 3341 24157 3375 24191
rect 3433 24157 3467 24191
rect 5089 24157 5123 24191
rect 5273 24157 5307 24191
rect 5457 24157 5491 24191
rect 5549 24157 5583 24191
rect 5917 24157 5951 24191
rect 6101 24157 6135 24191
rect 6469 24157 6503 24191
rect 6929 24157 6963 24191
rect 7021 24157 7055 24191
rect 7205 24157 7239 24191
rect 7481 24157 7515 24191
rect 7665 24157 7699 24191
rect 9597 24157 9631 24191
rect 10241 24157 10275 24191
rect 10333 24157 10367 24191
rect 10425 24157 10459 24191
rect 10609 24157 10643 24191
rect 11897 24157 11931 24191
rect 12265 24157 12299 24191
rect 12541 24157 12575 24191
rect 13921 24157 13955 24191
rect 15117 24157 15151 24191
rect 17325 24157 17359 24191
rect 19625 24157 19659 24191
rect 22661 24157 22695 24191
rect 23029 24157 23063 24191
rect 23673 24157 23707 24191
rect 24409 24157 24443 24191
rect 2881 24089 2915 24123
rect 5181 24089 5215 24123
rect 6193 24089 6227 24123
rect 7297 24089 7331 24123
rect 9413 24089 9447 24123
rect 9873 24089 9907 24123
rect 12173 24089 12207 24123
rect 13185 24089 13219 24123
rect 15653 24089 15687 24123
rect 15853 24089 15887 24123
rect 17592 24089 17626 24123
rect 19441 24089 19475 24123
rect 22753 24089 22787 24123
rect 22845 24089 22879 24123
rect 23121 24089 23155 24123
rect 24654 24089 24688 24123
rect 3065 24021 3099 24055
rect 3801 24021 3835 24055
rect 4169 24021 4203 24055
rect 4261 24021 4295 24055
rect 5641 24021 5675 24055
rect 6377 24021 6411 24055
rect 7665 24021 7699 24055
rect 9781 24021 9815 24055
rect 13737 24021 13771 24055
rect 14933 24021 14967 24055
rect 15485 24021 15519 24055
rect 18705 24021 18739 24055
rect 22477 24021 22511 24055
rect 23857 24021 23891 24055
rect 25789 24021 25823 24055
rect 3617 23817 3651 23851
rect 4537 23817 4571 23851
rect 4721 23817 4755 23851
rect 5365 23817 5399 23851
rect 6745 23817 6779 23851
rect 10333 23817 10367 23851
rect 12909 23817 12943 23851
rect 16129 23817 16163 23851
rect 17509 23817 17543 23851
rect 19825 23817 19859 23851
rect 21465 23817 21499 23851
rect 23213 23817 23247 23851
rect 24869 23817 24903 23851
rect 6377 23749 6411 23783
rect 7297 23749 7331 23783
rect 10701 23749 10735 23783
rect 13360 23749 13394 23783
rect 14924 23749 14958 23783
rect 18857 23749 18891 23783
rect 19073 23749 19107 23783
rect 19625 23749 19659 23783
rect 20545 23749 20579 23783
rect 22078 23749 22112 23783
rect 23581 23749 23615 23783
rect 23673 23749 23707 23783
rect 25206 23749 25240 23783
rect 1961 23681 1995 23715
rect 2145 23681 2179 23715
rect 2237 23681 2271 23715
rect 2329 23681 2363 23715
rect 2513 23681 2547 23715
rect 3801 23681 3835 23715
rect 3985 23681 4019 23715
rect 4169 23681 4203 23715
rect 4353 23681 4387 23715
rect 4718 23681 4752 23715
rect 6837 23681 6871 23715
rect 7113 23681 7147 23715
rect 7205 23681 7239 23715
rect 7481 23681 7515 23715
rect 7573 23681 7607 23715
rect 7757 23681 7791 23715
rect 8309 23681 8343 23715
rect 10517 23681 10551 23715
rect 10793 23681 10827 23715
rect 11069 23681 11103 23715
rect 11161 23681 11195 23715
rect 12817 23681 12851 23715
rect 13093 23681 13127 23715
rect 14657 23681 14691 23715
rect 16313 23681 16347 23715
rect 17325 23681 17359 23715
rect 21281 23681 21315 23715
rect 21833 23681 21867 23715
rect 23484 23681 23518 23715
rect 23801 23681 23835 23715
rect 23949 23681 23983 23715
rect 24685 23681 24719 23715
rect 4077 23613 4111 23647
rect 5181 23613 5215 23647
rect 5549 23613 5583 23647
rect 5641 23613 5675 23647
rect 5733 23613 5767 23647
rect 5825 23613 5859 23647
rect 6469 23613 6503 23647
rect 16497 23613 16531 23647
rect 16773 23613 16807 23647
rect 17233 23613 17267 23647
rect 24961 23613 24995 23647
rect 6929 23545 6963 23579
rect 17049 23545 17083 23579
rect 2421 23477 2455 23511
rect 5089 23477 5123 23511
rect 6561 23477 6595 23511
rect 7573 23477 7607 23511
rect 9597 23477 9631 23511
rect 10885 23477 10919 23511
rect 14473 23477 14507 23511
rect 16037 23477 16071 23511
rect 18705 23477 18739 23511
rect 18889 23477 18923 23511
rect 19809 23477 19843 23511
rect 19993 23477 20027 23511
rect 20821 23477 20855 23511
rect 23305 23477 23339 23511
rect 26341 23477 26375 23511
rect 5089 23273 5123 23307
rect 5825 23273 5859 23307
rect 8125 23273 8159 23307
rect 8309 23273 8343 23307
rect 9413 23273 9447 23307
rect 9597 23273 9631 23307
rect 10517 23273 10551 23307
rect 11253 23273 11287 23307
rect 14473 23273 14507 23307
rect 15577 23273 15611 23307
rect 18797 23273 18831 23307
rect 19441 23273 19475 23307
rect 19993 23273 20027 23307
rect 21465 23273 21499 23307
rect 23029 23273 23063 23307
rect 7389 23205 7423 23239
rect 8401 23205 8435 23239
rect 10057 23205 10091 23239
rect 14657 23205 14691 23239
rect 15669 23205 15703 23239
rect 15945 23205 15979 23239
rect 19257 23205 19291 23239
rect 20177 23205 20211 23239
rect 5733 23137 5767 23171
rect 5917 23137 5951 23171
rect 9229 23137 9263 23171
rect 18337 23137 18371 23171
rect 2329 23069 2363 23103
rect 2881 23069 2915 23103
rect 3065 23069 3099 23103
rect 3249 23069 3283 23103
rect 3801 23069 3835 23103
rect 6009 23069 6043 23103
rect 8401 23069 8435 23103
rect 8677 23069 8711 23103
rect 9137 23069 9171 23103
rect 9965 23069 9999 23103
rect 10057 23069 10091 23103
rect 10149 23069 10183 23103
rect 10333 23069 10367 23103
rect 10425 23069 10459 23103
rect 10609 23069 10643 23103
rect 10885 23069 10919 23103
rect 11069 23069 11103 23103
rect 12541 23069 12575 23103
rect 15209 23069 15243 23103
rect 15393 23069 15427 23103
rect 15485 23069 15519 23103
rect 16129 23069 16163 23103
rect 16221 23069 16255 23103
rect 17141 23069 17175 23103
rect 17325 23069 17359 23103
rect 17509 23069 17543 23103
rect 18061 23069 18095 23103
rect 18153 23069 18187 23103
rect 22293 23069 22327 23103
rect 22386 23069 22420 23103
rect 22569 23069 22603 23103
rect 22799 23069 22833 23103
rect 23213 23069 23247 23103
rect 23397 23069 23431 23103
rect 23581 23069 23615 23103
rect 24409 23069 24443 23103
rect 2605 23001 2639 23035
rect 6101 23001 6135 23035
rect 7941 23001 7975 23035
rect 9781 23001 9815 23035
rect 12808 23001 12842 23035
rect 14289 23001 14323 23035
rect 17233 23001 17267 23035
rect 18613 23001 18647 23035
rect 19579 23001 19613 23035
rect 19809 23001 19843 23035
rect 21097 23001 21131 23035
rect 21281 23001 21315 23035
rect 22661 23001 22695 23035
rect 23305 23001 23339 23035
rect 24654 23001 24688 23035
rect 8151 22933 8185 22967
rect 8585 22933 8619 22967
rect 13921 22933 13955 22967
rect 14499 22933 14533 22967
rect 16405 22933 16439 22967
rect 16957 22933 16991 22967
rect 18813 22933 18847 22967
rect 18981 22933 19015 22967
rect 19425 22933 19459 22967
rect 20019 22933 20053 22967
rect 22937 22933 22971 22967
rect 25789 22933 25823 22967
rect 2513 22729 2547 22763
rect 2605 22729 2639 22763
rect 3893 22729 3927 22763
rect 5457 22729 5491 22763
rect 9045 22729 9079 22763
rect 11529 22729 11563 22763
rect 12449 22729 12483 22763
rect 12909 22729 12943 22763
rect 15393 22729 15427 22763
rect 19717 22729 19751 22763
rect 23949 22729 23983 22763
rect 1961 22661 1995 22695
rect 2237 22661 2271 22695
rect 6837 22661 6871 22695
rect 6929 22661 6963 22695
rect 7665 22661 7699 22695
rect 15025 22661 15059 22695
rect 15241 22661 15275 22695
rect 20054 22661 20088 22695
rect 24501 22661 24535 22695
rect 25237 22661 25271 22695
rect 1593 22593 1627 22627
rect 2421 22593 2455 22627
rect 2789 22593 2823 22627
rect 3157 22593 3191 22627
rect 3249 22593 3283 22627
rect 3341 22593 3375 22627
rect 3525 22593 3559 22627
rect 5365 22593 5399 22627
rect 5733 22593 5767 22627
rect 5825 22593 5859 22627
rect 5917 22593 5951 22627
rect 6101 22593 6135 22627
rect 6740 22593 6774 22627
rect 7057 22593 7091 22627
rect 7205 22593 7239 22627
rect 7849 22593 7883 22627
rect 7941 22593 7975 22627
rect 8125 22593 8159 22627
rect 8217 22593 8251 22627
rect 8493 22593 8527 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 9137 22593 9171 22627
rect 11989 22593 12023 22627
rect 12081 22593 12115 22627
rect 12240 22593 12274 22627
rect 12357 22593 12391 22627
rect 12541 22593 12575 22627
rect 12725 22593 12759 22627
rect 13369 22593 13403 22627
rect 13461 22593 13495 22627
rect 16957 22593 16991 22627
rect 18889 22593 18923 22627
rect 19073 22593 19107 22627
rect 19165 22593 19199 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 23213 22593 23247 22627
rect 23765 22593 23799 22627
rect 2881 22525 2915 22559
rect 11621 22525 11655 22559
rect 11713 22525 11747 22559
rect 16773 22525 16807 22559
rect 18981 22525 19015 22559
rect 19809 22525 19843 22559
rect 23673 22525 23707 22559
rect 6561 22457 6595 22491
rect 8585 22457 8619 22491
rect 13185 22457 13219 22491
rect 23489 22457 23523 22491
rect 24869 22457 24903 22491
rect 25605 22457 25639 22491
rect 1961 22389 1995 22423
rect 2145 22389 2179 22423
rect 8309 22389 8343 22423
rect 11897 22389 11931 22423
rect 12173 22389 12207 22423
rect 13645 22389 13679 22423
rect 15209 22389 15243 22423
rect 17141 22389 17175 22423
rect 18613 22389 18647 22423
rect 21189 22389 21223 22423
rect 24961 22389 24995 22423
rect 25697 22389 25731 22423
rect 8309 22185 8343 22219
rect 10793 22185 10827 22219
rect 11529 22185 11563 22219
rect 12081 22185 12115 22219
rect 12265 22185 12299 22219
rect 17877 22185 17911 22219
rect 19625 22185 19659 22219
rect 22753 22185 22787 22219
rect 22845 22185 22879 22219
rect 23489 22185 23523 22219
rect 2697 22117 2731 22151
rect 4169 22117 4203 22151
rect 4537 22049 4571 22083
rect 5641 22049 5675 22083
rect 6193 22049 6227 22083
rect 11437 22049 11471 22083
rect 16037 22049 16071 22083
rect 16129 22049 16163 22083
rect 23213 22049 23247 22083
rect 1593 21981 1627 22015
rect 1777 21981 1811 22015
rect 1869 21981 1903 22015
rect 2513 21981 2547 22015
rect 3893 21981 3927 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 4445 21981 4479 22015
rect 4629 21981 4663 22015
rect 4813 21981 4847 22015
rect 5273 21981 5307 22015
rect 5549 21981 5583 22015
rect 5825 21981 5859 22015
rect 6009 21981 6043 22015
rect 6101 21981 6135 22015
rect 6377 21981 6411 22015
rect 6561 21981 6595 22015
rect 6653 21981 6687 22015
rect 10517 21981 10551 22015
rect 10977 21981 11011 22015
rect 11069 21981 11103 22015
rect 11161 21981 11195 22015
rect 11713 21981 11747 22015
rect 11989 21981 12023 22015
rect 12817 21981 12851 22015
rect 13461 21981 13495 22015
rect 14841 21981 14875 22015
rect 15853 21981 15887 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 19901 21981 19935 22015
rect 20361 21981 20395 22015
rect 20545 21981 20579 22015
rect 20821 21981 20855 22015
rect 21373 21981 21407 22015
rect 23029 21981 23063 22015
rect 24593 21981 24627 22015
rect 26249 21981 26283 22015
rect 26341 21981 26375 22015
rect 1409 21913 1443 21947
rect 2053 21913 2087 21947
rect 4169 21913 4203 21947
rect 5089 21913 5123 21947
rect 7021 21913 7055 21947
rect 10333 21913 10367 21947
rect 10701 21913 10735 21947
rect 11279 21913 11313 21947
rect 12449 21913 12483 21947
rect 13185 21913 13219 21947
rect 16396 21913 16430 21947
rect 17845 21913 17879 21947
rect 18061 21913 18095 21947
rect 19717 21913 19751 21947
rect 20085 21913 20119 21947
rect 20177 21913 20211 21947
rect 21618 21913 21652 21947
rect 23673 21913 23707 21947
rect 25982 21913 26016 21947
rect 26586 21913 26620 21947
rect 2145 21845 2179 21879
rect 4997 21845 5031 21879
rect 5457 21845 5491 21879
rect 11897 21845 11931 21879
rect 12249 21845 12283 21879
rect 13645 21845 13679 21879
rect 14657 21845 14691 21879
rect 15669 21845 15703 21879
rect 17509 21845 17543 21879
rect 17693 21845 17727 21879
rect 20637 21845 20671 21879
rect 23305 21845 23339 21879
rect 23463 21845 23497 21879
rect 24777 21845 24811 21879
rect 24869 21845 24903 21879
rect 27721 21845 27755 21879
rect 2697 21641 2731 21675
rect 3709 21641 3743 21675
rect 5641 21641 5675 21675
rect 6009 21641 6043 21675
rect 6469 21641 6503 21675
rect 8585 21641 8619 21675
rect 9505 21641 9539 21675
rect 12081 21641 12115 21675
rect 16681 21641 16715 21675
rect 19191 21641 19225 21675
rect 25973 21641 26007 21675
rect 2191 21573 2225 21607
rect 2778 21573 2812 21607
rect 2881 21573 2915 21607
rect 3249 21573 3283 21607
rect 4077 21573 4111 21607
rect 6193 21573 6227 21607
rect 6745 21573 6779 21607
rect 6837 21573 6871 21607
rect 7205 21573 7239 21607
rect 14810 21573 14844 21607
rect 16037 21573 16071 21607
rect 18981 21573 19015 21607
rect 20352 21573 20386 21607
rect 21925 21573 21959 21607
rect 22141 21573 22175 21607
rect 23213 21573 23247 21607
rect 1777 21505 1811 21539
rect 2421 21505 2455 21539
rect 2513 21505 2547 21539
rect 3157 21505 3191 21539
rect 3341 21505 3375 21539
rect 3888 21505 3922 21539
rect 3985 21505 4019 21539
rect 4260 21505 4294 21539
rect 4353 21505 4387 21539
rect 4629 21505 4663 21539
rect 5549 21505 5583 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6607 21505 6641 21539
rect 6965 21505 6999 21539
rect 7113 21505 7147 21539
rect 7389 21505 7423 21539
rect 7481 21505 7515 21539
rect 7665 21505 7699 21539
rect 7757 21505 7791 21539
rect 7941 21505 7975 21539
rect 8125 21505 8159 21539
rect 8217 21505 8251 21539
rect 8493 21505 8527 21539
rect 8677 21505 8711 21539
rect 8769 21505 8803 21539
rect 8953 21505 8987 21539
rect 9321 21505 9355 21539
rect 9781 21505 9815 21539
rect 10057 21505 10091 21539
rect 10241 21505 10275 21539
rect 10517 21505 10551 21539
rect 10701 21505 10735 21539
rect 10977 21505 11011 21539
rect 11529 21505 11563 21539
rect 12357 21505 12391 21539
rect 12909 21505 12943 21539
rect 13176 21505 13210 21539
rect 16221 21505 16255 21539
rect 16405 21505 16439 21539
rect 16865 21505 16899 21539
rect 17509 21505 17543 21539
rect 17785 21505 17819 21539
rect 18153 21505 18187 21539
rect 18613 21505 18647 21539
rect 19533 21505 19567 21539
rect 22937 21505 22971 21539
rect 23121 21505 23155 21539
rect 25789 21505 25823 21539
rect 4445 21437 4479 21471
rect 4905 21437 4939 21471
rect 6120 21437 6154 21471
rect 9137 21437 9171 21471
rect 9597 21437 9631 21471
rect 11805 21437 11839 21471
rect 14565 21437 14599 21471
rect 17601 21437 17635 21471
rect 19717 21437 19751 21471
rect 20085 21437 20119 21471
rect 3065 21369 3099 21403
rect 5825 21369 5859 21403
rect 7941 21369 7975 21403
rect 9873 21369 9907 21403
rect 9965 21369 9999 21403
rect 10609 21369 10643 21403
rect 15945 21369 15979 21403
rect 22293 21369 22327 21403
rect 22753 21369 22787 21403
rect 23489 21369 23523 21403
rect 2145 21301 2179 21335
rect 4813 21301 4847 21335
rect 8861 21301 8895 21335
rect 11621 21301 11655 21335
rect 12541 21301 12575 21335
rect 14289 21301 14323 21335
rect 17969 21301 18003 21335
rect 18337 21301 18371 21335
rect 18705 21301 18739 21335
rect 19165 21301 19199 21335
rect 19349 21301 19383 21335
rect 21465 21301 21499 21335
rect 22109 21301 22143 21335
rect 22385 21301 22419 21335
rect 22661 21301 22695 21335
rect 22845 21301 22879 21335
rect 23673 21301 23707 21335
rect 2237 21097 2271 21131
rect 4721 21097 4755 21131
rect 7021 21097 7055 21131
rect 8585 21097 8619 21131
rect 8769 21097 8803 21131
rect 9137 21097 9171 21131
rect 13369 21097 13403 21131
rect 14933 21097 14967 21131
rect 15209 21097 15243 21131
rect 15853 21097 15887 21131
rect 17141 21097 17175 21131
rect 18705 21097 18739 21131
rect 19533 21097 19567 21131
rect 20545 21097 20579 21131
rect 21465 21097 21499 21131
rect 22845 21097 22879 21131
rect 23029 21097 23063 21131
rect 3157 21029 3191 21063
rect 10885 21029 10919 21063
rect 19625 21029 19659 21063
rect 24961 21029 24995 21063
rect 2697 20961 2731 20995
rect 3249 20961 3283 20995
rect 7113 20961 7147 20995
rect 8217 20961 8251 20995
rect 9689 20961 9723 20995
rect 11161 20961 11195 20995
rect 12081 20961 12115 20995
rect 19073 20961 19107 20995
rect 24593 20961 24627 20995
rect 25053 20961 25087 20995
rect 2053 20893 2087 20927
rect 2329 20893 2363 20927
rect 2881 20893 2915 20927
rect 4859 20893 4893 20927
rect 5227 20893 5261 20927
rect 5365 20893 5399 20927
rect 6650 20893 6684 20927
rect 7343 20893 7377 20927
rect 7481 20893 7515 20927
rect 7701 20893 7735 20927
rect 7849 20893 7883 20927
rect 9505 20893 9539 20927
rect 10333 20893 10367 20927
rect 10701 20893 10735 20927
rect 11253 20893 11287 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 14749 20893 14783 20927
rect 15025 20893 15059 20927
rect 18889 20893 18923 20927
rect 19254 20893 19288 20927
rect 19717 20893 19751 20927
rect 20821 20893 20855 20927
rect 21189 20893 21223 20927
rect 21281 20893 21315 20927
rect 23581 20893 23615 20927
rect 25237 20893 25271 20927
rect 4997 20825 5031 20859
rect 5089 20825 5123 20859
rect 7573 20825 7607 20859
rect 10517 20825 10551 20859
rect 10609 20825 10643 20859
rect 12909 20825 12943 20859
rect 14565 20825 14599 20859
rect 15669 20825 15703 20859
rect 16957 20825 16991 20859
rect 20361 20825 20395 20859
rect 21005 20825 21039 20859
rect 23213 20825 23247 20859
rect 1869 20757 1903 20791
rect 6469 20757 6503 20791
rect 6653 20757 6687 20791
rect 7205 20757 7239 20791
rect 8585 20757 8619 20791
rect 9597 20757 9631 20791
rect 13001 20757 13035 20791
rect 14105 20757 14139 20791
rect 15869 20757 15903 20791
rect 16037 20757 16071 20791
rect 17157 20757 17191 20791
rect 17325 20757 17359 20791
rect 19349 20757 19383 20791
rect 19993 20757 20027 20791
rect 20561 20757 20595 20791
rect 20729 20757 20763 20791
rect 23003 20757 23037 20791
rect 23765 20757 23799 20791
rect 25421 20757 25455 20791
rect 3249 20553 3283 20587
rect 3893 20553 3927 20587
rect 5181 20553 5215 20587
rect 7665 20553 7699 20587
rect 10977 20553 11011 20587
rect 16329 20553 16363 20587
rect 18981 20553 19015 20587
rect 23397 20553 23431 20587
rect 6193 20485 6227 20519
rect 12449 20485 12483 20519
rect 13093 20485 13127 20519
rect 15577 20485 15611 20519
rect 16129 20485 16163 20519
rect 18613 20485 18647 20519
rect 18813 20485 18847 20519
rect 24510 20485 24544 20519
rect 26442 20485 26476 20519
rect 3433 20417 3467 20451
rect 3525 20417 3559 20451
rect 4261 20417 4295 20451
rect 4353 20417 4387 20451
rect 4537 20417 4571 20451
rect 4629 20417 4663 20451
rect 4721 20417 4755 20451
rect 4813 20417 4847 20451
rect 4997 20417 5031 20451
rect 5917 20417 5951 20451
rect 6009 20417 6043 20451
rect 6377 20417 6411 20451
rect 8217 20417 8251 20451
rect 8401 20417 8435 20451
rect 10885 20417 10919 20451
rect 11069 20417 11103 20451
rect 12541 20417 12575 20451
rect 12633 20417 12667 20451
rect 13277 20417 13311 20451
rect 13553 20417 13587 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 14841 20417 14875 20451
rect 15761 20417 15795 20451
rect 17233 20417 17267 20451
rect 17509 20417 17543 20451
rect 20361 20417 20395 20451
rect 21833 20417 21867 20451
rect 22006 20417 22040 20451
rect 22385 20417 22419 20451
rect 22569 20417 22603 20451
rect 22661 20417 22695 20451
rect 24777 20417 24811 20451
rect 26709 20417 26743 20451
rect 2881 20349 2915 20383
rect 2973 20349 3007 20383
rect 3617 20349 3651 20383
rect 13001 20349 13035 20383
rect 17325 20349 17359 20383
rect 22201 20349 22235 20383
rect 8217 20281 8251 20315
rect 14289 20281 14323 20315
rect 25329 20281 25363 20315
rect 3525 20213 3559 20247
rect 4077 20213 4111 20247
rect 6193 20213 6227 20247
rect 14933 20213 14967 20247
rect 15393 20213 15427 20247
rect 16313 20213 16347 20247
rect 16497 20213 16531 20247
rect 17049 20213 17083 20247
rect 17417 20213 17451 20247
rect 18797 20213 18831 20247
rect 20545 20213 20579 20247
rect 22845 20213 22879 20247
rect 3065 20009 3099 20043
rect 3985 20009 4019 20043
rect 4721 20009 4755 20043
rect 5365 20009 5399 20043
rect 8769 20009 8803 20043
rect 8953 20009 8987 20043
rect 9965 20009 9999 20043
rect 10333 20009 10367 20043
rect 11529 20009 11563 20043
rect 14105 20009 14139 20043
rect 17141 20009 17175 20043
rect 17969 20009 18003 20043
rect 18613 20009 18647 20043
rect 20269 20009 20303 20043
rect 21741 20009 21775 20043
rect 4997 19941 5031 19975
rect 17417 19941 17451 19975
rect 17601 19941 17635 19975
rect 18429 19941 18463 19975
rect 2881 19873 2915 19907
rect 4905 19873 4939 19907
rect 5825 19873 5859 19907
rect 5917 19873 5951 19907
rect 9505 19873 9539 19907
rect 10241 19873 10275 19907
rect 10793 19873 10827 19907
rect 10977 19873 11011 19907
rect 11161 19873 11195 19907
rect 14473 19873 14507 19907
rect 23213 19873 23247 19907
rect 1961 19805 1995 19839
rect 2237 19805 2271 19839
rect 2421 19805 2455 19839
rect 2789 19805 2823 19839
rect 3249 19805 3283 19839
rect 3617 19805 3651 19839
rect 3893 19805 3927 19839
rect 3985 19805 4019 19839
rect 4353 19805 4387 19839
rect 4629 19805 4663 19839
rect 5181 19805 5215 19839
rect 5273 19805 5307 19839
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 8585 19805 8619 19839
rect 9873 19805 9907 19839
rect 9965 19805 9999 19839
rect 10701 19805 10735 19839
rect 11345 19805 11379 19839
rect 14289 19805 14323 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 14749 19805 14783 19839
rect 15025 19805 15059 19839
rect 17509 19805 17543 19839
rect 17693 19805 17727 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18245 19805 18279 19839
rect 19257 19805 19291 19839
rect 20361 19805 20395 19839
rect 22946 19805 22980 19839
rect 23765 19805 23799 19839
rect 25789 19805 25823 19839
rect 1501 19737 1535 19771
rect 4997 19737 5031 19771
rect 9321 19737 9355 19771
rect 15270 19737 15304 19771
rect 18797 19737 18831 19771
rect 19901 19737 19935 19771
rect 20085 19737 20119 19771
rect 20628 19737 20662 19771
rect 25522 19737 25556 19771
rect 3433 19669 3467 19703
rect 4905 19669 4939 19703
rect 5733 19669 5767 19703
rect 6929 19669 6963 19703
rect 8401 19669 8435 19703
rect 9413 19669 9447 19703
rect 10057 19669 10091 19703
rect 14933 19669 14967 19703
rect 16405 19669 16439 19703
rect 18587 19669 18621 19703
rect 19441 19669 19475 19703
rect 21833 19669 21867 19703
rect 23581 19669 23615 19703
rect 24409 19669 24443 19703
rect 4353 19465 4387 19499
rect 4629 19465 4663 19499
rect 6561 19465 6595 19499
rect 7481 19465 7515 19499
rect 8217 19465 8251 19499
rect 9682 19465 9716 19499
rect 9965 19465 9999 19499
rect 10517 19465 10551 19499
rect 11345 19465 11379 19499
rect 17509 19465 17543 19499
rect 18613 19465 18647 19499
rect 18981 19465 19015 19499
rect 19901 19465 19935 19499
rect 25145 19465 25179 19499
rect 25421 19465 25455 19499
rect 1409 19397 1443 19431
rect 2421 19397 2455 19431
rect 3249 19397 3283 19431
rect 7573 19397 7607 19431
rect 10425 19397 10459 19431
rect 10977 19397 11011 19431
rect 14381 19397 14415 19431
rect 16037 19397 16071 19431
rect 17672 19397 17706 19431
rect 17877 19397 17911 19431
rect 18245 19397 18279 19431
rect 18461 19397 18495 19431
rect 19441 19397 19475 19431
rect 19809 19397 19843 19431
rect 23480 19397 23514 19431
rect 24685 19397 24719 19431
rect 2789 19329 2823 19363
rect 2881 19329 2915 19363
rect 3525 19329 3559 19363
rect 3617 19329 3651 19363
rect 3709 19329 3743 19363
rect 3893 19329 3927 19363
rect 4169 19329 4203 19363
rect 4445 19329 4479 19363
rect 4767 19329 4801 19363
rect 4905 19329 4939 19363
rect 4997 19329 5031 19363
rect 5125 19329 5159 19363
rect 5273 19329 5307 19363
rect 6377 19329 6411 19363
rect 7297 19329 7331 19363
rect 7849 19329 7883 19363
rect 7941 19329 7975 19363
rect 8033 19329 8067 19363
rect 8217 19329 8251 19363
rect 9505 19329 9539 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 10149 19329 10183 19363
rect 10701 19329 10735 19363
rect 11070 19351 11104 19385
rect 12633 19329 12667 19363
rect 13461 19329 13495 19363
rect 13921 19329 13955 19363
rect 14013 19329 14047 19363
rect 15577 19329 15611 19363
rect 15669 19329 15703 19363
rect 19993 19329 20027 19363
rect 20545 19329 20579 19363
rect 25237 19329 25271 19363
rect 26065 19329 26099 19363
rect 1593 19261 1627 19295
rect 1685 19261 1719 19295
rect 1777 19261 1811 19295
rect 2697 19261 2731 19295
rect 10333 19261 10367 19295
rect 10885 19261 10919 19295
rect 11345 19261 11379 19295
rect 12357 19261 12391 19295
rect 14473 19261 14507 19295
rect 15117 19261 15151 19295
rect 16129 19261 16163 19295
rect 16957 19261 16991 19295
rect 18889 19261 18923 19295
rect 20361 19261 20395 19295
rect 23213 19261 23247 19295
rect 2237 19193 2271 19227
rect 4169 19193 4203 19227
rect 17325 19193 17359 19227
rect 18705 19193 18739 19227
rect 19441 19193 19475 19227
rect 24961 19193 24995 19227
rect 7021 19125 7055 19159
rect 10149 19125 10183 19159
rect 10885 19125 10919 19159
rect 11161 19125 11195 19159
rect 12449 19125 12483 19159
rect 12541 19125 12575 19159
rect 17417 19125 17451 19159
rect 17693 19125 17727 19159
rect 18429 19125 18463 19159
rect 24593 19125 24627 19159
rect 26249 19125 26283 19159
rect 2513 18921 2547 18955
rect 4261 18921 4295 18955
rect 10609 18921 10643 18955
rect 11805 18921 11839 18955
rect 18613 18921 18647 18955
rect 19257 18921 19291 18955
rect 20177 18921 20211 18955
rect 22385 18921 22419 18955
rect 23765 18921 23799 18955
rect 24041 18921 24075 18955
rect 25881 18921 25915 18955
rect 27353 18921 27387 18955
rect 2053 18853 2087 18887
rect 4721 18853 4755 18887
rect 12541 18853 12575 18887
rect 23581 18853 23615 18887
rect 2329 18785 2363 18819
rect 2697 18785 2731 18819
rect 6929 18785 6963 18819
rect 7389 18785 7423 18819
rect 9413 18785 9447 18819
rect 10241 18785 10275 18819
rect 12449 18785 12483 18819
rect 13001 18785 13035 18819
rect 15209 18785 15243 18819
rect 19416 18785 19450 18819
rect 19901 18785 19935 18819
rect 20637 18785 20671 18819
rect 20729 18785 20763 18819
rect 21925 18785 21959 18819
rect 25973 18785 26007 18819
rect 1961 18717 1995 18751
rect 2605 18717 2639 18751
rect 2881 18717 2915 18751
rect 4445 18717 4479 18751
rect 4629 18717 4663 18751
rect 6653 18717 6687 18751
rect 6837 18717 6871 18751
rect 7113 18717 7147 18751
rect 9045 18717 9079 18751
rect 9229 18717 9263 18751
rect 9505 18717 9539 18751
rect 9689 18717 9723 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 10425 18717 10459 18751
rect 10609 18717 10643 18751
rect 11989 18717 12023 18751
rect 12265 18717 12299 18751
rect 12817 18717 12851 18751
rect 13277 18717 13311 18751
rect 13369 18717 13403 18751
rect 13921 18717 13955 18751
rect 14105 18717 14139 18751
rect 14381 18717 14415 18751
rect 14657 18717 14691 18751
rect 15117 18717 15151 18751
rect 15577 18717 15611 18751
rect 16037 18717 16071 18751
rect 16313 18717 16347 18751
rect 17325 18717 17359 18751
rect 21097 18717 21131 18751
rect 21193 18717 21227 18751
rect 22569 18717 22603 18751
rect 22661 18717 22695 18751
rect 25513 18717 25547 18751
rect 26240 18717 26274 18751
rect 3985 18649 4019 18683
rect 4169 18649 4203 18683
rect 8769 18649 8803 18683
rect 12173 18649 12207 18683
rect 13185 18649 13219 18683
rect 15393 18649 15427 18683
rect 18797 18649 18831 18683
rect 20161 18649 20195 18683
rect 20361 18649 20395 18683
rect 21281 18649 21315 18683
rect 21557 18649 21591 18683
rect 22017 18649 22051 18683
rect 22385 18649 22419 18683
rect 23305 18649 23339 18683
rect 24225 18649 24259 18683
rect 25697 18649 25731 18683
rect 1777 18581 1811 18615
rect 13737 18581 13771 18615
rect 14197 18581 14231 18615
rect 15485 18581 15519 18615
rect 15761 18581 15795 18615
rect 16221 18581 16255 18615
rect 17141 18581 17175 18615
rect 18429 18581 18463 18615
rect 18597 18581 18631 18615
rect 19533 18581 19567 18615
rect 19625 18581 19659 18615
rect 19993 18581 20027 18615
rect 21833 18581 21867 18615
rect 22201 18581 22235 18615
rect 22845 18581 22879 18615
rect 23857 18581 23891 18615
rect 24025 18581 24059 18615
rect 1777 18377 1811 18411
rect 2329 18377 2363 18411
rect 3525 18377 3559 18411
rect 4905 18377 4939 18411
rect 5181 18377 5215 18411
rect 7941 18377 7975 18411
rect 9413 18377 9447 18411
rect 9597 18377 9631 18411
rect 11713 18377 11747 18411
rect 12449 18377 12483 18411
rect 13921 18377 13955 18411
rect 21925 18377 21959 18411
rect 22569 18377 22603 18411
rect 24501 18377 24535 18411
rect 25973 18377 26007 18411
rect 26249 18377 26283 18411
rect 14381 18309 14415 18343
rect 14657 18309 14691 18343
rect 15485 18309 15519 18343
rect 15669 18309 15703 18343
rect 16037 18309 16071 18343
rect 16237 18309 16271 18343
rect 17121 18309 17155 18343
rect 20897 18309 20931 18343
rect 21097 18309 21131 18343
rect 22385 18309 22419 18343
rect 24838 18309 24872 18343
rect 27230 18309 27264 18343
rect 2053 18241 2087 18275
rect 2513 18241 2547 18275
rect 2881 18241 2915 18275
rect 2973 18241 3007 18275
rect 3341 18241 3375 18275
rect 3525 18241 3559 18275
rect 3617 18241 3651 18275
rect 3801 18241 3835 18275
rect 4353 18241 4387 18275
rect 5089 18241 5123 18275
rect 5365 18241 5399 18275
rect 5641 18241 5675 18275
rect 5917 18241 5951 18275
rect 6101 18241 6135 18275
rect 6653 18241 6687 18275
rect 8493 18241 8527 18275
rect 8769 18241 8803 18275
rect 8861 18241 8895 18275
rect 9045 18241 9079 18275
rect 9137 18241 9171 18275
rect 9505 18241 9539 18275
rect 9689 18241 9723 18275
rect 11897 18241 11931 18275
rect 12173 18241 12207 18275
rect 12357 18241 12391 18275
rect 12633 18241 12667 18275
rect 12817 18241 12851 18275
rect 14105 18241 14139 18275
rect 14933 18241 14967 18275
rect 15853 18241 15887 18275
rect 16865 18241 16899 18275
rect 18337 18241 18371 18275
rect 18521 18241 18555 18275
rect 19533 18241 19567 18275
rect 22116 18241 22150 18275
rect 22845 18241 22879 18275
rect 23121 18241 23155 18275
rect 23305 18241 23339 18275
rect 24317 18241 24351 18275
rect 26065 18241 26099 18275
rect 26341 18241 26375 18275
rect 26525 18241 26559 18275
rect 26709 18241 26743 18275
rect 2789 18173 2823 18207
rect 6193 18173 6227 18207
rect 6377 18173 6411 18207
rect 9413 18173 9447 18207
rect 12081 18173 12115 18207
rect 14841 18173 14875 18207
rect 18705 18173 18739 18207
rect 22293 18173 22327 18207
rect 23029 18173 23063 18207
rect 24593 18173 24627 18207
rect 26985 18173 27019 18207
rect 11989 18105 12023 18139
rect 14565 18105 14599 18139
rect 20729 18105 20763 18139
rect 3157 18037 3191 18071
rect 8585 18037 8619 18071
rect 9229 18037 9263 18071
rect 14657 18037 14691 18071
rect 15117 18037 15151 18071
rect 16221 18037 16255 18071
rect 16405 18037 16439 18071
rect 18245 18037 18279 18071
rect 19349 18037 19383 18071
rect 20913 18037 20947 18071
rect 22385 18037 22419 18071
rect 22937 18037 22971 18071
rect 28365 18037 28399 18071
rect 1869 17833 1903 17867
rect 3525 17833 3559 17867
rect 4261 17833 4295 17867
rect 10241 17833 10275 17867
rect 10885 17833 10919 17867
rect 11161 17833 11195 17867
rect 13277 17833 13311 17867
rect 14657 17833 14691 17867
rect 16773 17833 16807 17867
rect 19481 17833 19515 17867
rect 23029 17833 23063 17867
rect 24409 17833 24443 17867
rect 28549 17833 28583 17867
rect 4077 17765 4111 17799
rect 5089 17765 5123 17799
rect 7389 17765 7423 17799
rect 8585 17765 8619 17799
rect 9781 17765 9815 17799
rect 9873 17765 9907 17799
rect 10149 17765 10183 17799
rect 10517 17765 10551 17799
rect 14381 17765 14415 17799
rect 16681 17765 16715 17799
rect 19257 17765 19291 17799
rect 23949 17765 23983 17799
rect 26617 17765 26651 17799
rect 9965 17697 9999 17731
rect 10333 17697 10367 17731
rect 10977 17697 11011 17731
rect 13829 17697 13863 17731
rect 14933 17697 14967 17731
rect 16865 17697 16899 17731
rect 2605 17629 2639 17663
rect 3249 17629 3283 17663
rect 3341 17629 3375 17663
rect 3893 17629 3927 17663
rect 4445 17629 4479 17663
rect 4731 17629 4765 17663
rect 4905 17629 4939 17663
rect 5043 17629 5077 17663
rect 7021 17629 7055 17663
rect 8769 17629 8803 17663
rect 9689 17629 9723 17663
rect 10057 17629 10091 17663
rect 10425 17629 10459 17663
rect 10701 17629 10735 17663
rect 11437 17629 11471 17663
rect 11897 17629 11931 17663
rect 13553 17629 13587 17663
rect 14841 17629 14875 17663
rect 16405 17629 16439 17663
rect 16589 17629 16623 17663
rect 19993 17629 20027 17663
rect 21373 17629 21407 17663
rect 23208 17629 23242 17663
rect 23305 17629 23339 17663
rect 23580 17629 23614 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 24593 17629 24627 17663
rect 25237 17629 25271 17663
rect 26893 17629 26927 17663
rect 27169 17629 27203 17663
rect 19395 17595 19429 17629
rect 1685 17561 1719 17595
rect 7205 17561 7239 17595
rect 12164 17561 12198 17595
rect 14197 17561 14231 17595
rect 15200 17561 15234 17595
rect 19625 17561 19659 17595
rect 23397 17561 23431 17595
rect 24777 17561 24811 17595
rect 25504 17561 25538 17595
rect 26709 17561 26743 17595
rect 27436 17561 27470 17595
rect 1885 17493 1919 17527
rect 2053 17493 2087 17527
rect 4629 17493 4663 17527
rect 5733 17493 5767 17527
rect 16313 17493 16347 17527
rect 17141 17493 17175 17527
rect 20177 17493 20211 17527
rect 21557 17493 21591 17527
rect 27077 17493 27111 17527
rect 2145 17289 2179 17323
rect 2789 17289 2823 17323
rect 3065 17289 3099 17323
rect 3341 17289 3375 17323
rect 5273 17289 5307 17323
rect 7665 17289 7699 17323
rect 12173 17289 12207 17323
rect 13829 17289 13863 17323
rect 14565 17289 14599 17323
rect 15393 17289 15427 17323
rect 21373 17289 21407 17323
rect 23213 17289 23247 17323
rect 23489 17289 23523 17323
rect 25513 17289 25547 17323
rect 27445 17289 27479 17323
rect 1961 17221 1995 17255
rect 2605 17221 2639 17255
rect 7941 17221 7975 17255
rect 22293 17221 22327 17255
rect 24602 17221 24636 17255
rect 26985 17221 27019 17255
rect 2881 17153 2915 17187
rect 3249 17153 3283 17187
rect 3801 17153 3835 17187
rect 5641 17153 5675 17187
rect 5917 17153 5951 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 7021 17153 7055 17187
rect 8125 17153 8159 17187
rect 8861 17153 8895 17187
rect 12357 17153 12391 17187
rect 13001 17153 13035 17187
rect 13277 17153 13311 17187
rect 13645 17153 13679 17187
rect 13737 17153 13771 17187
rect 14381 17153 14415 17187
rect 14657 17153 14691 17187
rect 15577 17153 15611 17187
rect 18061 17153 18095 17187
rect 18245 17153 18279 17187
rect 18788 17153 18822 17187
rect 20249 17153 20283 17187
rect 22017 17153 22051 17187
rect 23029 17153 23063 17187
rect 24869 17153 24903 17187
rect 25329 17153 25363 17187
rect 27169 17153 27203 17187
rect 27353 17153 27387 17187
rect 27629 17153 27663 17187
rect 8585 17085 8619 17119
rect 13093 17085 13127 17119
rect 13185 17085 13219 17119
rect 14197 17085 14231 17119
rect 18521 17085 18555 17119
rect 19993 17085 20027 17119
rect 22201 17085 22235 17119
rect 22845 17085 22879 17119
rect 1593 17017 1627 17051
rect 2237 17017 2271 17051
rect 5917 17017 5951 17051
rect 6469 17017 6503 17051
rect 8493 17017 8527 17051
rect 21833 17017 21867 17051
rect 1961 16949 1995 16983
rect 2605 16949 2639 16983
rect 7113 16949 7147 16983
rect 8677 16949 8711 16983
rect 13461 16949 13495 16983
rect 18429 16949 18463 16983
rect 19901 16949 19935 16983
rect 22201 16949 22235 16983
rect 8769 16745 8803 16779
rect 10149 16745 10183 16779
rect 11161 16745 11195 16779
rect 13185 16745 13219 16779
rect 16405 16745 16439 16779
rect 16865 16745 16899 16779
rect 18797 16745 18831 16779
rect 19441 16745 19475 16779
rect 20085 16745 20119 16779
rect 20545 16745 20579 16779
rect 22845 16745 22879 16779
rect 24041 16745 24075 16779
rect 25329 16745 25363 16779
rect 9413 16677 9447 16711
rect 11253 16677 11287 16711
rect 11713 16677 11747 16711
rect 18245 16677 18279 16711
rect 19257 16677 19291 16711
rect 23857 16677 23891 16711
rect 25145 16677 25179 16711
rect 5365 16609 5399 16643
rect 5641 16609 5675 16643
rect 9689 16609 9723 16643
rect 12265 16609 12299 16643
rect 16773 16609 16807 16643
rect 17785 16609 17819 16643
rect 21373 16609 21407 16643
rect 25881 16609 25915 16643
rect 3500 16542 3534 16576
rect 3801 16541 3835 16575
rect 4261 16541 4295 16575
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 5549 16541 5583 16575
rect 5917 16541 5951 16575
rect 7389 16541 7423 16575
rect 9597 16541 9631 16575
rect 9873 16541 9907 16575
rect 9965 16541 9999 16575
rect 11437 16541 11471 16575
rect 11529 16541 11563 16575
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 12633 16541 12667 16575
rect 14381 16541 14415 16575
rect 16589 16541 16623 16575
rect 17877 16541 17911 16575
rect 18429 16541 18463 16575
rect 18613 16541 18647 16575
rect 19901 16541 19935 16575
rect 21097 16541 21131 16575
rect 23024 16541 23058 16575
rect 23396 16541 23430 16575
rect 23489 16541 23523 16575
rect 27353 16541 27387 16575
rect 3893 16473 3927 16507
rect 4629 16473 4663 16507
rect 5457 16473 5491 16507
rect 7656 16473 7690 16507
rect 9045 16473 9079 16507
rect 10793 16473 10827 16507
rect 10977 16473 11011 16507
rect 12817 16473 12851 16507
rect 13001 16473 13035 16507
rect 16865 16473 16899 16507
rect 17417 16473 17451 16507
rect 17601 16473 17635 16507
rect 19625 16473 19659 16507
rect 19717 16473 19751 16507
rect 20729 16473 20763 16507
rect 21618 16473 21652 16507
rect 23121 16473 23155 16507
rect 23213 16473 23247 16507
rect 23581 16473 23615 16507
rect 24869 16473 24903 16507
rect 26148 16473 26182 16507
rect 3571 16405 3605 16439
rect 7205 16405 7239 16439
rect 9505 16405 9539 16439
rect 14197 16405 14231 16439
rect 18061 16405 18095 16439
rect 19425 16405 19459 16439
rect 20361 16405 20395 16439
rect 20524 16405 20558 16439
rect 21281 16405 21315 16439
rect 22753 16405 22787 16439
rect 27261 16405 27295 16439
rect 27537 16405 27571 16439
rect 3617 16201 3651 16235
rect 3985 16201 4019 16235
rect 7573 16201 7607 16235
rect 9321 16201 9355 16235
rect 10977 16201 11011 16235
rect 13093 16201 13127 16235
rect 15301 16201 15335 16235
rect 17049 16201 17083 16235
rect 20729 16201 20763 16235
rect 26433 16201 26467 16235
rect 1685 16133 1719 16167
rect 6469 16133 6503 16167
rect 8208 16133 8242 16167
rect 11713 16133 11747 16167
rect 13912 16133 13946 16167
rect 21985 16133 22019 16167
rect 22201 16133 22235 16167
rect 25973 16133 26007 16167
rect 27436 16133 27470 16167
rect 1501 16065 1535 16099
rect 2228 16065 2262 16099
rect 3801 16065 3835 16099
rect 4721 16065 4755 16099
rect 4813 16065 4847 16099
rect 5365 16065 5399 16099
rect 5641 16065 5675 16099
rect 5917 16065 5951 16099
rect 6193 16065 6227 16099
rect 7297 16065 7331 16099
rect 7389 16065 7423 16099
rect 9864 16065 9898 16099
rect 11897 16065 11931 16099
rect 13277 16065 13311 16099
rect 15209 16065 15243 16099
rect 16221 16065 16255 16099
rect 16405 16065 16439 16099
rect 18162 16065 18196 16099
rect 18429 16065 18463 16099
rect 20361 16065 20395 16099
rect 20545 16065 20579 16099
rect 21097 16065 21131 16099
rect 24501 16065 24535 16099
rect 24768 16065 24802 16099
rect 26157 16065 26191 16099
rect 26341 16065 26375 16099
rect 26617 16065 26651 16099
rect 27169 16065 27203 16099
rect 1961 15997 1995 16031
rect 3893 15997 3927 16031
rect 4261 15997 4295 16031
rect 4353 15997 4387 16031
rect 6929 15997 6963 16031
rect 7941 15997 7975 16031
rect 9597 15997 9631 16031
rect 13645 15997 13679 16031
rect 15577 15997 15611 16031
rect 15669 15997 15703 16031
rect 3341 15929 3375 15963
rect 6101 15929 6135 15963
rect 6745 15929 6779 15963
rect 7113 15929 7147 15963
rect 16129 15929 16163 15963
rect 4537 15861 4571 15895
rect 11529 15861 11563 15895
rect 15025 15861 15059 15895
rect 15393 15861 15427 15895
rect 15485 15861 15519 15895
rect 15945 15861 15979 15895
rect 16037 15861 16071 15895
rect 21005 15861 21039 15895
rect 21833 15861 21867 15895
rect 22017 15861 22051 15895
rect 25881 15861 25915 15895
rect 28549 15861 28583 15895
rect 3893 15657 3927 15691
rect 9781 15657 9815 15691
rect 10793 15657 10827 15691
rect 12449 15657 12483 15691
rect 14657 15657 14691 15691
rect 15761 15657 15795 15691
rect 16221 15657 16255 15691
rect 17601 15657 17635 15691
rect 17693 15657 17727 15691
rect 17785 15657 17819 15691
rect 23121 15657 23155 15691
rect 23949 15657 23983 15691
rect 24593 15657 24627 15691
rect 24777 15657 24811 15691
rect 27077 15657 27111 15691
rect 13093 15589 13127 15623
rect 15117 15589 15151 15623
rect 17325 15589 17359 15623
rect 22937 15589 22971 15623
rect 23765 15589 23799 15623
rect 3571 15521 3605 15555
rect 4813 15521 4847 15555
rect 6101 15521 6135 15555
rect 11069 15521 11103 15555
rect 13369 15521 13403 15555
rect 1777 15453 1811 15487
rect 1869 15453 1903 15487
rect 2053 15453 2087 15487
rect 2237 15453 2271 15487
rect 3468 15447 3502 15481
rect 4077 15453 4111 15487
rect 4261 15453 4295 15487
rect 4353 15453 4387 15487
rect 4537 15453 4571 15487
rect 4997 15453 5031 15487
rect 7665 15453 7699 15487
rect 8401 15453 8435 15487
rect 9413 15453 9447 15487
rect 9597 15453 9631 15487
rect 10977 15453 11011 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 14381 15453 14415 15487
rect 14841 15453 14875 15487
rect 15485 15453 15519 15487
rect 17877 15453 17911 15487
rect 18061 15453 18095 15487
rect 18521 15453 18555 15487
rect 18613 15453 18647 15487
rect 19257 15453 19291 15487
rect 21189 15453 21223 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 22753 15453 22787 15487
rect 24409 15453 24443 15487
rect 24961 15453 24995 15487
rect 28457 15453 28491 15487
rect 4169 15385 4203 15419
rect 11314 15385 11348 15419
rect 13829 15385 13863 15419
rect 14197 15385 14231 15419
rect 14565 15385 14599 15419
rect 15025 15385 15059 15419
rect 15301 15385 15335 15419
rect 15945 15385 15979 15419
rect 16037 15385 16071 15419
rect 18153 15385 18187 15419
rect 18337 15385 18371 15419
rect 19502 15385 19536 15419
rect 20729 15385 20763 15419
rect 20913 15385 20947 15419
rect 23305 15385 23339 15419
rect 24133 15385 24167 15419
rect 28190 15385 28224 15419
rect 1593 15317 1627 15351
rect 5181 15317 5215 15351
rect 5549 15317 5583 15351
rect 7481 15317 7515 15351
rect 8217 15317 8251 15351
rect 9229 15317 9263 15351
rect 12909 15317 12943 15351
rect 15577 15317 15611 15351
rect 15745 15317 15779 15351
rect 16237 15317 16271 15351
rect 16405 15317 16439 15351
rect 18797 15317 18831 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 22661 15317 22695 15351
rect 23095 15317 23129 15351
rect 23923 15317 23957 15351
rect 6101 15113 6135 15147
rect 7757 15113 7791 15147
rect 9597 15113 9631 15147
rect 11161 15113 11195 15147
rect 12449 15113 12483 15147
rect 14657 15113 14691 15147
rect 18061 15113 18095 15147
rect 24961 15113 24995 15147
rect 27445 15113 27479 15147
rect 1676 15045 1710 15079
rect 8392 15045 8426 15079
rect 12265 15045 12299 15079
rect 20897 15045 20931 15079
rect 21097 15045 21131 15079
rect 22170 15045 22204 15079
rect 25421 15045 25455 15079
rect 3065 14977 3099 15011
rect 3249 14977 3283 15011
rect 3341 14977 3375 15011
rect 4169 14977 4203 15011
rect 4445 14977 4479 15011
rect 4629 14977 4663 15011
rect 4721 14977 4755 15011
rect 4977 14977 5011 15011
rect 6653 14977 6687 15011
rect 10701 14977 10735 15011
rect 11345 14977 11379 15011
rect 12081 14977 12115 15011
rect 13001 14977 13035 15011
rect 14841 14977 14875 15011
rect 16313 14977 16347 15011
rect 16937 14977 16971 15011
rect 20177 14977 20211 15011
rect 20361 14977 20395 15011
rect 21925 14977 21959 15011
rect 23489 14977 23523 15011
rect 23756 14977 23790 15011
rect 26157 14977 26191 15011
rect 27261 14977 27295 15011
rect 1409 14909 1443 14943
rect 6377 14909 6411 14943
rect 8125 14909 8159 14943
rect 10057 14909 10091 14943
rect 16681 14909 16715 14943
rect 25605 14909 25639 14943
rect 26065 14909 26099 14943
rect 4445 14841 4479 14875
rect 9689 14841 9723 14875
rect 25053 14841 25087 14875
rect 25881 14841 25915 14875
rect 2789 14773 2823 14807
rect 2881 14773 2915 14807
rect 9505 14773 9539 14807
rect 10885 14773 10919 14807
rect 12817 14773 12851 14807
rect 16497 14773 16531 14807
rect 19993 14773 20027 14807
rect 20729 14773 20763 14807
rect 20913 14773 20947 14807
rect 23305 14773 23339 14807
rect 24869 14773 24903 14807
rect 26341 14773 26375 14807
rect 1869 14569 1903 14603
rect 3801 14569 3835 14603
rect 4813 14569 4847 14603
rect 5365 14569 5399 14603
rect 15761 14569 15795 14603
rect 17417 14569 17451 14603
rect 19993 14569 20027 14603
rect 23857 14569 23891 14603
rect 27629 14569 27663 14603
rect 23489 14501 23523 14535
rect 27537 14501 27571 14535
rect 4077 14433 4111 14467
rect 4169 14433 4203 14467
rect 8953 14433 8987 14467
rect 23581 14433 23615 14467
rect 2145 14365 2179 14399
rect 3985 14365 4019 14399
rect 4261 14365 4295 14399
rect 4813 14365 4847 14399
rect 4997 14365 5031 14399
rect 5273 14365 5307 14399
rect 7113 14365 7147 14399
rect 7380 14365 7414 14399
rect 9220 14365 9254 14399
rect 10609 14365 10643 14399
rect 10876 14365 10910 14399
rect 12173 14365 12207 14399
rect 12440 14365 12474 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15577 14365 15611 14399
rect 18061 14365 18095 14399
rect 18153 14365 18187 14399
rect 20453 14365 20487 14399
rect 20821 14365 20855 14399
rect 23673 14365 23707 14399
rect 24777 14365 24811 14399
rect 26810 14365 26844 14399
rect 27077 14365 27111 14399
rect 1961 14297 1995 14331
rect 2412 14297 2446 14331
rect 14657 14297 14691 14331
rect 15301 14297 15335 14331
rect 15485 14297 15519 14331
rect 17233 14297 17267 14331
rect 17433 14297 17467 14331
rect 17693 14297 17727 14331
rect 17877 14297 17911 14331
rect 19809 14297 19843 14331
rect 20269 14297 20303 14331
rect 21066 14297 21100 14331
rect 23121 14297 23155 14331
rect 27169 14297 27203 14331
rect 3525 14229 3559 14263
rect 8493 14229 8527 14263
rect 10333 14229 10367 14263
rect 11989 14229 12023 14263
rect 13553 14229 13587 14263
rect 15117 14229 15151 14263
rect 17601 14229 17635 14263
rect 18337 14229 18371 14263
rect 20009 14229 20043 14263
rect 20177 14229 20211 14263
rect 20637 14229 20671 14263
rect 22201 14229 22235 14263
rect 24869 14229 24903 14263
rect 25697 14229 25731 14263
rect 1593 14025 1627 14059
rect 2973 14025 3007 14059
rect 3525 14025 3559 14059
rect 4445 14025 4479 14059
rect 10425 14025 10459 14059
rect 12173 14025 12207 14059
rect 14105 14025 14139 14059
rect 16129 14025 16163 14059
rect 17325 14025 17359 14059
rect 18153 14025 18187 14059
rect 19717 14025 19751 14059
rect 20453 14025 20487 14059
rect 20821 14025 20855 14059
rect 23949 14025 23983 14059
rect 2697 13957 2731 13991
rect 2881 13957 2915 13991
rect 4597 13957 4631 13991
rect 4813 13957 4847 13991
rect 7573 13957 7607 13991
rect 8953 13957 8987 13991
rect 10793 13957 10827 13991
rect 14381 13957 14415 13991
rect 14473 13957 14507 13991
rect 18582 13957 18616 13991
rect 22293 13957 22327 13991
rect 22063 13923 22097 13957
rect 1409 13889 1443 13923
rect 3065 13889 3099 13923
rect 3249 13889 3283 13923
rect 3617 13889 3651 13923
rect 10609 13889 10643 13923
rect 11989 13889 12023 13923
rect 13645 13889 13679 13923
rect 13737 13889 13771 13923
rect 13921 13889 13955 13923
rect 14013 13889 14047 13923
rect 14289 13889 14323 13923
rect 14657 13889 14691 13923
rect 15016 13889 15050 13923
rect 17417 13889 17451 13923
rect 17785 13889 17819 13923
rect 18245 13889 18279 13923
rect 20177 13889 20211 13923
rect 20545 13889 20579 13923
rect 20637 13889 20671 13923
rect 22569 13889 22603 13923
rect 23765 13889 23799 13923
rect 28282 13889 28316 13923
rect 28549 13889 28583 13923
rect 14749 13821 14783 13855
rect 17141 13821 17175 13855
rect 18337 13821 18371 13855
rect 25697 13821 25731 13855
rect 7941 13753 7975 13787
rect 9229 13753 9263 13787
rect 13461 13753 13495 13787
rect 16957 13753 16991 13787
rect 20085 13753 20119 13787
rect 21925 13753 21959 13787
rect 25973 13753 26007 13787
rect 27169 13753 27203 13787
rect 4629 13685 4663 13719
rect 8033 13685 8067 13719
rect 9413 13685 9447 13719
rect 16681 13685 16715 13719
rect 17049 13685 17083 13719
rect 17509 13685 17543 13719
rect 17877 13685 17911 13719
rect 17969 13685 18003 13719
rect 19809 13685 19843 13719
rect 20269 13685 20303 13719
rect 22109 13685 22143 13719
rect 22385 13685 22419 13719
rect 26157 13685 26191 13719
rect 2145 13481 2179 13515
rect 4721 13481 4755 13515
rect 6193 13481 6227 13515
rect 8769 13481 8803 13515
rect 13645 13481 13679 13515
rect 15025 13481 15059 13515
rect 16405 13481 16439 13515
rect 16681 13481 16715 13515
rect 17325 13481 17359 13515
rect 19901 13481 19935 13515
rect 20085 13481 20119 13515
rect 20729 13481 20763 13515
rect 20821 13481 20855 13515
rect 22017 13481 22051 13515
rect 24041 13481 24075 13515
rect 28089 13481 28123 13515
rect 4169 13413 4203 13447
rect 11069 13413 11103 13447
rect 21925 13413 21959 13447
rect 23949 13413 23983 13447
rect 27629 13413 27663 13447
rect 4813 13345 4847 13379
rect 7389 13345 7423 13379
rect 12265 13345 12299 13379
rect 19257 13345 19291 13379
rect 27261 13345 27295 13379
rect 27353 13345 27387 13379
rect 27813 13345 27847 13379
rect 2329 13277 2363 13311
rect 2605 13277 2639 13311
rect 2789 13277 2823 13311
rect 3893 13277 3927 13311
rect 3985 13277 4019 13311
rect 4261 13277 4295 13311
rect 4445 13277 4479 13311
rect 6837 13277 6871 13311
rect 8953 13277 8987 13311
rect 9046 13277 9080 13311
rect 9321 13277 9355 13311
rect 9459 13277 9493 13311
rect 9689 13277 9723 13311
rect 11345 13277 11379 13311
rect 11438 13277 11472 13311
rect 11621 13277 11655 13311
rect 11713 13277 11747 13311
rect 11851 13277 11885 13311
rect 12521 13277 12555 13311
rect 14565 13277 14599 13311
rect 15209 13277 15243 13311
rect 16589 13277 16623 13311
rect 16681 13277 16715 13311
rect 18797 13277 18831 13311
rect 18981 13277 19015 13311
rect 19625 13277 19659 13311
rect 19809 13277 19843 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 20913 13277 20947 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 22109 13277 22143 13311
rect 25522 13277 25556 13311
rect 25789 13277 25823 13311
rect 27905 13277 27939 13311
rect 2513 13209 2547 13243
rect 4169 13209 4203 13243
rect 5058 13209 5092 13243
rect 7656 13209 7690 13243
rect 9229 13209 9263 13243
rect 9934 13209 9968 13243
rect 14749 13209 14783 13243
rect 16865 13209 16899 13243
rect 17509 13209 17543 13243
rect 19441 13209 19475 13243
rect 19717 13209 19751 13243
rect 20085 13209 20119 13243
rect 22376 13209 22410 13243
rect 23581 13209 23615 13243
rect 26994 13209 27028 13243
rect 2605 13141 2639 13175
rect 4537 13141 4571 13175
rect 6653 13141 6687 13175
rect 9597 13141 9631 13175
rect 11989 13141 12023 13175
rect 14933 13141 14967 13175
rect 17141 13141 17175 13175
rect 17309 13141 17343 13175
rect 18613 13141 18647 13175
rect 23489 13141 23523 13175
rect 24409 13141 24443 13175
rect 25881 13141 25915 13175
rect 2789 12937 2823 12971
rect 3065 12937 3099 12971
rect 5181 12937 5215 12971
rect 9781 12937 9815 12971
rect 11989 12937 12023 12971
rect 12357 12937 12391 12971
rect 15025 12937 15059 12971
rect 19257 12937 19291 12971
rect 20269 12937 20303 12971
rect 20913 12937 20947 12971
rect 26249 12937 26283 12971
rect 28549 12937 28583 12971
rect 3862 12869 3896 12903
rect 6633 12869 6667 12903
rect 9229 12869 9263 12903
rect 12449 12869 12483 12903
rect 15362 12869 15396 12903
rect 18122 12869 18156 12903
rect 22109 12869 22143 12903
rect 23029 12869 23063 12903
rect 25697 12869 25731 12903
rect 1409 12801 1443 12835
rect 1676 12801 1710 12835
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 3525 12801 3559 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 8033 12801 8067 12835
rect 8953 12801 8987 12835
rect 9137 12801 9171 12835
rect 9321 12801 9355 12835
rect 9597 12801 9631 12835
rect 11529 12801 11563 12835
rect 12173 12801 12207 12835
rect 13001 12801 13035 12835
rect 13257 12801 13291 12835
rect 14841 12801 14875 12835
rect 15117 12801 15151 12835
rect 17049 12801 17083 12835
rect 17141 12801 17175 12835
rect 17279 12801 17313 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 17877 12801 17911 12835
rect 21008 12801 21042 12835
rect 21097 12801 21131 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 22319 12801 22353 12835
rect 24786 12801 24820 12835
rect 25053 12801 25087 12835
rect 26065 12801 26099 12835
rect 27169 12801 27203 12835
rect 27436 12801 27470 12835
rect 3617 12733 3651 12767
rect 6377 12733 6411 12767
rect 12081 12733 12115 12767
rect 20729 12733 20763 12767
rect 22477 12733 22511 12767
rect 23489 12733 23523 12767
rect 4997 12665 5031 12699
rect 7849 12665 7883 12699
rect 11805 12665 11839 12699
rect 16497 12665 16531 12699
rect 17785 12665 17819 12699
rect 20545 12665 20579 12699
rect 20637 12665 20671 12699
rect 23397 12665 23431 12699
rect 23673 12665 23707 12699
rect 25329 12665 25363 12699
rect 6193 12597 6227 12631
rect 7757 12597 7791 12631
rect 9505 12597 9539 12631
rect 12265 12597 12299 12631
rect 14381 12597 14415 12631
rect 16681 12597 16715 12631
rect 16957 12597 16991 12631
rect 21281 12597 21315 12631
rect 21833 12597 21867 12631
rect 25237 12597 25271 12631
rect 1869 12393 1903 12427
rect 2789 12393 2823 12427
rect 13001 12393 13035 12427
rect 15485 12393 15519 12427
rect 15669 12393 15703 12427
rect 16129 12393 16163 12427
rect 16313 12393 16347 12427
rect 17417 12393 17451 12427
rect 18245 12393 18279 12427
rect 19625 12393 19659 12427
rect 23857 12393 23891 12427
rect 27537 12393 27571 12427
rect 1593 12325 1627 12359
rect 7757 12325 7791 12359
rect 12541 12325 12575 12359
rect 18153 12325 18187 12359
rect 19993 12325 20027 12359
rect 21281 12325 21315 12359
rect 6377 12257 6411 12291
rect 12173 12257 12207 12291
rect 12633 12257 12667 12291
rect 17785 12257 17819 12291
rect 20085 12257 20119 12291
rect 20913 12257 20947 12291
rect 1409 12189 1443 12223
rect 2053 12189 2087 12223
rect 2329 12189 2363 12223
rect 3801 12189 3835 12223
rect 5549 12189 5583 12223
rect 6101 12189 6135 12223
rect 12817 12189 12851 12223
rect 14381 12189 14415 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 17233 12189 17267 12223
rect 18061 12189 18095 12223
rect 18337 12189 18371 12223
rect 18521 12189 18555 12223
rect 18613 12189 18647 12223
rect 18797 12189 18831 12223
rect 19901 12189 19935 12223
rect 20361 12189 20395 12223
rect 21097 12189 21131 12223
rect 23673 12189 23707 12223
rect 25053 12189 25087 12223
rect 26709 12189 26743 12223
rect 27353 12189 27387 12223
rect 2513 12121 2547 12155
rect 6622 12121 6656 12155
rect 15301 12121 15335 12155
rect 15945 12121 15979 12155
rect 17049 12121 17083 12155
rect 26442 12121 26476 12155
rect 2237 12053 2271 12087
rect 6285 12053 6319 12087
rect 14197 12053 14231 12087
rect 15501 12053 15535 12087
rect 16145 12053 16179 12087
rect 18981 12053 19015 12087
rect 20269 12053 20303 12087
rect 25237 12053 25271 12087
rect 25329 12053 25363 12087
rect 3801 11849 3835 11883
rect 4353 11849 4387 11883
rect 6377 11849 6411 11883
rect 9597 11849 9631 11883
rect 12173 11849 12207 11883
rect 19273 11849 19307 11883
rect 19441 11849 19475 11883
rect 6837 11781 6871 11815
rect 9934 11781 9968 11815
rect 11713 11781 11747 11815
rect 19073 11781 19107 11815
rect 21281 11781 21315 11815
rect 22569 11781 22603 11815
rect 23055 11781 23089 11815
rect 24869 11781 24903 11815
rect 2237 11713 2271 11747
rect 3985 11713 4019 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 4445 11713 4479 11747
rect 4721 11713 4755 11747
rect 5641 11713 5675 11747
rect 8033 11713 8067 11747
rect 9413 11713 9447 11747
rect 9689 11713 9723 11747
rect 12817 11713 12851 11747
rect 20177 11713 20211 11747
rect 21005 11713 21039 11747
rect 21098 11713 21132 11747
rect 21373 11713 21407 11747
rect 21470 11713 21504 11747
rect 21833 11713 21867 11747
rect 21926 11713 21960 11747
rect 22109 11713 22143 11747
rect 22201 11713 22235 11747
rect 22298 11713 22332 11747
rect 22753 11713 22787 11747
rect 22845 11713 22879 11747
rect 22937 11713 22971 11747
rect 23213 11713 23247 11747
rect 25421 11713 25455 11747
rect 27436 11713 27470 11747
rect 2329 11645 2363 11679
rect 5273 11645 5307 11679
rect 8125 11645 8159 11679
rect 8585 11645 8619 11679
rect 8769 11645 8803 11679
rect 9229 11645 9263 11679
rect 25329 11645 25363 11679
rect 27169 11645 27203 11679
rect 2697 11577 2731 11611
rect 6561 11577 6595 11611
rect 8309 11577 8343 11611
rect 9045 11577 9079 11611
rect 11069 11577 11103 11611
rect 11989 11577 12023 11611
rect 21649 11577 21683 11611
rect 25145 11577 25179 11611
rect 1961 11509 1995 11543
rect 2513 11509 2547 11543
rect 5825 11509 5859 11543
rect 7849 11509 7883 11543
rect 13001 11509 13035 11543
rect 19257 11509 19291 11543
rect 20361 11509 20395 11543
rect 22477 11509 22511 11543
rect 25605 11509 25639 11543
rect 28549 11509 28583 11543
rect 5365 11305 5399 11339
rect 6837 11305 6871 11339
rect 10057 11305 10091 11339
rect 14289 11305 14323 11339
rect 14749 11305 14783 11339
rect 27353 11305 27387 11339
rect 27445 11305 27479 11339
rect 5181 11237 5215 11271
rect 8769 11237 8803 11271
rect 10793 11237 10827 11271
rect 14105 11237 14139 11271
rect 18521 11237 18555 11271
rect 23581 11237 23615 11271
rect 24777 11237 24811 11271
rect 27169 11237 27203 11271
rect 9045 11169 9079 11203
rect 9873 11169 9907 11203
rect 13645 11169 13679 11203
rect 23121 11169 23155 11203
rect 23489 11169 23523 11203
rect 3249 11101 3283 11135
rect 3617 11101 3651 11135
rect 3801 11101 3835 11135
rect 5457 11101 5491 11135
rect 5724 11101 5758 11135
rect 7297 11101 7331 11135
rect 7389 11101 7423 11135
rect 7656 11101 7690 11135
rect 9203 11101 9237 11135
rect 9413 11101 9447 11135
rect 9505 11101 9539 11135
rect 9689 11101 9723 11135
rect 10057 11101 10091 11135
rect 10977 11101 11011 11135
rect 11069 11101 11103 11135
rect 13378 11101 13412 11135
rect 15945 11101 15979 11135
rect 17877 11101 17911 11135
rect 18061 11101 18095 11135
rect 18337 11101 18371 11135
rect 19257 11101 19291 11135
rect 19513 11101 19547 11135
rect 20729 11101 20763 11135
rect 20985 11101 21019 11135
rect 23305 11101 23339 11135
rect 23719 11101 23753 11135
rect 23949 11101 23983 11135
rect 24132 11101 24166 11135
rect 24225 11101 24259 11135
rect 25890 11101 25924 11135
rect 26157 11101 26191 11135
rect 27629 11101 27663 11135
rect 3157 11033 3191 11067
rect 3433 11033 3467 11067
rect 4905 11033 4939 11067
rect 9321 11033 9355 11067
rect 9781 11033 9815 11067
rect 14273 11033 14307 11067
rect 14473 11033 14507 11067
rect 14733 11033 14767 11067
rect 14933 11033 14967 11067
rect 15485 11033 15519 11067
rect 15669 11033 15703 11067
rect 16212 11033 16246 11067
rect 23857 11033 23891 11067
rect 26893 11033 26927 11067
rect 1869 10965 1903 10999
rect 3985 10965 4019 10999
rect 7113 10965 7147 10999
rect 10241 10965 10275 10999
rect 12265 10965 12299 10999
rect 14565 10965 14599 10999
rect 15853 10965 15887 10999
rect 17325 10965 17359 10999
rect 18245 10965 18279 10999
rect 20637 10965 20671 10999
rect 22109 10965 22143 10999
rect 2973 10761 3007 10795
rect 6009 10761 6043 10795
rect 9873 10761 9907 10795
rect 10517 10761 10551 10795
rect 10701 10761 10735 10795
rect 12265 10761 12299 10795
rect 12909 10761 12943 10795
rect 14473 10761 14507 10795
rect 15945 10761 15979 10795
rect 16221 10761 16255 10795
rect 17049 10761 17083 10795
rect 17693 10761 17727 10795
rect 18337 10761 18371 10795
rect 18781 10761 18815 10795
rect 20361 10761 20395 10795
rect 22109 10761 22143 10795
rect 22753 10761 22787 10795
rect 27445 10761 27479 10795
rect 4086 10693 4120 10727
rect 5672 10693 5706 10727
rect 7012 10693 7046 10727
rect 8835 10693 8869 10727
rect 8953 10693 8987 10727
rect 11161 10693 11195 10727
rect 11805 10693 11839 10727
rect 14810 10693 14844 10727
rect 18981 10693 19015 10727
rect 20913 10693 20947 10727
rect 21097 10693 21131 10727
rect 23673 10693 23707 10727
rect 24409 10693 24443 10727
rect 25329 10693 25363 10727
rect 26985 10693 27019 10727
rect 1501 10625 1535 10659
rect 2421 10625 2455 10659
rect 2605 10625 2639 10659
rect 4353 10625 4387 10659
rect 6193 10625 6227 10659
rect 6745 10625 6779 10659
rect 8677 10625 8711 10659
rect 9045 10625 9079 10659
rect 9137 10625 9171 10659
rect 10241 10625 10275 10659
rect 10609 10625 10643 10659
rect 10885 10625 10919 10659
rect 11529 10625 11563 10659
rect 11677 10625 11711 10659
rect 11897 10625 11931 10659
rect 11994 10625 12028 10659
rect 12449 10625 12483 10659
rect 12725 10625 12759 10659
rect 13093 10625 13127 10659
rect 13277 10625 13311 10659
rect 13369 10625 13403 10659
rect 14289 10625 14323 10659
rect 16037 10625 16071 10659
rect 17509 10625 17543 10659
rect 17722 10625 17756 10659
rect 19993 10625 20027 10659
rect 20177 10625 20211 10659
rect 22845 10625 22879 10659
rect 23484 10625 23518 10659
rect 23581 10625 23615 10659
rect 23801 10625 23835 10659
rect 23949 10625 23983 10659
rect 24041 10625 24075 10659
rect 24225 10625 24259 10659
rect 24317 10625 24351 10659
rect 24527 10625 24561 10659
rect 26065 10625 26099 10659
rect 5917 10557 5951 10591
rect 10149 10557 10183 10591
rect 11069 10557 11103 10591
rect 12633 10557 12667 10591
rect 14565 10557 14599 10591
rect 17877 10557 17911 10591
rect 24685 10557 24719 10591
rect 25789 10557 25823 10591
rect 12173 10489 12207 10523
rect 17325 10489 17359 10523
rect 18153 10489 18187 10523
rect 23305 10489 23339 10523
rect 25697 10489 25731 10523
rect 27261 10489 27295 10523
rect 1593 10421 1627 10455
rect 4537 10421 4571 10455
rect 8125 10421 8159 10455
rect 9321 10421 9355 10455
rect 10333 10421 10367 10455
rect 10885 10421 10919 10455
rect 12449 10421 12483 10455
rect 13553 10421 13587 10455
rect 17417 10421 17451 10455
rect 18613 10421 18647 10455
rect 18797 10421 18831 10455
rect 21281 10421 21315 10455
rect 22385 10421 22419 10455
rect 22477 10421 22511 10455
rect 22569 10421 22603 10455
rect 25881 10421 25915 10455
rect 5181 10217 5215 10251
rect 5733 10217 5767 10251
rect 7573 10217 7607 10251
rect 9229 10217 9263 10251
rect 9505 10217 9539 10251
rect 10793 10217 10827 10251
rect 10977 10217 11011 10251
rect 14657 10217 14691 10251
rect 15485 10217 15519 10251
rect 15761 10217 15795 10251
rect 20453 10217 20487 10251
rect 20637 10217 20671 10251
rect 22201 10217 22235 10251
rect 22385 10217 22419 10251
rect 24409 10217 24443 10251
rect 28549 10217 28583 10251
rect 2329 10149 2363 10183
rect 5641 10149 5675 10183
rect 5825 10149 5859 10183
rect 7481 10149 7515 10183
rect 11989 10149 12023 10183
rect 14473 10149 14507 10183
rect 23581 10149 23615 10183
rect 12173 10081 12207 10115
rect 16681 10081 16715 10115
rect 25605 10081 25639 10115
rect 27169 10081 27203 10115
rect 1593 10013 1627 10047
rect 1869 10013 1903 10047
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 3065 10013 3099 10047
rect 3157 10013 3191 10047
rect 3801 10013 3835 10047
rect 6009 10013 6043 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 12265 10013 12299 10047
rect 14197 10013 14231 10047
rect 15853 10013 15887 10047
rect 15945 10013 15979 10047
rect 16221 10013 16255 10047
rect 17233 10013 17267 10047
rect 20729 10013 20763 10047
rect 22845 10013 22879 10047
rect 23029 10013 23063 10047
rect 23305 10013 23339 10047
rect 23673 10013 23707 10047
rect 23765 10013 23799 10047
rect 23857 10013 23891 10047
rect 24041 10013 24075 10047
rect 24593 10013 24627 10047
rect 24895 10013 24929 10047
rect 25053 10013 25087 10047
rect 25872 10013 25906 10047
rect 2697 9945 2731 9979
rect 2881 9945 2915 9979
rect 4046 9945 4080 9979
rect 5273 9945 5307 9979
rect 7113 9945 7147 9979
rect 9045 9945 9079 9979
rect 10609 9945 10643 9979
rect 11713 9945 11747 9979
rect 16865 9945 16899 9979
rect 19441 9945 19475 9979
rect 19625 9945 19659 9979
rect 20269 9945 20303 9979
rect 20996 9945 21030 9979
rect 22569 9945 22603 9979
rect 23213 9945 23247 9979
rect 24685 9945 24719 9979
rect 24777 9945 24811 9979
rect 27436 9945 27470 9979
rect 2053 9877 2087 9911
rect 3341 9877 3375 9911
rect 10809 9877 10843 9911
rect 12449 9877 12483 9911
rect 16129 9877 16163 9911
rect 17049 9877 17083 9911
rect 19257 9877 19291 9911
rect 20469 9877 20503 9911
rect 22109 9877 22143 9911
rect 22359 9877 22393 9911
rect 26985 9877 27019 9911
rect 10609 9673 10643 9707
rect 14197 9673 14231 9707
rect 14933 9673 14967 9707
rect 18061 9673 18095 9707
rect 21097 9673 21131 9707
rect 21189 9673 21223 9707
rect 22201 9673 22235 9707
rect 23029 9673 23063 9707
rect 27537 9673 27571 9707
rect 5080 9605 5114 9639
rect 10333 9605 10367 9639
rect 15285 9605 15319 9639
rect 15485 9605 15519 9639
rect 16497 9605 16531 9639
rect 16948 9605 16982 9639
rect 21833 9605 21867 9639
rect 22033 9605 22067 9639
rect 24593 9605 24627 9639
rect 26985 9605 27019 9639
rect 1409 9537 1443 9571
rect 1593 9537 1627 9571
rect 1685 9537 1719 9571
rect 1869 9537 1903 9571
rect 2237 9537 2271 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 3709 9537 3743 9571
rect 4813 9537 4847 9571
rect 6745 9537 6779 9571
rect 8125 9537 8159 9571
rect 9965 9537 9999 9571
rect 10058 9537 10092 9571
rect 10241 9537 10275 9571
rect 10471 9537 10505 9571
rect 11529 9537 11563 9571
rect 12817 9537 12851 9571
rect 13073 9537 13107 9571
rect 15025 9537 15059 9571
rect 16037 9537 16071 9571
rect 16129 9537 16163 9571
rect 16313 9537 16347 9571
rect 19358 9537 19392 9571
rect 19973 9537 20007 9571
rect 21373 9537 21407 9571
rect 22937 9537 22971 9571
rect 27721 9537 27755 9571
rect 12081 9469 12115 9503
rect 14565 9469 14599 9503
rect 16681 9469 16715 9503
rect 19625 9469 19659 9503
rect 19717 9469 19751 9503
rect 27445 9469 27479 9503
rect 2421 9401 2455 9435
rect 3893 9401 3927 9435
rect 6193 9401 6227 9435
rect 11713 9401 11747 9435
rect 12357 9401 12391 9435
rect 18245 9401 18279 9435
rect 27261 9401 27295 9435
rect 1961 9333 1995 9367
rect 2605 9333 2639 9367
rect 2881 9333 2915 9367
rect 6561 9333 6595 9367
rect 7941 9333 7975 9367
rect 12541 9333 12575 9367
rect 14289 9333 14323 9367
rect 14657 9333 14691 9367
rect 14749 9333 14783 9367
rect 15117 9333 15151 9367
rect 15301 9333 15335 9367
rect 15853 9333 15887 9367
rect 22017 9333 22051 9367
rect 24685 9333 24719 9367
rect 5733 9129 5767 9163
rect 7297 9129 7331 9163
rect 8769 9129 8803 9163
rect 9597 9129 9631 9163
rect 9781 9129 9815 9163
rect 10609 9129 10643 9163
rect 10885 9129 10919 9163
rect 12909 9129 12943 9163
rect 13369 9129 13403 9163
rect 15209 9129 15243 9163
rect 15669 9129 15703 9163
rect 15853 9129 15887 9163
rect 16129 9129 16163 9163
rect 16957 9129 16991 9163
rect 17141 9129 17175 9163
rect 18981 9129 19015 9163
rect 22845 9129 22879 9163
rect 23029 9129 23063 9163
rect 23581 9129 23615 9163
rect 23765 9129 23799 9163
rect 25789 9129 25823 9163
rect 28273 9129 28307 9163
rect 13553 9061 13587 9095
rect 15393 9061 15427 9095
rect 17969 9061 18003 9095
rect 18705 9061 18739 9095
rect 25973 9061 26007 9095
rect 5917 8993 5951 9027
rect 9965 8993 9999 9027
rect 13185 8993 13219 9027
rect 18153 8993 18187 9027
rect 26893 8993 26927 9027
rect 1501 8925 1535 8959
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 3801 8925 3835 8959
rect 5365 8925 5399 8959
rect 6184 8925 6218 8959
rect 7389 8925 7423 8959
rect 7656 8925 7690 8959
rect 10103 8925 10137 8959
rect 10216 8925 10250 8959
rect 10425 8925 10459 8959
rect 12285 8925 12319 8959
rect 12541 8925 12575 8959
rect 12725 8925 12759 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 17693 8925 17727 8959
rect 18521 8925 18555 8959
rect 18797 8925 18831 8959
rect 20821 8925 20855 8959
rect 21005 8925 21039 8959
rect 21373 8925 21407 8959
rect 24041 8925 24075 8959
rect 24409 8925 24443 8959
rect 26617 8925 26651 8959
rect 4046 8857 4080 8891
rect 5549 8857 5583 8891
rect 9413 8857 9447 8891
rect 9629 8857 9663 8891
rect 10333 8857 10367 8891
rect 10701 8857 10735 8891
rect 10901 8857 10935 8891
rect 13093 8857 13127 8891
rect 15025 8857 15059 8891
rect 15241 8857 15275 8891
rect 15485 8857 15519 8891
rect 15685 8857 15719 8891
rect 16313 8857 16347 8891
rect 16773 8857 16807 8891
rect 20637 8857 20671 8891
rect 22661 8857 22695 8891
rect 23397 8857 23431 8891
rect 24654 8857 24688 8891
rect 26341 8857 26375 8891
rect 27138 8857 27172 8891
rect 3157 8789 3191 8823
rect 5181 8789 5215 8823
rect 11069 8789 11103 8823
rect 11161 8789 11195 8823
rect 14105 8789 14139 8823
rect 15945 8789 15979 8823
rect 16113 8789 16147 8823
rect 16973 8789 17007 8823
rect 21557 8789 21591 8823
rect 22861 8789 22895 8823
rect 23607 8789 23641 8823
rect 24225 8789 24259 8823
rect 25881 8789 25915 8823
rect 26801 8789 26835 8823
rect 1593 8585 1627 8619
rect 2881 8585 2915 8619
rect 6837 8585 6871 8619
rect 8033 8585 8067 8619
rect 10901 8585 10935 8619
rect 14657 8585 14691 8619
rect 17141 8585 17175 8619
rect 18061 8585 18095 8619
rect 20611 8585 20645 8619
rect 21205 8585 21239 8619
rect 21373 8585 21407 8619
rect 23213 8585 23247 8619
rect 23305 8585 23339 8619
rect 24409 8585 24443 8619
rect 25329 8585 25363 8619
rect 26985 8585 27019 8619
rect 4169 8517 4203 8551
rect 7849 8517 7883 8551
rect 8309 8517 8343 8551
rect 8852 8517 8886 8551
rect 10701 8517 10735 8551
rect 11897 8517 11931 8551
rect 14289 8517 14323 8551
rect 15853 8517 15887 8551
rect 16069 8517 16103 8551
rect 16773 8517 16807 8551
rect 16973 8517 17007 8551
rect 17785 8517 17819 8551
rect 18213 8517 18247 8551
rect 18429 8517 18463 8551
rect 20821 8517 20855 8551
rect 21031 8517 21065 8551
rect 23457 8517 23491 8551
rect 23673 8517 23707 8551
rect 23765 8517 23799 8551
rect 23949 8517 23983 8551
rect 25666 8517 25700 8551
rect 27445 8517 27479 8551
rect 14519 8483 14553 8517
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1869 8449 1903 8483
rect 1961 8449 1995 8483
rect 5089 8449 5123 8483
rect 5917 8449 5951 8483
rect 7665 8449 7699 8483
rect 8125 8449 8159 8483
rect 11529 8449 11563 8483
rect 11677 8449 11711 8483
rect 11805 8449 11839 8483
rect 11994 8449 12028 8483
rect 17601 8449 17635 8483
rect 19809 8449 19843 8483
rect 22100 8449 22134 8483
rect 24869 8449 24903 8483
rect 25145 8449 25179 8483
rect 4813 8381 4847 8415
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 6377 8381 6411 8415
rect 8493 8381 8527 8415
rect 8585 8381 8619 8415
rect 21833 8381 21867 8415
rect 25421 8381 25455 8415
rect 5457 8313 5491 8347
rect 6653 8313 6687 8347
rect 11069 8313 11103 8347
rect 12173 8313 12207 8347
rect 20453 8313 20487 8347
rect 24593 8313 24627 8347
rect 27077 8313 27111 8347
rect 5733 8245 5767 8279
rect 9965 8245 9999 8279
rect 10885 8245 10919 8279
rect 14473 8245 14507 8279
rect 16037 8245 16071 8279
rect 16221 8245 16255 8279
rect 16957 8245 16991 8279
rect 18245 8245 18279 8279
rect 19993 8245 20027 8279
rect 20637 8245 20671 8279
rect 21189 8245 21223 8279
rect 23489 8245 23523 8279
rect 24133 8245 24167 8279
rect 26801 8245 26835 8279
rect 3341 8041 3375 8075
rect 8953 8041 8987 8075
rect 12265 8041 12299 8075
rect 12541 8041 12575 8075
rect 15853 8041 15887 8075
rect 16129 8041 16163 8075
rect 16313 8041 16347 8075
rect 19441 8041 19475 8075
rect 19625 8041 19659 8075
rect 21097 8041 21131 8075
rect 22477 8041 22511 8075
rect 22661 8041 22695 8075
rect 24225 8041 24259 8075
rect 4353 7973 4387 8007
rect 5917 7973 5951 8007
rect 6377 7973 6411 8007
rect 10333 7973 10367 8007
rect 12449 7973 12483 8007
rect 12817 7973 12851 8007
rect 17693 7973 17727 8007
rect 4537 7905 4571 7939
rect 6469 7905 6503 7939
rect 1593 7837 1627 7871
rect 1777 7837 1811 7871
rect 1869 7837 1903 7871
rect 2329 7837 2363 7871
rect 2513 7837 2547 7871
rect 2605 7837 2639 7871
rect 2789 7837 2823 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 6561 7837 6595 7871
rect 9137 7837 9171 7871
rect 10057 7837 10091 7871
rect 10793 7837 10827 7871
rect 11529 7837 11563 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 13277 7837 13311 7871
rect 14105 7837 14139 7871
rect 16221 7837 16255 7871
rect 16589 7837 16623 7871
rect 16773 7837 16807 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17325 7837 17359 7871
rect 19073 7837 19107 7871
rect 19717 7837 19751 7871
rect 19984 7837 20018 7871
rect 21373 7837 21407 7871
rect 22845 7837 22879 7871
rect 26801 7837 26835 7871
rect 3249 7769 3283 7803
rect 3985 7769 4019 7803
rect 4804 7769 4838 7803
rect 6009 7769 6043 7803
rect 12081 7769 12115 7803
rect 12281 7769 12315 7803
rect 14350 7769 14384 7803
rect 18806 7769 18840 7803
rect 19257 7769 19291 7803
rect 19457 7769 19491 7803
rect 21557 7769 21591 7803
rect 22293 7769 22327 7803
rect 23112 7769 23146 7803
rect 4445 7701 4479 7735
rect 6745 7701 6779 7735
rect 10517 7701 10551 7735
rect 10701 7701 10735 7735
rect 11713 7701 11747 7735
rect 13185 7701 13219 7735
rect 15485 7701 15519 7735
rect 16497 7701 16531 7735
rect 17509 7701 17543 7735
rect 21189 7701 21223 7735
rect 22493 7701 22527 7735
rect 26985 7701 27019 7735
rect 3433 7497 3467 7531
rect 4905 7497 4939 7531
rect 11345 7497 11379 7531
rect 12909 7497 12943 7531
rect 13093 7497 13127 7531
rect 14381 7497 14415 7531
rect 15853 7497 15887 7531
rect 16313 7497 16347 7531
rect 18061 7497 18095 7531
rect 18705 7497 18739 7531
rect 19901 7497 19935 7531
rect 23305 7497 23339 7531
rect 24317 7497 24351 7531
rect 25789 7497 25823 7531
rect 26801 7497 26835 7531
rect 28365 7497 28399 7531
rect 6644 7429 6678 7463
rect 13261 7429 13295 7463
rect 13461 7429 13495 7463
rect 13737 7429 13771 7463
rect 14718 7429 14752 7463
rect 15945 7429 15979 7463
rect 16161 7429 16195 7463
rect 16957 7429 16991 7463
rect 19441 7429 19475 7463
rect 23857 7429 23891 7463
rect 24654 7429 24688 7463
rect 26341 7429 26375 7463
rect 27230 7429 27264 7463
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 2329 7361 2363 7395
rect 2881 7361 2915 7395
rect 4557 7361 4591 7395
rect 5089 7361 5123 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 8309 7361 8343 7395
rect 8585 7361 8619 7395
rect 10232 7361 10266 7395
rect 11529 7361 11563 7395
rect 11785 7361 11819 7395
rect 13553 7361 13587 7395
rect 14197 7361 14231 7395
rect 17141 7361 17175 7395
rect 17509 7361 17543 7395
rect 17785 7361 17819 7395
rect 18245 7361 18279 7395
rect 18521 7361 18555 7395
rect 22569 7361 22603 7395
rect 23489 7361 23523 7395
rect 26985 7361 27019 7395
rect 1777 7293 1811 7327
rect 2421 7293 2455 7327
rect 2973 7293 3007 7327
rect 4813 7293 4847 7327
rect 6377 7293 6411 7327
rect 9965 7293 9999 7327
rect 14473 7293 14507 7327
rect 17325 7293 17359 7327
rect 24409 7293 24443 7327
rect 17693 7225 17727 7259
rect 17969 7225 18003 7259
rect 19809 7225 19843 7259
rect 24225 7225 24259 7259
rect 26617 7225 26651 7259
rect 7757 7157 7791 7191
rect 8401 7157 8435 7191
rect 13277 7157 13311 7191
rect 13921 7157 13955 7191
rect 16129 7157 16163 7191
rect 22385 7157 22419 7191
rect 10333 6953 10367 6987
rect 11529 6953 11563 6987
rect 14473 6953 14507 6987
rect 18521 6953 18555 6987
rect 22661 6953 22695 6987
rect 24685 6953 24719 6987
rect 27169 6953 27203 6987
rect 6837 6885 6871 6919
rect 11345 6885 11379 6919
rect 14657 6885 14691 6919
rect 21005 6885 21039 6919
rect 22845 6885 22879 6919
rect 6653 6817 6687 6851
rect 7389 6817 7423 6851
rect 9597 6817 9631 6851
rect 11069 6817 11103 6851
rect 1593 6749 1627 6783
rect 1777 6749 1811 6783
rect 3617 6749 3651 6783
rect 3918 6757 3952 6791
rect 6377 6749 6411 6783
rect 7656 6749 7690 6783
rect 8953 6749 8987 6783
rect 9413 6749 9447 6783
rect 10517 6749 10551 6783
rect 13185 6749 13219 6783
rect 17141 6749 17175 6783
rect 21189 6749 21223 6783
rect 23213 6749 23247 6783
rect 24869 6749 24903 6783
rect 25789 6749 25823 6783
rect 1869 6681 1903 6715
rect 7113 6681 7147 6715
rect 9111 6681 9145 6715
rect 9229 6681 9263 6715
rect 9321 6681 9355 6715
rect 9873 6681 9907 6715
rect 10057 6681 10091 6715
rect 14933 6681 14967 6715
rect 17408 6681 17442 6715
rect 20637 6681 20671 6715
rect 21456 6681 21490 6715
rect 23121 6681 23155 6715
rect 26056 6681 26090 6715
rect 3847 6613 3881 6647
rect 6561 6613 6595 6647
rect 8769 6613 8803 6647
rect 9689 6613 9723 6647
rect 13369 6613 13403 6647
rect 21097 6613 21131 6647
rect 22569 6613 22603 6647
rect 23397 6613 23431 6647
rect 4629 6409 4663 6443
rect 6101 6409 6135 6443
rect 8125 6409 8159 6443
rect 8953 6409 8987 6443
rect 17785 6409 17819 6443
rect 20085 6409 20119 6443
rect 21833 6409 21867 6443
rect 23673 6409 23707 6443
rect 25329 6409 25363 6443
rect 26157 6409 26191 6443
rect 4966 6341 5000 6375
rect 6990 6341 7024 6375
rect 9290 6341 9324 6375
rect 12541 6341 12575 6375
rect 12746 6341 12780 6375
rect 14473 6341 14507 6375
rect 16037 6341 16071 6375
rect 16237 6341 16271 6375
rect 22538 6341 22572 6375
rect 23765 6341 23799 6375
rect 24593 6341 24627 6375
rect 25605 6341 25639 6375
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 2237 6273 2271 6307
rect 3224 6273 3258 6307
rect 4445 6273 4479 6307
rect 6745 6273 6779 6307
rect 8769 6273 8803 6307
rect 13001 6273 13035 6307
rect 13185 6273 13219 6307
rect 17601 6273 17635 6307
rect 18337 6273 18371 6307
rect 18889 6273 18923 6307
rect 20637 6273 20671 6307
rect 20821 6273 20855 6307
rect 21097 6273 21131 6307
rect 22017 6273 22051 6307
rect 24317 6273 24351 6307
rect 25237 6273 25271 6307
rect 26341 6273 26375 6307
rect 4721 6205 4755 6239
rect 9045 6205 9079 6239
rect 18797 6205 18831 6239
rect 20453 6205 20487 6239
rect 20913 6205 20947 6239
rect 21281 6205 21315 6239
rect 22293 6205 22327 6239
rect 24225 6205 24259 6239
rect 26065 6205 26099 6239
rect 1593 6137 1627 6171
rect 14841 6137 14875 6171
rect 18613 6137 18647 6171
rect 24041 6137 24075 6171
rect 24869 6137 24903 6171
rect 25881 6137 25915 6171
rect 3295 6069 3329 6103
rect 10425 6069 10459 6103
rect 12725 6069 12759 6103
rect 12909 6069 12943 6103
rect 13369 6069 13403 6103
rect 14933 6069 14967 6103
rect 16221 6069 16255 6103
rect 16405 6069 16439 6103
rect 19073 6069 19107 6103
rect 20361 6069 20395 6103
rect 20545 6069 20579 6103
rect 24501 6069 24535 6103
rect 25053 6069 25087 6103
rect 5641 5865 5675 5899
rect 12725 5865 12759 5899
rect 13185 5865 13219 5899
rect 13553 5865 13587 5899
rect 16957 5865 16991 5899
rect 17233 5865 17267 5899
rect 17693 5865 17727 5899
rect 17877 5865 17911 5899
rect 17969 5865 18003 5899
rect 18153 5865 18187 5899
rect 18613 5865 18647 5899
rect 20729 5865 20763 5899
rect 20913 5865 20947 5899
rect 24409 5865 24443 5899
rect 7849 5797 7883 5831
rect 10241 5797 10275 5831
rect 11989 5797 12023 5831
rect 13645 5797 13679 5831
rect 15761 5797 15795 5831
rect 16497 5797 16531 5831
rect 17049 5797 17083 5831
rect 18429 5797 18463 5831
rect 20637 5797 20671 5831
rect 4261 5729 4295 5763
rect 8125 5729 8159 5763
rect 10609 5729 10643 5763
rect 16589 5729 16623 5763
rect 3985 5661 4019 5695
rect 6101 5661 6135 5695
rect 9597 5661 9631 5695
rect 10057 5661 10091 5695
rect 10333 5661 10367 5695
rect 12081 5661 12115 5695
rect 12357 5661 12391 5695
rect 12449 5661 12483 5695
rect 12541 5661 12575 5695
rect 13461 5661 13495 5695
rect 13737 5661 13771 5695
rect 13921 5661 13955 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 16221 5661 16255 5695
rect 16681 5661 16715 5695
rect 19257 5661 19291 5695
rect 19513 5661 19547 5695
rect 25522 5661 25556 5695
rect 25789 5661 25823 5695
rect 25881 5661 25915 5695
rect 17739 5627 17773 5661
rect 4506 5593 4540 5627
rect 6368 5593 6402 5627
rect 9755 5593 9789 5627
rect 9873 5593 9907 5627
rect 9965 5593 9999 5627
rect 10854 5593 10888 5627
rect 12239 5593 12273 5627
rect 14648 5593 14682 5627
rect 17417 5593 17451 5627
rect 17509 5593 17543 5627
rect 18337 5593 18371 5627
rect 18797 5593 18831 5627
rect 21097 5593 21131 5627
rect 4169 5525 4203 5559
rect 7481 5525 7515 5559
rect 7665 5525 7699 5559
rect 10517 5525 10551 5559
rect 14105 5525 14139 5559
rect 16313 5525 16347 5559
rect 17207 5525 17241 5559
rect 18137 5525 18171 5559
rect 18597 5525 18631 5559
rect 20887 5525 20921 5559
rect 26065 5525 26099 5559
rect 4721 5321 4755 5355
rect 5273 5321 5307 5355
rect 7021 5321 7055 5355
rect 7757 5321 7791 5355
rect 10609 5321 10643 5355
rect 12909 5321 12943 5355
rect 14657 5321 14691 5355
rect 14749 5321 14783 5355
rect 15837 5321 15871 5355
rect 16329 5321 16363 5355
rect 16497 5321 16531 5355
rect 18500 5321 18534 5355
rect 20545 5321 20579 5355
rect 22645 5321 22679 5355
rect 24133 5321 24167 5355
rect 24961 5321 24995 5355
rect 5733 5253 5767 5287
rect 6745 5253 6779 5287
rect 6929 5253 6963 5287
rect 8094 5253 8128 5287
rect 10425 5253 10459 5287
rect 11621 5253 11655 5287
rect 11805 5253 11839 5287
rect 12541 5253 12575 5287
rect 12757 5253 12791 5287
rect 13544 5253 13578 5287
rect 16037 5253 16071 5287
rect 16129 5253 16163 5287
rect 18705 5253 18739 5287
rect 20177 5253 20211 5287
rect 20393 5253 20427 5287
rect 22845 5253 22879 5287
rect 26074 5253 26108 5287
rect 5181 5185 5215 5219
rect 7205 5185 7239 5219
rect 7573 5185 7607 5219
rect 7849 5185 7883 5219
rect 10241 5185 10275 5219
rect 13277 5185 13311 5219
rect 14933 5185 14967 5219
rect 17785 5185 17819 5219
rect 18061 5185 18095 5219
rect 20637 5185 20671 5219
rect 20821 5185 20855 5219
rect 22201 5185 22235 5219
rect 23121 5185 23155 5219
rect 23213 5185 23247 5219
rect 23857 5185 23891 5219
rect 26341 5185 26375 5219
rect 6561 5117 6595 5151
rect 17877 5117 17911 5151
rect 21925 5117 21959 5151
rect 22017 5117 22051 5151
rect 22109 5117 22143 5151
rect 22385 5117 22419 5151
rect 23305 5117 23339 5151
rect 23397 5117 23431 5151
rect 4905 5049 4939 5083
rect 5457 5049 5491 5083
rect 15669 5049 15703 5083
rect 17601 5049 17635 5083
rect 18337 5049 18371 5083
rect 22477 5049 22511 5083
rect 22937 5049 22971 5083
rect 9229 4981 9263 5015
rect 11989 4981 12023 5015
rect 12725 4981 12759 5015
rect 15853 4981 15887 5015
rect 16313 4981 16347 5015
rect 18521 4981 18555 5015
rect 20361 4981 20395 5015
rect 21005 4981 21039 5015
rect 22661 4981 22695 5015
rect 5365 4777 5399 4811
rect 9321 4777 9355 4811
rect 13645 4777 13679 4811
rect 16681 4777 16715 4811
rect 18061 4777 18095 4811
rect 20637 4777 20671 4811
rect 23029 4777 23063 4811
rect 23213 4777 23247 4811
rect 7389 4709 7423 4743
rect 12725 4709 12759 4743
rect 17141 4709 17175 4743
rect 22109 4709 22143 4743
rect 12357 4641 12391 4675
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 7113 4573 7147 4607
rect 9505 4573 9539 4607
rect 9689 4573 9723 4607
rect 9965 4573 9999 4607
rect 10333 4573 10367 4607
rect 11897 4573 11931 4607
rect 13461 4573 13495 4607
rect 14289 4573 14323 4607
rect 15669 4573 15703 4607
rect 16865 4573 16899 4607
rect 16957 4573 16991 4607
rect 17877 4573 17911 4607
rect 19257 4573 19291 4607
rect 20729 4573 20763 4607
rect 22201 4573 22235 4607
rect 22385 4573 22419 4607
rect 23489 4573 23523 4607
rect 23949 4573 23983 4607
rect 1501 4505 1535 4539
rect 1685 4505 1719 4539
rect 7297 4505 7331 4539
rect 7573 4505 7607 4539
rect 9597 4505 9631 4539
rect 9807 4505 9841 4539
rect 10793 4505 10827 4539
rect 19524 4505 19558 4539
rect 20996 4505 21030 4539
rect 22569 4505 22603 4539
rect 22845 4505 22879 4539
rect 23061 4505 23095 4539
rect 23305 4505 23339 4539
rect 5641 4437 5675 4471
rect 6929 4437 6963 4471
rect 10149 4437 10183 4471
rect 11069 4437 11103 4471
rect 11713 4437 11747 4471
rect 12817 4437 12851 4471
rect 14105 4437 14139 4471
rect 15485 4437 15519 4471
rect 23673 4437 23707 4471
rect 23765 4437 23799 4471
rect 6193 4233 6227 4267
rect 9045 4233 9079 4267
rect 15025 4233 15059 4267
rect 16497 4233 16531 4267
rect 16681 4233 16715 4267
rect 19717 4233 19751 4267
rect 20913 4233 20947 4267
rect 23581 4233 23615 4267
rect 9413 4165 9447 4199
rect 9505 4165 9539 4199
rect 9643 4165 9677 4199
rect 9873 4165 9907 4199
rect 11069 4165 11103 4199
rect 11713 4165 11747 4199
rect 13912 4165 13946 4199
rect 15384 4165 15418 4199
rect 17794 4165 17828 4199
rect 19165 4165 19199 4199
rect 5080 4097 5114 4131
rect 6929 4097 6963 4131
rect 7665 4097 7699 4131
rect 7932 4097 7966 4131
rect 9137 4097 9171 4131
rect 9321 4097 9355 4131
rect 12173 4097 12207 4131
rect 12440 4097 12474 4131
rect 13645 4097 13679 4131
rect 18061 4097 18095 4131
rect 19901 4097 19935 4131
rect 20729 4097 20763 4131
rect 22468 4097 22502 4131
rect 24786 4097 24820 4131
rect 4813 4029 4847 4063
rect 9781 4029 9815 4063
rect 15117 4029 15151 4063
rect 19625 4029 19659 4063
rect 22201 4029 22235 4063
rect 25053 4029 25087 4063
rect 10149 3961 10183 3995
rect 10701 3961 10735 3995
rect 19441 3961 19475 3995
rect 6745 3893 6779 3927
rect 10333 3893 10367 3927
rect 10609 3893 10643 3927
rect 11621 3893 11655 3927
rect 13553 3893 13587 3927
rect 23673 3893 23707 3927
rect 5733 3689 5767 3723
rect 8125 3689 8159 3723
rect 11345 3689 11379 3723
rect 12817 3689 12851 3723
rect 12909 3689 12943 3723
rect 14105 3689 14139 3723
rect 15761 3689 15795 3723
rect 17141 3689 17175 3723
rect 19073 3689 19107 3723
rect 23857 3689 23891 3723
rect 5641 3621 5675 3655
rect 14197 3621 14231 3655
rect 15577 3621 15611 3655
rect 16037 3621 16071 3655
rect 16957 3621 16991 3655
rect 19533 3621 19567 3655
rect 21465 3621 21499 3655
rect 5273 3553 5307 3587
rect 6285 3553 6319 3587
rect 14565 3553 14599 3587
rect 19717 3553 19751 3587
rect 6552 3485 6586 3519
rect 8309 3485 8343 3519
rect 9689 3485 9723 3519
rect 9873 3485 9907 3519
rect 9965 3485 9999 3519
rect 11437 3485 11471 3519
rect 11704 3485 11738 3519
rect 13093 3485 13127 3519
rect 17417 3485 17451 3519
rect 17693 3485 17727 3519
rect 19809 3485 19843 3519
rect 20085 3485 20119 3519
rect 22661 3485 22695 3519
rect 23673 3485 23707 3519
rect 10232 3417 10266 3451
rect 15301 3417 15335 3451
rect 16313 3417 16347 3451
rect 16681 3417 16715 3451
rect 17938 3417 17972 3451
rect 19257 3417 19291 3451
rect 20330 3417 20364 3451
rect 7665 3349 7699 3383
rect 15853 3349 15887 3383
rect 17601 3349 17635 3383
rect 19993 3349 20027 3383
rect 22845 3349 22879 3383
rect 10149 3145 10183 3179
rect 16221 3145 16255 3179
rect 17693 3145 17727 3179
rect 22477 3145 22511 3179
rect 9781 3077 9815 3111
rect 18153 3077 18187 3111
rect 19993 3077 20027 3111
rect 22385 3077 22419 3111
rect 23590 3077 23624 3111
rect 8677 3009 8711 3043
rect 9965 3009 9999 3043
rect 12357 3009 12391 3043
rect 15108 3009 15142 3043
rect 21005 3009 21039 3043
rect 9321 2941 9355 2975
rect 12081 2941 12115 2975
rect 12173 2941 12207 2975
rect 14841 2941 14875 2975
rect 21925 2941 21959 2975
rect 23857 2941 23891 2975
rect 9505 2873 9539 2907
rect 11713 2873 11747 2907
rect 17877 2873 17911 2907
rect 19717 2873 19751 2907
rect 22109 2873 22143 2907
rect 8493 2805 8527 2839
rect 11621 2805 11655 2839
rect 19533 2805 19567 2839
rect 20821 2805 20855 2839
rect 8125 2601 8159 2635
rect 13369 2601 13403 2635
rect 15393 2601 15427 2635
rect 18245 2601 18279 2635
rect 22109 2601 22143 2635
rect 22753 2601 22787 2635
rect 9229 2533 9263 2567
rect 10977 2533 11011 2567
rect 13737 2533 13771 2567
rect 19257 2533 19291 2567
rect 22569 2533 22603 2567
rect 6745 2465 6779 2499
rect 8953 2465 8987 2499
rect 9413 2465 9447 2499
rect 11253 2465 11287 2499
rect 11989 2465 12023 2499
rect 13921 2465 13955 2499
rect 9689 2397 9723 2431
rect 10057 2397 10091 2431
rect 11713 2397 11747 2431
rect 14105 2397 14139 2431
rect 15577 2397 15611 2431
rect 16865 2397 16899 2431
rect 20637 2397 20671 2431
rect 20729 2397 20763 2431
rect 20985 2397 21019 2431
rect 7012 2329 7046 2363
rect 12234 2329 12268 2363
rect 13461 2329 13495 2363
rect 17110 2329 17144 2363
rect 20370 2329 20404 2363
rect 22293 2329 22327 2363
rect 9505 2261 9539 2295
rect 10241 2261 10275 2295
rect 10793 2261 10827 2295
rect 11897 2261 11931 2295
rect 14289 2261 14323 2295
rect 7205 2057 7239 2091
rect 9321 2057 9355 2091
rect 9873 2057 9907 2091
rect 14565 2057 14599 2091
rect 16497 2057 16531 2091
rect 18705 2057 18739 2091
rect 19625 2057 19659 2091
rect 21649 2057 21683 2091
rect 23213 2057 23247 2091
rect 8208 1989 8242 2023
rect 9413 1989 9447 2023
rect 10232 1989 10266 2023
rect 11529 1989 11563 2023
rect 14994 1989 15028 2023
rect 22078 1989 22112 2023
rect 7389 1921 7423 1955
rect 9965 1921 9999 1955
rect 12081 1921 12115 1955
rect 12337 1921 12371 1955
rect 13645 1921 13679 1955
rect 14381 1921 14415 1955
rect 16313 1921 16347 1955
rect 17325 1921 17359 1955
rect 17581 1921 17615 1955
rect 18797 1921 18831 1955
rect 19441 1921 19475 1955
rect 20157 1921 20191 1955
rect 21465 1921 21499 1955
rect 21833 1921 21867 1955
rect 7941 1853 7975 1887
rect 14105 1853 14139 1887
rect 14749 1853 14783 1887
rect 16681 1853 16715 1887
rect 17141 1853 17175 1887
rect 19901 1853 19935 1887
rect 9781 1785 9815 1819
rect 11345 1785 11379 1819
rect 11897 1785 11931 1819
rect 13921 1785 13955 1819
rect 16773 1785 16807 1819
rect 19073 1785 19107 1819
rect 11989 1717 12023 1751
rect 13461 1717 13495 1751
rect 16129 1717 16163 1751
rect 19257 1717 19291 1751
rect 21281 1717 21315 1751
rect 10333 1513 10367 1547
rect 12173 1513 12207 1547
rect 15485 1513 15519 1547
rect 17417 1513 17451 1547
rect 19625 1513 19659 1547
rect 21833 1513 21867 1547
rect 17049 1445 17083 1479
rect 22017 1445 22051 1479
rect 8953 1377 8987 1411
rect 22293 1377 22327 1411
rect 9220 1309 9254 1343
rect 11989 1309 12023 1343
rect 14105 1309 14139 1343
rect 14372 1309 14406 1343
rect 16681 1309 16715 1343
rect 17233 1309 17267 1343
rect 19441 1309 19475 1343
rect 17141 1173 17175 1207
<< metal1 >>
rect 1104 32666 29048 32688
rect 1104 32614 7896 32666
rect 7948 32614 7960 32666
rect 8012 32614 8024 32666
rect 8076 32614 8088 32666
rect 8140 32614 8152 32666
rect 8204 32614 14842 32666
rect 14894 32614 14906 32666
rect 14958 32614 14970 32666
rect 15022 32614 15034 32666
rect 15086 32614 15098 32666
rect 15150 32614 21788 32666
rect 21840 32614 21852 32666
rect 21904 32614 21916 32666
rect 21968 32614 21980 32666
rect 22032 32614 22044 32666
rect 22096 32614 28734 32666
rect 28786 32614 28798 32666
rect 28850 32614 28862 32666
rect 28914 32614 28926 32666
rect 28978 32614 28990 32666
rect 29042 32614 29048 32666
rect 1104 32592 29048 32614
rect 4709 32419 4767 32425
rect 4709 32416 4721 32419
rect 3988 32388 4721 32416
rect 3988 32360 4016 32388
rect 4709 32385 4721 32388
rect 4755 32416 4767 32419
rect 4801 32419 4859 32425
rect 4801 32416 4813 32419
rect 4755 32388 4813 32416
rect 4755 32385 4767 32388
rect 4709 32379 4767 32385
rect 4801 32385 4813 32388
rect 4847 32385 4859 32419
rect 8573 32419 8631 32425
rect 8573 32416 8585 32419
rect 4801 32379 4859 32385
rect 8128 32388 8585 32416
rect 3881 32351 3939 32357
rect 3881 32317 3893 32351
rect 3927 32348 3939 32351
rect 3970 32348 3976 32360
rect 3927 32320 3976 32348
rect 3927 32317 3939 32320
rect 3881 32311 3939 32317
rect 3970 32308 3976 32320
rect 4028 32308 4034 32360
rect 4246 32308 4252 32360
rect 4304 32348 4310 32360
rect 4341 32351 4399 32357
rect 4341 32348 4353 32351
rect 4304 32320 4353 32348
rect 4304 32308 4310 32320
rect 4341 32317 4353 32320
rect 4387 32348 4399 32351
rect 5169 32351 5227 32357
rect 5169 32348 5181 32351
rect 4387 32320 5181 32348
rect 4387 32317 4399 32320
rect 4341 32311 4399 32317
rect 5169 32317 5181 32320
rect 5215 32317 5227 32351
rect 5169 32311 5227 32317
rect 6365 32351 6423 32357
rect 6365 32317 6377 32351
rect 6411 32317 6423 32351
rect 6365 32311 6423 32317
rect 4249 32215 4307 32221
rect 4249 32181 4261 32215
rect 4295 32212 4307 32215
rect 4338 32212 4344 32224
rect 4295 32184 4344 32212
rect 4295 32181 4307 32184
rect 4249 32175 4307 32181
rect 4338 32172 4344 32184
rect 4396 32212 4402 32224
rect 6380 32221 6408 32311
rect 6454 32308 6460 32360
rect 6512 32348 6518 32360
rect 6733 32351 6791 32357
rect 6733 32348 6745 32351
rect 6512 32320 6745 32348
rect 6512 32308 6518 32320
rect 6733 32317 6745 32320
rect 6779 32348 6791 32351
rect 6825 32351 6883 32357
rect 6825 32348 6837 32351
rect 6779 32320 6837 32348
rect 6779 32317 6791 32320
rect 6733 32311 6791 32317
rect 6825 32317 6837 32320
rect 6871 32317 6883 32351
rect 6825 32311 6883 32317
rect 7193 32351 7251 32357
rect 7193 32317 7205 32351
rect 7239 32317 7251 32351
rect 7193 32311 7251 32317
rect 7745 32351 7803 32357
rect 7745 32317 7757 32351
rect 7791 32317 7803 32351
rect 7745 32311 7803 32317
rect 7208 32221 7236 32311
rect 7760 32221 7788 32311
rect 7834 32308 7840 32360
rect 7892 32348 7898 32360
rect 8128 32357 8156 32388
rect 8573 32385 8585 32388
rect 8619 32385 8631 32419
rect 8573 32379 8631 32385
rect 8113 32351 8171 32357
rect 8113 32348 8125 32351
rect 7892 32320 8125 32348
rect 7892 32308 7898 32320
rect 8113 32317 8125 32320
rect 8159 32317 8171 32351
rect 8113 32311 8171 32317
rect 8205 32351 8263 32357
rect 8205 32317 8217 32351
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 9309 32351 9367 32357
rect 9309 32317 9321 32351
rect 9355 32317 9367 32351
rect 9309 32311 9367 32317
rect 8220 32221 8248 32311
rect 9324 32221 9352 32311
rect 9582 32308 9588 32360
rect 9640 32348 9646 32360
rect 9677 32351 9735 32357
rect 9677 32348 9689 32351
rect 9640 32320 9689 32348
rect 9640 32308 9646 32320
rect 9677 32317 9689 32320
rect 9723 32317 9735 32351
rect 9677 32311 9735 32317
rect 5169 32215 5227 32221
rect 5169 32212 5181 32215
rect 4396 32184 5181 32212
rect 4396 32172 4402 32184
rect 5169 32181 5181 32184
rect 5215 32212 5227 32215
rect 6365 32215 6423 32221
rect 6365 32212 6377 32215
rect 5215 32184 6377 32212
rect 5215 32181 5227 32184
rect 5169 32175 5227 32181
rect 6365 32181 6377 32184
rect 6411 32212 6423 32215
rect 7193 32215 7251 32221
rect 7193 32212 7205 32215
rect 6411 32184 7205 32212
rect 6411 32181 6423 32184
rect 6365 32175 6423 32181
rect 7193 32181 7205 32184
rect 7239 32212 7251 32215
rect 7745 32215 7803 32221
rect 7745 32212 7757 32215
rect 7239 32184 7757 32212
rect 7239 32181 7251 32184
rect 7193 32175 7251 32181
rect 7745 32181 7757 32184
rect 7791 32212 7803 32215
rect 8205 32215 8263 32221
rect 8205 32212 8217 32215
rect 7791 32184 8217 32212
rect 7791 32181 7803 32184
rect 7745 32175 7803 32181
rect 8205 32181 8217 32184
rect 8251 32212 8263 32215
rect 9309 32215 9367 32221
rect 9309 32212 9321 32215
rect 8251 32184 9321 32212
rect 8251 32181 8263 32184
rect 8205 32175 8263 32181
rect 9309 32181 9321 32184
rect 9355 32181 9367 32215
rect 9309 32175 9367 32181
rect 11054 32172 11060 32224
rect 11112 32172 11118 32224
rect 1104 32122 28888 32144
rect 1104 32070 4423 32122
rect 4475 32070 4487 32122
rect 4539 32070 4551 32122
rect 4603 32070 4615 32122
rect 4667 32070 4679 32122
rect 4731 32070 11369 32122
rect 11421 32070 11433 32122
rect 11485 32070 11497 32122
rect 11549 32070 11561 32122
rect 11613 32070 11625 32122
rect 11677 32070 18315 32122
rect 18367 32070 18379 32122
rect 18431 32070 18443 32122
rect 18495 32070 18507 32122
rect 18559 32070 18571 32122
rect 18623 32070 25261 32122
rect 25313 32070 25325 32122
rect 25377 32070 25389 32122
rect 25441 32070 25453 32122
rect 25505 32070 25517 32122
rect 25569 32070 28888 32122
rect 1104 32048 28888 32070
rect 11054 31968 11060 32020
rect 11112 31968 11118 32020
rect 4246 31900 4252 31952
rect 4304 31940 4310 31952
rect 4709 31943 4767 31949
rect 4709 31940 4721 31943
rect 4304 31912 4721 31940
rect 4304 31900 4310 31912
rect 4709 31909 4721 31912
rect 4755 31909 4767 31943
rect 4709 31903 4767 31909
rect 4341 31875 4399 31881
rect 4341 31841 4353 31875
rect 4387 31841 4399 31875
rect 5537 31875 5595 31881
rect 5537 31872 5549 31875
rect 4341 31835 4399 31841
rect 5092 31844 5549 31872
rect 3881 31807 3939 31813
rect 3881 31773 3893 31807
rect 3927 31804 3939 31807
rect 3970 31804 3976 31816
rect 3927 31776 3976 31804
rect 3927 31773 3939 31776
rect 3881 31767 3939 31773
rect 3970 31764 3976 31776
rect 4028 31804 4034 31816
rect 4356 31804 4384 31835
rect 4028 31776 4384 31804
rect 4028 31764 4034 31776
rect 4982 31764 4988 31816
rect 5040 31804 5046 31816
rect 5092 31813 5120 31844
rect 5537 31841 5549 31844
rect 5583 31872 5595 31875
rect 5997 31875 6055 31881
rect 5997 31872 6009 31875
rect 5583 31844 6009 31872
rect 5583 31841 5595 31844
rect 5537 31835 5595 31841
rect 5997 31841 6009 31844
rect 6043 31872 6055 31875
rect 6454 31872 6460 31884
rect 6043 31844 6460 31872
rect 6043 31841 6055 31844
rect 5997 31835 6055 31841
rect 6454 31832 6460 31844
rect 6512 31832 6518 31884
rect 7834 31872 7840 31884
rect 7392 31844 7840 31872
rect 5077 31807 5135 31813
rect 5077 31804 5089 31807
rect 5040 31776 5089 31804
rect 5040 31764 5046 31776
rect 5077 31773 5089 31776
rect 5123 31773 5135 31807
rect 5077 31767 5135 31773
rect 5445 31807 5503 31813
rect 5445 31773 5457 31807
rect 5491 31773 5503 31807
rect 5445 31767 5503 31773
rect 5905 31807 5963 31813
rect 5905 31773 5917 31807
rect 5951 31773 5963 31807
rect 5905 31767 5963 31773
rect 6365 31807 6423 31813
rect 6365 31773 6377 31807
rect 6411 31773 6423 31807
rect 6365 31767 6423 31773
rect 6825 31807 6883 31813
rect 6825 31773 6837 31807
rect 6871 31804 6883 31807
rect 6917 31807 6975 31813
rect 6917 31804 6929 31807
rect 6871 31776 6929 31804
rect 6871 31773 6883 31776
rect 6825 31767 6883 31773
rect 6917 31773 6929 31776
rect 6963 31773 6975 31807
rect 6917 31767 6975 31773
rect 5460 31736 5488 31767
rect 5920 31736 5948 31767
rect 6380 31736 6408 31767
rect 6840 31736 6868 31767
rect 7282 31764 7288 31816
rect 7340 31804 7346 31816
rect 7392 31813 7420 31844
rect 7834 31832 7840 31844
rect 7892 31832 7898 31884
rect 8757 31875 8815 31881
rect 8757 31841 8769 31875
rect 8803 31872 8815 31875
rect 9582 31872 9588 31884
rect 8803 31844 9588 31872
rect 8803 31841 8815 31844
rect 8757 31835 8815 31841
rect 9324 31816 9352 31844
rect 9582 31832 9588 31844
rect 9640 31872 9646 31884
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 9640 31844 9781 31872
rect 9640 31832 9646 31844
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 10229 31875 10287 31881
rect 10229 31872 10241 31875
rect 9769 31835 9827 31841
rect 9876 31844 10241 31872
rect 7377 31807 7435 31813
rect 7377 31804 7389 31807
rect 7340 31776 7389 31804
rect 7340 31764 7346 31776
rect 7377 31773 7389 31776
rect 7423 31773 7435 31807
rect 7377 31767 7435 31773
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31773 7803 31807
rect 7745 31767 7803 31773
rect 8205 31807 8263 31813
rect 8205 31773 8217 31807
rect 8251 31804 8263 31807
rect 8389 31807 8447 31813
rect 8389 31804 8401 31807
rect 8251 31776 8401 31804
rect 8251 31773 8263 31776
rect 8205 31767 8263 31773
rect 8389 31773 8401 31776
rect 8435 31773 8447 31807
rect 8389 31767 8447 31773
rect 7760 31736 7788 31767
rect 8220 31736 8248 31767
rect 8662 31764 8668 31816
rect 8720 31804 8726 31816
rect 8941 31807 8999 31813
rect 8941 31804 8953 31807
rect 8720 31776 8953 31804
rect 8720 31764 8726 31776
rect 8941 31773 8953 31776
rect 8987 31773 8999 31807
rect 8941 31767 8999 31773
rect 9306 31764 9312 31816
rect 9364 31764 9370 31816
rect 9674 31764 9680 31816
rect 9732 31764 9738 31816
rect 9876 31804 9904 31844
rect 10229 31841 10241 31844
rect 10275 31841 10287 31875
rect 11072 31872 11100 31968
rect 11149 31875 11207 31881
rect 11149 31872 11161 31875
rect 11072 31844 11161 31872
rect 10229 31835 10287 31841
rect 11149 31841 11161 31844
rect 11195 31841 11207 31875
rect 11149 31835 11207 31841
rect 9784 31776 9904 31804
rect 10137 31807 10195 31813
rect 9784 31736 9812 31776
rect 10137 31773 10149 31807
rect 10183 31773 10195 31807
rect 10137 31767 10195 31773
rect 10597 31807 10655 31813
rect 10597 31773 10609 31807
rect 10643 31804 10655 31807
rect 10781 31807 10839 31813
rect 10781 31804 10793 31807
rect 10643 31776 10793 31804
rect 10643 31773 10655 31776
rect 10597 31767 10655 31773
rect 10781 31773 10793 31776
rect 10827 31773 10839 31807
rect 10781 31767 10839 31773
rect 5460 31708 8248 31736
rect 4249 31671 4307 31677
rect 4249 31637 4261 31671
rect 4295 31668 4307 31671
rect 4338 31668 4344 31680
rect 4295 31640 4344 31668
rect 4295 31637 4307 31640
rect 4249 31631 4307 31637
rect 4338 31628 4344 31640
rect 4396 31668 4402 31680
rect 5460 31677 5488 31708
rect 5920 31677 5948 31708
rect 6380 31677 6408 31708
rect 6840 31677 6868 31708
rect 7760 31677 7788 31708
rect 8220 31677 8248 31708
rect 9600 31708 9812 31736
rect 10152 31736 10180 31767
rect 10612 31736 10640 31767
rect 10152 31708 10640 31736
rect 9600 31680 9628 31708
rect 4709 31671 4767 31677
rect 4709 31668 4721 31671
rect 4396 31640 4721 31668
rect 4396 31628 4402 31640
rect 4709 31637 4721 31640
rect 4755 31668 4767 31671
rect 5445 31671 5503 31677
rect 5445 31668 5457 31671
rect 4755 31640 5457 31668
rect 4755 31637 4767 31640
rect 4709 31631 4767 31637
rect 5445 31637 5457 31640
rect 5491 31637 5503 31671
rect 5445 31631 5503 31637
rect 5905 31671 5963 31677
rect 5905 31637 5917 31671
rect 5951 31668 5963 31671
rect 6365 31671 6423 31677
rect 5951 31640 5985 31668
rect 5951 31637 5963 31640
rect 5905 31631 5963 31637
rect 6365 31637 6377 31671
rect 6411 31668 6423 31671
rect 6825 31671 6883 31677
rect 6411 31640 6445 31668
rect 6411 31637 6423 31640
rect 6365 31631 6423 31637
rect 6825 31637 6837 31671
rect 6871 31668 6883 31671
rect 6917 31671 6975 31677
rect 6917 31668 6929 31671
rect 6871 31640 6929 31668
rect 6871 31637 6883 31640
rect 6825 31631 6883 31637
rect 6917 31637 6929 31640
rect 6963 31637 6975 31671
rect 6917 31631 6975 31637
rect 7745 31671 7803 31677
rect 7745 31637 7757 31671
rect 7791 31668 7803 31671
rect 8205 31671 8263 31677
rect 7791 31640 7825 31668
rect 7791 31637 7803 31640
rect 7745 31631 7803 31637
rect 8205 31637 8217 31671
rect 8251 31668 8263 31671
rect 8389 31671 8447 31677
rect 8389 31668 8401 31671
rect 8251 31640 8401 31668
rect 8251 31637 8263 31640
rect 8205 31631 8263 31637
rect 8389 31637 8401 31640
rect 8435 31637 8447 31671
rect 8389 31631 8447 31637
rect 9125 31671 9183 31677
rect 9125 31637 9137 31671
rect 9171 31668 9183 31671
rect 9582 31668 9588 31680
rect 9171 31640 9588 31668
rect 9171 31637 9183 31640
rect 9125 31631 9183 31637
rect 9582 31628 9588 31640
rect 9640 31628 9646 31680
rect 9674 31628 9680 31680
rect 9732 31668 9738 31680
rect 10152 31677 10180 31708
rect 10612 31677 10640 31708
rect 10137 31671 10195 31677
rect 10137 31668 10149 31671
rect 9732 31640 10149 31668
rect 9732 31628 9738 31640
rect 10137 31637 10149 31640
rect 10183 31637 10195 31671
rect 10137 31631 10195 31637
rect 10597 31671 10655 31677
rect 10597 31637 10609 31671
rect 10643 31668 10655 31671
rect 10781 31671 10839 31677
rect 10781 31668 10793 31671
rect 10643 31640 10793 31668
rect 10643 31637 10655 31640
rect 10597 31631 10655 31637
rect 10781 31637 10793 31640
rect 10827 31637 10839 31671
rect 10781 31631 10839 31637
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 1949 31467 2007 31473
rect 1949 31433 1961 31467
rect 1995 31464 2007 31467
rect 2406 31464 2412 31476
rect 1995 31436 2412 31464
rect 1995 31433 2007 31436
rect 1949 31427 2007 31433
rect 1964 31337 1992 31427
rect 2406 31424 2412 31436
rect 2464 31424 2470 31476
rect 3237 31467 3295 31473
rect 3237 31464 3249 31467
rect 3068 31436 3249 31464
rect 1949 31331 2007 31337
rect 1949 31297 1961 31331
rect 1995 31297 2007 31331
rect 1949 31291 2007 31297
rect 2317 31331 2375 31337
rect 2317 31297 2329 31331
rect 2363 31328 2375 31331
rect 2498 31328 2504 31340
rect 2363 31300 2504 31328
rect 2363 31297 2375 31300
rect 2317 31291 2375 31297
rect 2498 31288 2504 31300
rect 2556 31328 2562 31340
rect 2777 31331 2835 31337
rect 2777 31328 2789 31331
rect 2556 31300 2789 31328
rect 2556 31288 2562 31300
rect 2777 31297 2789 31300
rect 2823 31328 2835 31331
rect 2869 31331 2927 31337
rect 2869 31328 2881 31331
rect 2823 31300 2881 31328
rect 2823 31297 2835 31300
rect 2777 31291 2835 31297
rect 2869 31297 2881 31300
rect 2915 31297 2927 31331
rect 2869 31291 2927 31297
rect 2409 31263 2467 31269
rect 2409 31229 2421 31263
rect 2455 31260 2467 31263
rect 3068 31260 3096 31436
rect 3237 31433 3249 31436
rect 3283 31464 3295 31467
rect 4249 31467 4307 31473
rect 4249 31464 4261 31467
rect 3283 31436 4261 31464
rect 3283 31433 3295 31436
rect 3237 31427 3295 31433
rect 4249 31433 4261 31436
rect 4295 31464 4307 31467
rect 4338 31464 4344 31476
rect 4295 31436 4344 31464
rect 4295 31433 4307 31436
rect 4249 31427 4307 31433
rect 4338 31424 4344 31436
rect 4396 31464 4402 31476
rect 5169 31467 5227 31473
rect 5169 31464 5181 31467
rect 4396 31436 5181 31464
rect 4396 31424 4402 31436
rect 5169 31433 5181 31436
rect 5215 31464 5227 31467
rect 6181 31467 6239 31473
rect 6181 31464 6193 31467
rect 5215 31436 6193 31464
rect 5215 31433 5227 31436
rect 5169 31427 5227 31433
rect 6181 31433 6193 31436
rect 6227 31433 6239 31467
rect 6181 31427 6239 31433
rect 6733 31467 6791 31473
rect 6733 31433 6745 31467
rect 6779 31464 6791 31467
rect 7561 31467 7619 31473
rect 7561 31464 7573 31467
rect 6779 31436 7573 31464
rect 6779 31433 6791 31436
rect 6733 31427 6791 31433
rect 7561 31433 7573 31436
rect 7607 31464 7619 31467
rect 8021 31467 8079 31473
rect 8021 31464 8033 31467
rect 7607 31436 8033 31464
rect 7607 31433 7619 31436
rect 7561 31427 7619 31433
rect 8021 31433 8033 31436
rect 8067 31464 8079 31467
rect 8481 31467 8539 31473
rect 8481 31464 8493 31467
rect 8067 31436 8493 31464
rect 8067 31433 8079 31436
rect 8021 31427 8079 31433
rect 8481 31433 8493 31436
rect 8527 31433 8539 31467
rect 8481 31427 8539 31433
rect 4264 31368 5212 31396
rect 4264 31340 4292 31368
rect 3881 31331 3939 31337
rect 3881 31297 3893 31331
rect 3927 31328 3939 31331
rect 3970 31328 3976 31340
rect 3927 31300 3976 31328
rect 3927 31297 3939 31300
rect 3881 31291 3939 31297
rect 3970 31288 3976 31300
rect 4028 31288 4034 31340
rect 4246 31288 4252 31340
rect 4304 31288 4310 31340
rect 4433 31331 4491 31337
rect 4433 31297 4445 31331
rect 4479 31297 4491 31331
rect 4433 31291 4491 31297
rect 4525 31331 4583 31337
rect 4525 31297 4537 31331
rect 4571 31328 4583 31331
rect 4982 31328 4988 31340
rect 4571 31300 4988 31328
rect 4571 31297 4583 31300
rect 4525 31291 4583 31297
rect 2455 31232 3096 31260
rect 4448 31260 4476 31291
rect 4982 31288 4988 31300
rect 5040 31288 5046 31340
rect 5184 31337 5212 31368
rect 6196 31337 6224 31427
rect 6748 31337 6776 31427
rect 5169 31331 5227 31337
rect 5169 31297 5181 31331
rect 5215 31297 5227 31331
rect 5169 31291 5227 31297
rect 6181 31331 6239 31337
rect 6181 31297 6193 31331
rect 6227 31328 6239 31331
rect 6733 31331 6791 31337
rect 6733 31328 6745 31331
rect 6227 31300 6745 31328
rect 6227 31297 6239 31300
rect 6181 31291 6239 31297
rect 6733 31297 6745 31300
rect 6779 31297 6791 31331
rect 6733 31291 6791 31297
rect 7193 31331 7251 31337
rect 7193 31297 7205 31331
rect 7239 31328 7251 31331
rect 7282 31328 7288 31340
rect 7239 31300 7288 31328
rect 7239 31297 7251 31300
rect 7193 31291 7251 31297
rect 4709 31263 4767 31269
rect 4448 31232 4568 31260
rect 2455 31229 2467 31232
rect 2409 31223 2467 31229
rect 3068 31204 3096 31232
rect 1872 31164 2912 31192
rect 1872 31136 1900 31164
rect 1854 31084 1860 31136
rect 1912 31084 1918 31136
rect 2406 31084 2412 31136
rect 2464 31124 2470 31136
rect 2774 31124 2780 31136
rect 2464 31096 2780 31124
rect 2464 31084 2470 31096
rect 2774 31084 2780 31096
rect 2832 31084 2838 31136
rect 2884 31124 2912 31164
rect 3050 31152 3056 31204
rect 3108 31192 3114 31204
rect 3237 31195 3295 31201
rect 3237 31192 3249 31195
rect 3108 31164 3249 31192
rect 3108 31152 3114 31164
rect 3237 31161 3249 31164
rect 3283 31161 3295 31195
rect 3237 31155 3295 31161
rect 4540 31192 4568 31232
rect 4709 31229 4721 31263
rect 4755 31260 4767 31263
rect 4798 31260 4804 31272
rect 4755 31232 4804 31260
rect 4755 31229 4767 31232
rect 4709 31223 4767 31229
rect 4798 31220 4804 31232
rect 4856 31220 4862 31272
rect 5000 31260 5028 31288
rect 5813 31263 5871 31269
rect 5813 31260 5825 31263
rect 5000 31232 5825 31260
rect 5813 31229 5825 31232
rect 5859 31260 5871 31263
rect 6365 31263 6423 31269
rect 6365 31260 6377 31263
rect 5859 31232 6377 31260
rect 5859 31229 5871 31232
rect 5813 31223 5871 31229
rect 6365 31229 6377 31232
rect 6411 31229 6423 31263
rect 6748 31260 6776 31291
rect 7282 31288 7288 31300
rect 7340 31328 7346 31340
rect 7653 31331 7711 31337
rect 7653 31328 7665 31331
rect 7340 31300 7665 31328
rect 7340 31288 7346 31300
rect 7653 31297 7665 31300
rect 7699 31328 7711 31331
rect 8113 31331 8171 31337
rect 8113 31328 8125 31331
rect 7699 31300 8125 31328
rect 7699 31297 7711 31300
rect 7653 31291 7711 31297
rect 8113 31297 8125 31300
rect 8159 31328 8171 31331
rect 9582 31328 9588 31340
rect 8159 31300 9588 31328
rect 8159 31297 8171 31300
rect 8113 31291 8171 31297
rect 9582 31288 9588 31300
rect 9640 31288 9646 31340
rect 9674 31288 9680 31340
rect 9732 31288 9738 31340
rect 10318 31288 10324 31340
rect 10376 31288 10382 31340
rect 11057 31331 11115 31337
rect 11057 31297 11069 31331
rect 11103 31328 11115 31331
rect 11103 31300 11284 31328
rect 11103 31297 11115 31300
rect 11057 31291 11115 31297
rect 7561 31263 7619 31269
rect 7561 31260 7573 31263
rect 6748 31232 7573 31260
rect 6365 31223 6423 31229
rect 7561 31229 7573 31232
rect 7607 31260 7619 31263
rect 8021 31263 8079 31269
rect 8021 31260 8033 31263
rect 7607 31232 8033 31260
rect 7607 31229 7619 31232
rect 7561 31223 7619 31229
rect 8021 31229 8033 31232
rect 8067 31260 8079 31263
rect 8478 31260 8484 31272
rect 8067 31232 8484 31260
rect 8067 31229 8079 31232
rect 8021 31223 8079 31229
rect 8478 31220 8484 31232
rect 8536 31220 8542 31272
rect 9306 31220 9312 31272
rect 9364 31260 9370 31272
rect 9769 31263 9827 31269
rect 9769 31260 9781 31263
rect 9364 31232 9781 31260
rect 9364 31220 9370 31232
rect 9769 31229 9781 31232
rect 9815 31229 9827 31263
rect 9769 31223 9827 31229
rect 10137 31263 10195 31269
rect 10137 31229 10149 31263
rect 10183 31229 10195 31263
rect 10137 31223 10195 31229
rect 4540 31164 8984 31192
rect 4540 31124 4568 31164
rect 8956 31136 8984 31164
rect 2884 31096 4568 31124
rect 8938 31084 8944 31136
rect 8996 31084 9002 31136
rect 9398 31084 9404 31136
rect 9456 31124 9462 31136
rect 9674 31124 9680 31136
rect 9456 31096 9680 31124
rect 9456 31084 9462 31096
rect 9674 31084 9680 31096
rect 9732 31124 9738 31136
rect 10152 31133 10180 31223
rect 11256 31136 11284 31300
rect 10137 31127 10195 31133
rect 10137 31124 10149 31127
rect 9732 31096 10149 31124
rect 9732 31084 9738 31096
rect 10137 31093 10149 31096
rect 10183 31093 10195 31127
rect 10137 31087 10195 31093
rect 10410 31084 10416 31136
rect 10468 31084 10474 31136
rect 10870 31084 10876 31136
rect 10928 31084 10934 31136
rect 11238 31084 11244 31136
rect 11296 31084 11302 31136
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 1026 30880 1032 30932
rect 1084 30920 1090 30932
rect 1949 30923 2007 30929
rect 1949 30920 1961 30923
rect 1084 30892 1961 30920
rect 1084 30880 1090 30892
rect 1949 30889 1961 30892
rect 1995 30889 2007 30923
rect 1949 30883 2007 30889
rect 3970 30880 3976 30932
rect 4028 30880 4034 30932
rect 4157 30923 4215 30929
rect 4157 30889 4169 30923
rect 4203 30920 4215 30923
rect 4246 30920 4252 30932
rect 4203 30892 4252 30920
rect 4203 30889 4215 30892
rect 4157 30883 4215 30889
rect 4246 30880 4252 30892
rect 4304 30880 4310 30932
rect 4982 30880 4988 30932
rect 5040 30880 5046 30932
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 9217 30923 9275 30929
rect 9217 30920 9229 30923
rect 8536 30892 9229 30920
rect 8536 30880 8542 30892
rect 9217 30889 9229 30892
rect 9263 30889 9275 30923
rect 9217 30883 9275 30889
rect 1946 30784 1952 30796
rect 1688 30756 1952 30784
rect 1688 30725 1716 30756
rect 1946 30744 1952 30756
rect 2004 30784 2010 30796
rect 2409 30787 2467 30793
rect 2409 30784 2421 30787
rect 2004 30756 2421 30784
rect 2004 30744 2010 30756
rect 2409 30753 2421 30756
rect 2455 30784 2467 30787
rect 2498 30784 2504 30796
rect 2455 30756 2504 30784
rect 2455 30753 2467 30756
rect 2409 30747 2467 30753
rect 2498 30744 2504 30756
rect 2556 30744 2562 30796
rect 3988 30784 4016 30880
rect 4264 30852 4292 30880
rect 4341 30855 4399 30861
rect 4341 30852 4353 30855
rect 4264 30824 4353 30852
rect 4341 30821 4353 30824
rect 4387 30821 4399 30855
rect 4798 30852 4804 30864
rect 4341 30815 4399 30821
rect 4724 30824 4804 30852
rect 4724 30793 4752 30824
rect 4798 30812 4804 30824
rect 4856 30812 4862 30864
rect 9232 30852 9260 30883
rect 9232 30824 9444 30852
rect 4709 30787 4767 30793
rect 4709 30784 4721 30787
rect 3988 30756 4721 30784
rect 4709 30753 4721 30756
rect 4755 30753 4767 30787
rect 4709 30747 4767 30753
rect 8481 30787 8539 30793
rect 8481 30753 8493 30787
rect 8527 30784 8539 30787
rect 9306 30784 9312 30796
rect 8527 30756 9312 30784
rect 8527 30753 8539 30756
rect 8481 30747 8539 30753
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 1854 30676 1860 30728
rect 1912 30676 1918 30728
rect 2133 30719 2191 30725
rect 2133 30685 2145 30719
rect 2179 30685 2191 30719
rect 2133 30679 2191 30685
rect 2148 30648 2176 30679
rect 2774 30676 2780 30728
rect 2832 30716 2838 30728
rect 4065 30719 4123 30725
rect 4065 30716 4077 30719
rect 2832 30688 3004 30716
rect 2832 30676 2838 30688
rect 2866 30648 2872 30660
rect 2148 30620 2872 30648
rect 2866 30608 2872 30620
rect 2924 30608 2930 30660
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 1854 30580 1860 30592
rect 1811 30552 1860 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 1854 30540 1860 30552
rect 1912 30540 1918 30592
rect 2777 30583 2835 30589
rect 2777 30549 2789 30583
rect 2823 30580 2835 30583
rect 2976 30580 3004 30688
rect 3436 30688 4077 30716
rect 3436 30592 3464 30688
rect 4065 30685 4077 30688
rect 4111 30685 4123 30719
rect 4065 30679 4123 30685
rect 4338 30676 4344 30728
rect 4396 30676 4402 30728
rect 4798 30676 4804 30728
rect 4856 30676 4862 30728
rect 5718 30676 5724 30728
rect 5776 30716 5782 30728
rect 6825 30719 6883 30725
rect 6825 30716 6837 30719
rect 5776 30688 6837 30716
rect 5776 30676 5782 30688
rect 6825 30685 6837 30688
rect 6871 30685 6883 30719
rect 6825 30679 6883 30685
rect 8662 30676 8668 30728
rect 8720 30676 8726 30728
rect 8938 30676 8944 30728
rect 8996 30676 9002 30728
rect 9140 30725 9168 30756
rect 9306 30744 9312 30756
rect 9364 30744 9370 30796
rect 9416 30728 9444 30824
rect 9950 30812 9956 30864
rect 10008 30852 10014 30864
rect 10045 30855 10103 30861
rect 10045 30852 10057 30855
rect 10008 30824 10057 30852
rect 10008 30812 10014 30824
rect 10045 30821 10057 30824
rect 10091 30852 10103 30855
rect 10410 30852 10416 30864
rect 10091 30824 10416 30852
rect 10091 30821 10103 30824
rect 10045 30815 10103 30821
rect 10410 30812 10416 30824
rect 10468 30852 10474 30864
rect 11977 30855 12035 30861
rect 11977 30852 11989 30855
rect 10468 30824 11989 30852
rect 10468 30812 10474 30824
rect 11977 30821 11989 30824
rect 12023 30852 12035 30855
rect 12066 30852 12072 30864
rect 12023 30824 12072 30852
rect 12023 30821 12035 30824
rect 11977 30815 12035 30821
rect 12066 30812 12072 30824
rect 12124 30812 12130 30864
rect 9582 30744 9588 30796
rect 9640 30744 9646 30796
rect 11149 30787 11207 30793
rect 11149 30784 11161 30787
rect 10704 30756 11161 30784
rect 9125 30719 9183 30725
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 9217 30719 9275 30725
rect 9217 30685 9229 30719
rect 9263 30716 9275 30719
rect 9398 30716 9404 30728
rect 9263 30688 9404 30716
rect 9263 30685 9275 30688
rect 9217 30679 9275 30685
rect 9398 30676 9404 30688
rect 9456 30676 9462 30728
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30716 9735 30719
rect 9858 30716 9864 30728
rect 9723 30688 9864 30716
rect 9723 30685 9735 30688
rect 9677 30679 9735 30685
rect 9858 30676 9864 30688
rect 9916 30676 9922 30728
rect 10226 30676 10232 30728
rect 10284 30676 10290 30728
rect 10594 30676 10600 30728
rect 10652 30716 10658 30728
rect 10704 30725 10732 30756
rect 11149 30753 11161 30756
rect 11195 30753 11207 30787
rect 11149 30747 11207 30753
rect 11238 30744 11244 30796
rect 11296 30784 11302 30796
rect 11296 30756 11652 30784
rect 11296 30744 11302 30756
rect 11624 30725 11652 30756
rect 10689 30719 10747 30725
rect 10689 30716 10701 30719
rect 10652 30688 10701 30716
rect 10652 30676 10658 30688
rect 10689 30685 10701 30688
rect 10735 30685 10747 30719
rect 10689 30679 10747 30685
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30716 11115 30719
rect 11517 30719 11575 30725
rect 11517 30716 11529 30719
rect 11103 30688 11529 30716
rect 11103 30685 11115 30688
rect 11057 30679 11115 30685
rect 11517 30685 11529 30688
rect 11563 30685 11575 30719
rect 11517 30679 11575 30685
rect 11609 30719 11667 30725
rect 11609 30685 11621 30719
rect 11655 30716 11667 30719
rect 11655 30688 12204 30716
rect 11655 30685 11667 30688
rect 11609 30679 11667 30685
rect 3050 30580 3056 30592
rect 2823 30552 3056 30580
rect 2823 30549 2835 30552
rect 2777 30543 2835 30549
rect 3050 30540 3056 30552
rect 3108 30540 3114 30592
rect 3418 30540 3424 30592
rect 3476 30540 3482 30592
rect 4356 30589 4384 30676
rect 4341 30583 4399 30589
rect 4341 30549 4353 30583
rect 4387 30549 4399 30583
rect 4341 30543 4399 30549
rect 7009 30583 7067 30589
rect 7009 30549 7021 30583
rect 7055 30580 7067 30583
rect 8680 30580 8708 30676
rect 9033 30651 9091 30657
rect 9033 30617 9045 30651
rect 9079 30648 9091 30651
rect 9766 30648 9772 30660
rect 9079 30620 9772 30648
rect 9079 30617 9091 30620
rect 9033 30611 9091 30617
rect 9766 30608 9772 30620
rect 9824 30608 9830 30660
rect 10244 30648 10272 30676
rect 10870 30648 10876 30660
rect 10244 30620 10876 30648
rect 10870 30608 10876 30620
rect 10928 30648 10934 30660
rect 11072 30648 11100 30679
rect 10928 30620 11100 30648
rect 10928 30608 10934 30620
rect 12176 30592 12204 30688
rect 7055 30552 8708 30580
rect 7055 30549 7067 30552
rect 7009 30543 7067 30549
rect 10042 30540 10048 30592
rect 10100 30580 10106 30592
rect 10597 30583 10655 30589
rect 10597 30580 10609 30583
rect 10100 30552 10609 30580
rect 10100 30540 10106 30552
rect 10597 30549 10609 30552
rect 10643 30580 10655 30583
rect 10689 30583 10747 30589
rect 10689 30580 10701 30583
rect 10643 30552 10701 30580
rect 10643 30549 10655 30552
rect 10597 30543 10655 30549
rect 10689 30549 10701 30552
rect 10735 30580 10747 30583
rect 11149 30583 11207 30589
rect 11149 30580 11161 30583
rect 10735 30552 11161 30580
rect 10735 30549 10747 30552
rect 10689 30543 10747 30549
rect 11149 30549 11161 30552
rect 11195 30580 11207 30583
rect 11977 30583 12035 30589
rect 11977 30580 11989 30583
rect 11195 30552 11989 30580
rect 11195 30549 11207 30552
rect 11149 30543 11207 30549
rect 11977 30549 11989 30552
rect 12023 30549 12035 30583
rect 11977 30543 12035 30549
rect 12158 30540 12164 30592
rect 12216 30540 12222 30592
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 3050 30336 3056 30388
rect 3108 30376 3114 30388
rect 3605 30379 3663 30385
rect 3605 30376 3617 30379
rect 3108 30348 3617 30376
rect 3108 30336 3114 30348
rect 3605 30345 3617 30348
rect 3651 30345 3663 30379
rect 3605 30339 3663 30345
rect 4433 30379 4491 30385
rect 4433 30345 4445 30379
rect 4479 30376 4491 30379
rect 4798 30376 4804 30388
rect 4479 30348 4804 30376
rect 4479 30345 4491 30348
rect 4433 30339 4491 30345
rect 4798 30336 4804 30348
rect 4856 30336 4862 30388
rect 9398 30336 9404 30388
rect 9456 30376 9462 30388
rect 9493 30379 9551 30385
rect 9493 30376 9505 30379
rect 9456 30348 9505 30376
rect 9456 30336 9462 30348
rect 9493 30345 9505 30348
rect 9539 30376 9551 30379
rect 9953 30379 10011 30385
rect 9953 30376 9965 30379
rect 9539 30348 9965 30376
rect 9539 30345 9551 30348
rect 9493 30339 9551 30345
rect 9953 30345 9965 30348
rect 9999 30376 10011 30379
rect 10042 30376 10048 30388
rect 9999 30348 10048 30376
rect 9999 30345 10011 30348
rect 9953 30339 10011 30345
rect 10042 30336 10048 30348
rect 10100 30376 10106 30388
rect 10413 30379 10471 30385
rect 10413 30376 10425 30379
rect 10100 30348 10425 30376
rect 10100 30336 10106 30348
rect 10413 30345 10425 30348
rect 10459 30376 10471 30379
rect 10686 30376 10692 30388
rect 10459 30348 10692 30376
rect 10459 30345 10471 30348
rect 10413 30339 10471 30345
rect 10686 30336 10692 30348
rect 10744 30376 10750 30388
rect 10873 30379 10931 30385
rect 10873 30376 10885 30379
rect 10744 30348 10885 30376
rect 10744 30336 10750 30348
rect 10873 30345 10885 30348
rect 10919 30376 10931 30379
rect 11333 30379 11391 30385
rect 11333 30376 11345 30379
rect 10919 30348 11345 30376
rect 10919 30345 10931 30348
rect 10873 30339 10931 30345
rect 11333 30345 11345 30348
rect 11379 30376 11391 30379
rect 11977 30379 12035 30385
rect 11977 30376 11989 30379
rect 11379 30348 11989 30376
rect 11379 30345 11391 30348
rect 11333 30339 11391 30345
rect 11977 30345 11989 30348
rect 12023 30376 12035 30379
rect 12069 30379 12127 30385
rect 12069 30376 12081 30379
rect 12023 30348 12081 30376
rect 12023 30345 12035 30348
rect 11977 30339 12035 30345
rect 12069 30345 12081 30348
rect 12115 30376 12127 30379
rect 12529 30379 12587 30385
rect 12529 30376 12541 30379
rect 12115 30348 12541 30376
rect 12115 30345 12127 30348
rect 12069 30339 12127 30345
rect 12529 30345 12541 30348
rect 12575 30345 12587 30379
rect 12529 30339 12587 30345
rect 2685 30311 2743 30317
rect 2685 30277 2697 30311
rect 2731 30308 2743 30311
rect 2731 30280 3924 30308
rect 2731 30277 2743 30280
rect 2685 30271 2743 30277
rect 2777 30243 2835 30249
rect 2777 30209 2789 30243
rect 2823 30240 2835 30243
rect 2823 30212 3004 30240
rect 2823 30209 2835 30212
rect 2777 30203 2835 30209
rect 2976 30184 3004 30212
rect 3896 30184 3924 30280
rect 4062 30268 4068 30320
rect 4120 30268 4126 30320
rect 6825 30311 6883 30317
rect 6825 30277 6837 30311
rect 6871 30308 6883 30311
rect 6871 30280 7236 30308
rect 6871 30277 6883 30280
rect 6825 30271 6883 30277
rect 7208 30252 7236 30280
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7009 30243 7067 30249
rect 7009 30240 7021 30243
rect 6972 30212 7021 30240
rect 6972 30200 6978 30212
rect 7009 30209 7021 30212
rect 7055 30209 7067 30243
rect 7009 30203 7067 30209
rect 7190 30200 7196 30252
rect 7248 30200 7254 30252
rect 9493 30243 9551 30249
rect 9493 30209 9505 30243
rect 9539 30240 9551 30243
rect 9950 30240 9956 30252
rect 9539 30212 9956 30240
rect 9539 30209 9551 30212
rect 9493 30203 9551 30209
rect 9950 30200 9956 30212
rect 10008 30200 10014 30252
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30240 10471 30243
rect 10594 30240 10600 30252
rect 10459 30212 10600 30240
rect 10459 30209 10471 30212
rect 10413 30203 10471 30209
rect 10594 30200 10600 30212
rect 10652 30240 10658 30252
rect 10873 30243 10931 30249
rect 10873 30240 10885 30243
rect 10652 30212 10885 30240
rect 10652 30200 10658 30212
rect 10873 30209 10885 30212
rect 10919 30240 10931 30243
rect 11333 30243 11391 30249
rect 11333 30240 11345 30243
rect 10919 30212 11345 30240
rect 10919 30209 10931 30212
rect 10873 30203 10931 30209
rect 11333 30209 11345 30212
rect 11379 30240 11391 30243
rect 11977 30243 12035 30249
rect 11977 30240 11989 30243
rect 11379 30212 11989 30240
rect 11379 30209 11391 30212
rect 11333 30203 11391 30209
rect 11977 30209 11989 30212
rect 12023 30240 12035 30243
rect 12529 30243 12587 30249
rect 12529 30240 12541 30243
rect 12023 30212 12541 30240
rect 12023 30209 12035 30212
rect 11977 30203 12035 30209
rect 12529 30209 12541 30212
rect 12575 30209 12587 30243
rect 12529 30203 12587 30209
rect 15838 30200 15844 30252
rect 15896 30200 15902 30252
rect 1946 30132 1952 30184
rect 2004 30132 2010 30184
rect 2225 30175 2283 30181
rect 2225 30141 2237 30175
rect 2271 30172 2283 30175
rect 2869 30175 2927 30181
rect 2271 30144 2360 30172
rect 2271 30141 2283 30144
rect 2225 30135 2283 30141
rect 2332 30113 2360 30144
rect 2869 30141 2881 30175
rect 2915 30141 2927 30175
rect 2869 30135 2927 30141
rect 2317 30107 2375 30113
rect 2317 30073 2329 30107
rect 2363 30073 2375 30107
rect 2884 30104 2912 30135
rect 2958 30132 2964 30184
rect 3016 30132 3022 30184
rect 3234 30132 3240 30184
rect 3292 30132 3298 30184
rect 3418 30132 3424 30184
rect 3476 30172 3482 30184
rect 3789 30175 3847 30181
rect 3789 30172 3801 30175
rect 3476 30144 3801 30172
rect 3476 30132 3482 30144
rect 3789 30141 3801 30144
rect 3835 30141 3847 30175
rect 3789 30135 3847 30141
rect 3878 30132 3884 30184
rect 3936 30172 3942 30184
rect 3973 30175 4031 30181
rect 3973 30172 3985 30175
rect 3936 30144 3985 30172
rect 3936 30132 3942 30144
rect 3973 30141 3985 30144
rect 4019 30141 4031 30175
rect 3973 30135 4031 30141
rect 4525 30175 4583 30181
rect 4525 30141 4537 30175
rect 4571 30141 4583 30175
rect 4525 30135 4583 30141
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 9585 30175 9643 30181
rect 9585 30172 9597 30175
rect 9171 30144 9597 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 9585 30141 9597 30144
rect 9631 30172 9643 30175
rect 9858 30172 9864 30184
rect 9631 30144 9864 30172
rect 9631 30141 9643 30144
rect 9585 30135 9643 30141
rect 2317 30067 2375 30073
rect 2746 30076 2912 30104
rect 3605 30107 3663 30113
rect 2746 30048 2774 30076
rect 3605 30073 3617 30107
rect 3651 30104 3663 30107
rect 4540 30104 4568 30135
rect 9858 30132 9864 30144
rect 9916 30132 9922 30184
rect 10045 30175 10103 30181
rect 10045 30141 10057 30175
rect 10091 30172 10103 30175
rect 10226 30172 10232 30184
rect 10091 30144 10232 30172
rect 10091 30141 10103 30144
rect 10045 30135 10103 30141
rect 10226 30132 10232 30144
rect 10284 30172 10290 30184
rect 10505 30175 10563 30181
rect 10505 30172 10517 30175
rect 10284 30144 10517 30172
rect 10284 30132 10290 30144
rect 10505 30141 10517 30144
rect 10551 30172 10563 30175
rect 10962 30172 10968 30184
rect 10551 30144 10968 30172
rect 10551 30141 10563 30144
rect 10505 30135 10563 30141
rect 10962 30132 10968 30144
rect 11020 30172 11026 30184
rect 11609 30175 11667 30181
rect 11609 30172 11621 30175
rect 11020 30144 11621 30172
rect 11020 30132 11026 30144
rect 11609 30141 11621 30144
rect 11655 30141 11667 30175
rect 11609 30135 11667 30141
rect 3651 30076 4568 30104
rect 11624 30104 11652 30135
rect 12066 30132 12072 30184
rect 12124 30132 12130 30184
rect 12158 30132 12164 30184
rect 12216 30172 12222 30184
rect 12437 30175 12495 30181
rect 12437 30172 12449 30175
rect 12216 30144 12449 30172
rect 12216 30132 12222 30144
rect 12437 30141 12449 30144
rect 12483 30141 12495 30175
rect 12437 30135 12495 30141
rect 12897 30175 12955 30181
rect 12897 30141 12909 30175
rect 12943 30141 12955 30175
rect 12897 30135 12955 30141
rect 12912 30104 12940 30135
rect 11624 30076 12940 30104
rect 3651 30073 3663 30076
rect 3605 30067 3663 30073
rect 2682 29996 2688 30048
rect 2740 30008 2774 30048
rect 2740 29996 2746 30008
rect 6638 29996 6644 30048
rect 6696 29996 6702 30048
rect 15654 29996 15660 30048
rect 15712 29996 15718 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 3234 29792 3240 29844
rect 3292 29832 3298 29844
rect 3421 29835 3479 29841
rect 3421 29832 3433 29835
rect 3292 29804 3433 29832
rect 3292 29792 3298 29804
rect 3421 29801 3433 29804
rect 3467 29801 3479 29835
rect 3421 29795 3479 29801
rect 4798 29792 4804 29844
rect 4856 29832 4862 29844
rect 10137 29835 10195 29841
rect 4856 29804 10088 29832
rect 4856 29792 4862 29804
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 1854 29696 1860 29708
rect 1443 29668 1860 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 1854 29656 1860 29668
rect 1912 29696 1918 29708
rect 2130 29696 2136 29708
rect 1912 29668 2136 29696
rect 1912 29656 1918 29668
rect 2130 29656 2136 29668
rect 2188 29696 2194 29708
rect 2317 29699 2375 29705
rect 2317 29696 2329 29699
rect 2188 29668 2329 29696
rect 2188 29656 2194 29668
rect 2317 29665 2329 29668
rect 2363 29665 2375 29699
rect 2317 29659 2375 29665
rect 1762 29588 1768 29640
rect 1820 29628 1826 29640
rect 2225 29631 2283 29637
rect 2225 29628 2237 29631
rect 1820 29600 2237 29628
rect 1820 29588 1826 29600
rect 2225 29597 2237 29600
rect 2271 29628 2283 29631
rect 2682 29628 2688 29640
rect 2271 29600 2688 29628
rect 2271 29597 2283 29600
rect 2225 29591 2283 29597
rect 2682 29588 2688 29600
rect 2740 29588 2746 29640
rect 3513 29631 3571 29637
rect 3513 29597 3525 29631
rect 3559 29597 3571 29631
rect 3513 29591 3571 29597
rect 3528 29504 3556 29591
rect 4246 29588 4252 29640
rect 4304 29628 4310 29640
rect 4433 29631 4491 29637
rect 4433 29628 4445 29631
rect 4304 29600 4445 29628
rect 4304 29588 4310 29600
rect 4433 29597 4445 29600
rect 4479 29628 4491 29631
rect 5905 29631 5963 29637
rect 5905 29628 5917 29631
rect 4479 29600 5917 29628
rect 4479 29597 4491 29600
rect 4433 29591 4491 29597
rect 5905 29597 5917 29600
rect 5951 29628 5963 29631
rect 7377 29631 7435 29637
rect 7377 29628 7389 29631
rect 5951 29600 7389 29628
rect 5951 29597 5963 29600
rect 5905 29591 5963 29597
rect 7377 29597 7389 29600
rect 7423 29597 7435 29631
rect 7377 29591 7435 29597
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29597 9551 29631
rect 9493 29591 9551 29597
rect 4700 29563 4758 29569
rect 4700 29529 4712 29563
rect 4746 29560 4758 29563
rect 5074 29560 5080 29572
rect 4746 29532 5080 29560
rect 4746 29529 4758 29532
rect 4700 29523 4758 29529
rect 5074 29520 5080 29532
rect 5132 29520 5138 29572
rect 6172 29563 6230 29569
rect 6172 29529 6184 29563
rect 6218 29560 6230 29563
rect 6362 29560 6368 29572
rect 6218 29532 6368 29560
rect 6218 29529 6230 29532
rect 6172 29523 6230 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 7650 29569 7656 29572
rect 7644 29523 7656 29569
rect 7650 29520 7656 29523
rect 7708 29520 7714 29572
rect 8294 29520 8300 29572
rect 8352 29560 8358 29572
rect 8941 29563 8999 29569
rect 8941 29560 8953 29563
rect 8352 29532 8953 29560
rect 8352 29520 8358 29532
rect 8941 29529 8953 29532
rect 8987 29529 8999 29563
rect 8941 29523 8999 29529
rect 1765 29495 1823 29501
rect 1765 29461 1777 29495
rect 1811 29492 1823 29495
rect 1854 29492 1860 29504
rect 1811 29464 1860 29492
rect 1811 29461 1823 29464
rect 1765 29455 1823 29461
rect 1854 29452 1860 29464
rect 1912 29492 1918 29504
rect 2225 29495 2283 29501
rect 2225 29492 2237 29495
rect 1912 29464 2237 29492
rect 1912 29452 1918 29464
rect 2225 29461 2237 29464
rect 2271 29492 2283 29495
rect 2685 29495 2743 29501
rect 2685 29492 2697 29495
rect 2271 29464 2697 29492
rect 2271 29461 2283 29464
rect 2225 29455 2283 29461
rect 2685 29461 2697 29464
rect 2731 29492 2743 29495
rect 3050 29492 3056 29504
rect 2731 29464 3056 29492
rect 2731 29461 2743 29464
rect 2685 29455 2743 29461
rect 3050 29452 3056 29464
rect 3108 29452 3114 29504
rect 3510 29452 3516 29504
rect 3568 29452 3574 29504
rect 5813 29495 5871 29501
rect 5813 29461 5825 29495
rect 5859 29492 5871 29495
rect 5994 29492 6000 29504
rect 5859 29464 6000 29492
rect 5859 29461 5871 29464
rect 5813 29455 5871 29461
rect 5994 29452 6000 29464
rect 6052 29452 6058 29504
rect 7190 29452 7196 29504
rect 7248 29492 7254 29504
rect 7285 29495 7343 29501
rect 7285 29492 7297 29495
rect 7248 29464 7297 29492
rect 7248 29452 7254 29464
rect 7285 29461 7297 29464
rect 7331 29461 7343 29495
rect 7285 29455 7343 29461
rect 7558 29452 7564 29504
rect 7616 29492 7622 29504
rect 8757 29495 8815 29501
rect 8757 29492 8769 29495
rect 7616 29464 8769 29492
rect 7616 29452 7622 29464
rect 8757 29461 8769 29464
rect 8803 29492 8815 29495
rect 9508 29492 9536 29591
rect 9766 29588 9772 29640
rect 9824 29588 9830 29640
rect 10060 29637 10088 29804
rect 10137 29801 10149 29835
rect 10183 29832 10195 29835
rect 10318 29832 10324 29844
rect 10183 29804 10324 29832
rect 10183 29801 10195 29804
rect 10137 29795 10195 29801
rect 10318 29792 10324 29804
rect 10376 29792 10382 29844
rect 12066 29792 12072 29844
rect 12124 29792 12130 29844
rect 12158 29792 12164 29844
rect 12216 29792 12222 29844
rect 15838 29792 15844 29844
rect 15896 29832 15902 29844
rect 16117 29835 16175 29841
rect 16117 29832 16129 29835
rect 15896 29804 16129 29832
rect 15896 29792 15902 29804
rect 16117 29801 16129 29804
rect 16163 29801 16175 29835
rect 16117 29795 16175 29801
rect 10594 29724 10600 29776
rect 10652 29764 10658 29776
rect 11057 29767 11115 29773
rect 11057 29764 11069 29767
rect 10652 29736 11069 29764
rect 10652 29724 10658 29736
rect 11057 29733 11069 29736
rect 11103 29764 11115 29767
rect 11146 29764 11152 29776
rect 11103 29736 11152 29764
rect 11103 29733 11115 29736
rect 11057 29727 11115 29733
rect 11146 29724 11152 29736
rect 11204 29724 11210 29776
rect 11885 29767 11943 29773
rect 11885 29733 11897 29767
rect 11931 29764 11943 29767
rect 12084 29764 12112 29792
rect 11931 29736 12112 29764
rect 11931 29733 11943 29736
rect 11885 29727 11943 29733
rect 10962 29656 10968 29708
rect 11020 29696 11026 29708
rect 11425 29699 11483 29705
rect 11425 29696 11437 29699
rect 11020 29668 11437 29696
rect 11020 29656 11026 29668
rect 11425 29665 11437 29668
rect 11471 29665 11483 29699
rect 11425 29659 11483 29665
rect 11517 29699 11575 29705
rect 11517 29665 11529 29699
rect 11563 29696 11575 29699
rect 12176 29696 12204 29792
rect 14277 29767 14335 29773
rect 14277 29733 14289 29767
rect 14323 29733 14335 29767
rect 14277 29727 14335 29733
rect 11563 29668 12204 29696
rect 14292 29696 14320 29727
rect 14642 29724 14648 29776
rect 14700 29724 14706 29776
rect 15746 29724 15752 29776
rect 15804 29764 15810 29776
rect 16209 29767 16267 29773
rect 16209 29764 16221 29767
rect 15804 29736 16221 29764
rect 15804 29724 15810 29736
rect 16209 29733 16221 29736
rect 16255 29764 16267 29767
rect 16853 29767 16911 29773
rect 16853 29764 16865 29767
rect 16255 29736 16865 29764
rect 16255 29733 16267 29736
rect 16209 29727 16267 29733
rect 16853 29733 16865 29736
rect 16899 29733 16911 29767
rect 16853 29727 16911 29733
rect 14660 29696 14688 29724
rect 14292 29668 14780 29696
rect 11563 29665 11575 29668
rect 11517 29659 11575 29665
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29597 10103 29631
rect 10045 29591 10103 29597
rect 9858 29520 9864 29572
rect 9916 29560 9922 29572
rect 9953 29563 10011 29569
rect 9953 29560 9965 29563
rect 9916 29532 9965 29560
rect 9916 29520 9922 29532
rect 9953 29529 9965 29532
rect 9999 29560 10011 29563
rect 11532 29560 11560 29659
rect 14458 29588 14464 29640
rect 14516 29628 14522 29640
rect 14645 29631 14703 29637
rect 14645 29628 14657 29631
rect 14516 29600 14657 29628
rect 14516 29588 14522 29600
rect 14645 29597 14657 29600
rect 14691 29597 14703 29631
rect 14752 29628 14780 29668
rect 18233 29631 18291 29637
rect 14752 29600 16160 29628
rect 14645 29591 14703 29597
rect 9999 29532 11560 29560
rect 9999 29529 10011 29532
rect 9953 29523 10011 29529
rect 14366 29520 14372 29572
rect 14424 29560 14430 29572
rect 14553 29563 14611 29569
rect 14553 29560 14565 29563
rect 14424 29532 14565 29560
rect 14424 29520 14430 29532
rect 14553 29529 14565 29532
rect 14599 29529 14611 29563
rect 14553 29523 14611 29529
rect 14734 29520 14740 29572
rect 14792 29560 14798 29572
rect 14890 29563 14948 29569
rect 14890 29560 14902 29563
rect 14792 29532 14902 29560
rect 14792 29520 14798 29532
rect 14890 29529 14902 29532
rect 14936 29529 14948 29563
rect 14890 29523 14948 29529
rect 8803 29464 9536 29492
rect 10597 29495 10655 29501
rect 8803 29461 8815 29464
rect 8757 29455 8815 29461
rect 10597 29461 10609 29495
rect 10643 29492 10655 29495
rect 10686 29492 10692 29504
rect 10643 29464 10692 29492
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 10686 29452 10692 29464
rect 10744 29492 10750 29504
rect 11057 29495 11115 29501
rect 11057 29492 11069 29495
rect 10744 29464 11069 29492
rect 10744 29452 10750 29464
rect 11057 29461 11069 29464
rect 11103 29492 11115 29495
rect 11885 29495 11943 29501
rect 11885 29492 11897 29495
rect 11103 29464 11897 29492
rect 11103 29461 11115 29464
rect 11057 29455 11115 29461
rect 11885 29461 11897 29464
rect 11931 29461 11943 29495
rect 11885 29455 11943 29461
rect 14090 29452 14096 29504
rect 14148 29452 14154 29504
rect 15470 29452 15476 29504
rect 15528 29492 15534 29504
rect 16025 29495 16083 29501
rect 16025 29492 16037 29495
rect 15528 29464 16037 29492
rect 15528 29452 15534 29464
rect 16025 29461 16037 29464
rect 16071 29461 16083 29495
rect 16132 29492 16160 29600
rect 18233 29597 18245 29631
rect 18279 29628 18291 29631
rect 18782 29628 18788 29640
rect 18279 29600 18788 29628
rect 18279 29597 18291 29600
rect 18233 29591 18291 29597
rect 18782 29588 18788 29600
rect 18840 29588 18846 29640
rect 16482 29520 16488 29572
rect 16540 29560 16546 29572
rect 16577 29563 16635 29569
rect 16577 29560 16589 29563
rect 16540 29532 16589 29560
rect 16540 29520 16546 29532
rect 16577 29529 16589 29532
rect 16623 29529 16635 29563
rect 16577 29523 16635 29529
rect 17954 29520 17960 29572
rect 18012 29569 18018 29572
rect 18012 29523 18024 29569
rect 18012 29520 18018 29523
rect 20806 29492 20812 29504
rect 16132 29464 20812 29492
rect 16025 29455 16083 29461
rect 20806 29452 20812 29464
rect 20864 29452 20870 29504
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 1854 29248 1860 29300
rect 1912 29248 1918 29300
rect 3050 29248 3056 29300
rect 3108 29288 3114 29300
rect 3237 29291 3295 29297
rect 3237 29288 3249 29291
rect 3108 29260 3249 29288
rect 3108 29248 3114 29260
rect 3237 29257 3249 29260
rect 3283 29257 3295 29291
rect 3237 29251 3295 29257
rect 5074 29248 5080 29300
rect 5132 29248 5138 29300
rect 6089 29291 6147 29297
rect 6089 29288 6101 29291
rect 5276 29260 6101 29288
rect 3510 29220 3516 29232
rect 2976 29192 3516 29220
rect 2976 29164 3004 29192
rect 3510 29180 3516 29192
rect 3568 29220 3574 29232
rect 4062 29220 4068 29232
rect 3568 29192 4068 29220
rect 3568 29180 3574 29192
rect 4062 29180 4068 29192
rect 4120 29220 4126 29232
rect 4249 29223 4307 29229
rect 4249 29220 4261 29223
rect 4120 29192 4261 29220
rect 4120 29180 4126 29192
rect 4249 29189 4261 29192
rect 4295 29189 4307 29223
rect 4249 29183 4307 29189
rect 2130 29112 2136 29164
rect 2188 29152 2194 29164
rect 2225 29155 2283 29161
rect 2225 29152 2237 29155
rect 2188 29124 2237 29152
rect 2188 29112 2194 29124
rect 2225 29121 2237 29124
rect 2271 29121 2283 29155
rect 2225 29115 2283 29121
rect 2958 29112 2964 29164
rect 3016 29112 3022 29164
rect 3234 29112 3240 29164
rect 3292 29152 3298 29164
rect 3878 29152 3884 29164
rect 3292 29124 3884 29152
rect 3292 29112 3298 29124
rect 3878 29112 3884 29124
rect 3936 29152 3942 29164
rect 4157 29155 4215 29161
rect 4157 29152 4169 29155
rect 3936 29124 4169 29152
rect 3936 29112 3942 29124
rect 4157 29121 4169 29124
rect 4203 29121 4215 29155
rect 4157 29115 4215 29121
rect 5166 29112 5172 29164
rect 5224 29112 5230 29164
rect 5276 29152 5304 29260
rect 6089 29257 6101 29260
rect 6135 29288 6147 29291
rect 6914 29288 6920 29300
rect 6135 29260 6920 29288
rect 6135 29257 6147 29260
rect 6089 29251 6147 29257
rect 6914 29248 6920 29260
rect 6972 29288 6978 29300
rect 8037 29291 8095 29297
rect 8037 29288 8049 29291
rect 6972 29260 8049 29288
rect 6972 29248 6978 29260
rect 8037 29257 8049 29260
rect 8083 29257 8095 29291
rect 8037 29251 8095 29257
rect 11146 29248 11152 29300
rect 11204 29248 11210 29300
rect 12066 29248 12072 29300
rect 12124 29248 12130 29300
rect 14458 29248 14464 29300
rect 14516 29248 14522 29300
rect 15654 29248 15660 29300
rect 15712 29248 15718 29300
rect 20806 29248 20812 29300
rect 20864 29248 20870 29300
rect 5442 29180 5448 29232
rect 5500 29220 5506 29232
rect 7837 29223 7895 29229
rect 7837 29220 7849 29223
rect 5500 29192 5672 29220
rect 5500 29180 5506 29192
rect 5644 29161 5672 29192
rect 7208 29192 7849 29220
rect 5353 29155 5411 29161
rect 5353 29152 5365 29155
rect 5276 29124 5365 29152
rect 5353 29121 5365 29124
rect 5399 29121 5411 29155
rect 5353 29115 5411 29121
rect 5629 29155 5687 29161
rect 5629 29121 5641 29155
rect 5675 29121 5687 29155
rect 5629 29115 5687 29121
rect 5813 29155 5871 29161
rect 5813 29121 5825 29155
rect 5859 29152 5871 29155
rect 5905 29155 5963 29161
rect 5905 29152 5917 29155
rect 5859 29124 5917 29152
rect 5859 29121 5871 29124
rect 5813 29115 5871 29121
rect 5905 29121 5917 29124
rect 5951 29121 5963 29155
rect 5905 29115 5963 29121
rect 7208 29096 7236 29192
rect 7837 29189 7849 29192
rect 7883 29189 7895 29223
rect 7837 29183 7895 29189
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 10146 29155 10204 29161
rect 10146 29152 10158 29155
rect 9732 29124 10158 29152
rect 9732 29112 9738 29124
rect 10146 29121 10158 29124
rect 10192 29121 10204 29155
rect 10146 29115 10204 29121
rect 10318 29112 10324 29164
rect 10376 29152 10382 29164
rect 10413 29155 10471 29161
rect 10413 29152 10425 29155
rect 10376 29124 10425 29152
rect 10376 29112 10382 29124
rect 10413 29121 10425 29124
rect 10459 29121 10471 29155
rect 10413 29115 10471 29121
rect 11333 29155 11391 29161
rect 11333 29121 11345 29155
rect 11379 29152 11391 29155
rect 12084 29152 12112 29248
rect 14476 29220 14504 29248
rect 13280 29192 14504 29220
rect 11379 29124 12112 29152
rect 11379 29121 11391 29124
rect 11333 29115 11391 29121
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 13280 29161 13308 29192
rect 13538 29161 13544 29164
rect 13265 29155 13323 29161
rect 13265 29152 13277 29155
rect 12492 29124 13277 29152
rect 12492 29112 12498 29124
rect 13265 29121 13277 29124
rect 13311 29121 13323 29155
rect 13265 29115 13323 29121
rect 13532 29115 13544 29161
rect 13538 29112 13544 29115
rect 13596 29112 13602 29164
rect 14476 29152 14504 29192
rect 15188 29223 15246 29229
rect 15188 29189 15200 29223
rect 15234 29220 15246 29223
rect 15672 29220 15700 29248
rect 15234 29192 15700 29220
rect 15234 29189 15246 29192
rect 15188 29183 15246 29189
rect 16482 29180 16488 29232
rect 16540 29220 16546 29232
rect 17681 29223 17739 29229
rect 17681 29220 17693 29223
rect 16540 29192 17693 29220
rect 16540 29180 16546 29192
rect 17681 29189 17693 29192
rect 17727 29189 17739 29223
rect 17681 29183 17739 29189
rect 14921 29155 14979 29161
rect 14921 29152 14933 29155
rect 14476 29124 14933 29152
rect 14921 29121 14933 29124
rect 14967 29121 14979 29155
rect 14921 29115 14979 29121
rect 15470 29112 15476 29164
rect 15528 29152 15534 29164
rect 18046 29161 18052 29164
rect 15528 29124 16988 29152
rect 15528 29112 15534 29124
rect 2774 29044 2780 29096
rect 2832 29084 2838 29096
rect 2869 29087 2927 29093
rect 2869 29084 2881 29087
rect 2832 29056 2881 29084
rect 2832 29044 2838 29056
rect 2869 29053 2881 29056
rect 2915 29053 2927 29087
rect 2869 29047 2927 29053
rect 4065 29087 4123 29093
rect 4065 29053 4077 29087
rect 4111 29084 4123 29087
rect 4338 29084 4344 29096
rect 4111 29056 4344 29084
rect 4111 29053 4123 29056
rect 4065 29047 4123 29053
rect 4338 29044 4344 29056
rect 4396 29084 4402 29096
rect 4798 29084 4804 29096
rect 4396 29056 4804 29084
rect 4396 29044 4402 29056
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 4982 29084 4988 29096
rect 4908 29056 4988 29084
rect 1854 28976 1860 29028
rect 1912 28976 1918 29028
rect 3050 28976 3056 29028
rect 3108 29016 3114 29028
rect 4908 29025 4936 29056
rect 4982 29044 4988 29056
rect 5040 29044 5046 29096
rect 5445 29087 5503 29093
rect 5445 29053 5457 29087
rect 5491 29084 5503 29087
rect 5994 29084 6000 29096
rect 5491 29056 6000 29084
rect 5491 29053 5503 29056
rect 5445 29047 5503 29053
rect 5994 29044 6000 29056
rect 6052 29084 6058 29096
rect 6917 29087 6975 29093
rect 6917 29084 6929 29087
rect 6052 29056 6929 29084
rect 6052 29044 6058 29056
rect 6917 29053 6929 29056
rect 6963 29053 6975 29087
rect 6917 29047 6975 29053
rect 7190 29044 7196 29096
rect 7248 29044 7254 29096
rect 8386 29044 8392 29096
rect 8444 29084 8450 29096
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 8444 29056 9076 29084
rect 8444 29044 8450 29056
rect 3237 29019 3295 29025
rect 3237 29016 3249 29019
rect 3108 28988 3249 29016
rect 3108 28976 3114 28988
rect 3237 28985 3249 28988
rect 3283 28985 3295 29019
rect 3237 28979 3295 28985
rect 4617 29019 4675 29025
rect 4617 28985 4629 29019
rect 4663 29016 4675 29019
rect 4893 29019 4951 29025
rect 4663 28988 4844 29016
rect 4663 28985 4675 28988
rect 4617 28979 4675 28985
rect 4816 28948 4844 28988
rect 4893 28985 4905 29019
rect 4939 28985 4951 29019
rect 5718 29016 5724 29028
rect 4893 28979 4951 28985
rect 5000 28988 5724 29016
rect 5000 28948 5028 28988
rect 5718 28976 5724 28988
rect 5776 28976 5782 29028
rect 9048 29025 9076 29056
rect 16500 29056 16681 29084
rect 9033 29019 9091 29025
rect 7576 28988 8064 29016
rect 7576 28960 7604 28988
rect 4816 28920 5028 28948
rect 6178 28908 6184 28960
rect 6236 28948 6242 28960
rect 6365 28951 6423 28957
rect 6365 28948 6377 28951
rect 6236 28920 6377 28948
rect 6236 28908 6242 28920
rect 6365 28917 6377 28920
rect 6411 28917 6423 28951
rect 6365 28911 6423 28917
rect 7558 28908 7564 28960
rect 7616 28908 7622 28960
rect 7742 28908 7748 28960
rect 7800 28908 7806 28960
rect 8036 28957 8064 28988
rect 9033 28985 9045 29019
rect 9079 28985 9091 29019
rect 9033 28979 9091 28985
rect 16298 28976 16304 29028
rect 16356 28976 16362 29028
rect 16500 28960 16528 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16669 29047 16727 29053
rect 16960 29025 16988 29124
rect 18040 29115 18052 29161
rect 18046 29112 18052 29115
rect 18104 29112 18110 29164
rect 19702 29161 19708 29164
rect 19696 29115 19708 29161
rect 19702 29112 19708 29115
rect 19760 29112 19766 29164
rect 17773 29087 17831 29093
rect 17773 29053 17785 29087
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 19429 29087 19487 29093
rect 19429 29053 19441 29087
rect 19475 29053 19487 29087
rect 19429 29047 19487 29053
rect 16945 29019 17003 29025
rect 16945 28985 16957 29019
rect 16991 28985 17003 29019
rect 16945 28979 17003 28985
rect 17402 28976 17408 29028
rect 17460 28976 17466 29028
rect 8021 28951 8079 28957
rect 8021 28917 8033 28951
rect 8067 28917 8079 28951
rect 8021 28911 8079 28917
rect 8205 28951 8263 28957
rect 8205 28917 8217 28951
rect 8251 28948 8263 28951
rect 8478 28948 8484 28960
rect 8251 28920 8484 28948
rect 8251 28917 8263 28920
rect 8205 28911 8263 28917
rect 8478 28908 8484 28920
rect 8536 28908 8542 28960
rect 8846 28908 8852 28960
rect 8904 28948 8910 28960
rect 8941 28951 8999 28957
rect 8941 28948 8953 28951
rect 8904 28920 8953 28948
rect 8904 28908 8910 28920
rect 8941 28917 8953 28920
rect 8987 28917 8999 28951
rect 8941 28911 8999 28917
rect 14550 28908 14556 28960
rect 14608 28948 14614 28960
rect 14645 28951 14703 28957
rect 14645 28948 14657 28951
rect 14608 28920 14657 28948
rect 14608 28908 14614 28920
rect 14645 28917 14657 28920
rect 14691 28917 14703 28951
rect 14645 28911 14703 28917
rect 15286 28908 15292 28960
rect 15344 28948 15350 28960
rect 16482 28948 16488 28960
rect 15344 28920 16488 28948
rect 15344 28908 15350 28920
rect 16482 28908 16488 28920
rect 16540 28908 16546 28960
rect 17126 28908 17132 28960
rect 17184 28908 17190 28960
rect 17218 28908 17224 28960
rect 17276 28908 17282 28960
rect 17788 28948 17816 29047
rect 19058 28976 19064 29028
rect 19116 29016 19122 29028
rect 19153 29019 19211 29025
rect 19153 29016 19165 29019
rect 19116 28988 19165 29016
rect 19116 28976 19122 28988
rect 19153 28985 19165 28988
rect 19199 28985 19211 29019
rect 19153 28979 19211 28985
rect 18874 28948 18880 28960
rect 17788 28920 18880 28948
rect 18874 28908 18880 28920
rect 18932 28948 18938 28960
rect 19444 28948 19472 29047
rect 18932 28920 19472 28948
rect 18932 28908 18938 28920
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 1578 28704 1584 28756
rect 1636 28704 1642 28756
rect 2317 28747 2375 28753
rect 2317 28713 2329 28747
rect 2363 28744 2375 28747
rect 2774 28744 2780 28756
rect 2363 28716 2780 28744
rect 2363 28713 2375 28716
rect 2317 28707 2375 28713
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 2038 28500 2044 28552
rect 2096 28500 2102 28552
rect 2225 28543 2283 28549
rect 2225 28509 2237 28543
rect 2271 28540 2283 28543
rect 2332 28540 2360 28707
rect 2774 28704 2780 28716
rect 2832 28704 2838 28756
rect 5166 28704 5172 28756
rect 5224 28744 5230 28756
rect 5261 28747 5319 28753
rect 5261 28744 5273 28747
rect 5224 28716 5273 28744
rect 5224 28704 5230 28716
rect 5261 28713 5273 28716
rect 5307 28713 5319 28747
rect 5261 28707 5319 28713
rect 6362 28704 6368 28756
rect 6420 28704 6426 28756
rect 7650 28704 7656 28756
rect 7708 28744 7714 28756
rect 7745 28747 7803 28753
rect 7745 28744 7757 28747
rect 7708 28716 7757 28744
rect 7708 28704 7714 28716
rect 7745 28713 7757 28716
rect 7791 28713 7803 28747
rect 7745 28707 7803 28713
rect 9125 28747 9183 28753
rect 9125 28713 9137 28747
rect 9171 28744 9183 28747
rect 9674 28744 9680 28756
rect 9171 28716 9680 28744
rect 9171 28713 9183 28716
rect 9125 28707 9183 28713
rect 9674 28704 9680 28716
rect 9732 28704 9738 28756
rect 13538 28704 13544 28756
rect 13596 28744 13602 28756
rect 13633 28747 13691 28753
rect 13633 28744 13645 28747
rect 13596 28716 13645 28744
rect 13596 28704 13602 28716
rect 13633 28713 13645 28716
rect 13679 28713 13691 28747
rect 14366 28744 14372 28756
rect 13633 28707 13691 28713
rect 14200 28716 14372 28744
rect 5442 28636 5448 28688
rect 5500 28636 5506 28688
rect 7377 28679 7435 28685
rect 7377 28645 7389 28679
rect 7423 28645 7435 28679
rect 9493 28679 9551 28685
rect 9493 28676 9505 28679
rect 7377 28639 7435 28645
rect 9232 28648 9505 28676
rect 3237 28611 3295 28617
rect 3237 28577 3249 28611
rect 3283 28608 3295 28611
rect 5460 28608 5488 28636
rect 3283 28580 3464 28608
rect 3283 28577 3295 28580
rect 3237 28571 3295 28577
rect 3436 28549 3464 28580
rect 5276 28580 5488 28608
rect 7392 28608 7420 28639
rect 8665 28611 8723 28617
rect 7392 28580 7788 28608
rect 5276 28549 5304 28580
rect 2271 28512 2360 28540
rect 2501 28543 2559 28549
rect 2271 28509 2283 28512
rect 2225 28503 2283 28509
rect 2501 28509 2513 28543
rect 2547 28540 2559 28543
rect 3421 28543 3479 28549
rect 2547 28512 2636 28540
rect 2547 28509 2559 28512
rect 2501 28503 2559 28509
rect 2130 28364 2136 28416
rect 2188 28364 2194 28416
rect 2608 28413 2636 28512
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 5261 28543 5319 28549
rect 3467 28512 3832 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3804 28416 3832 28512
rect 5261 28509 5273 28543
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 5445 28543 5503 28549
rect 5445 28509 5457 28543
rect 5491 28509 5503 28543
rect 5445 28503 5503 28509
rect 5460 28472 5488 28503
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5629 28543 5687 28549
rect 5629 28540 5641 28543
rect 5592 28512 5641 28540
rect 5592 28500 5598 28512
rect 5629 28509 5641 28512
rect 5675 28509 5687 28543
rect 5629 28503 5687 28509
rect 6178 28500 6184 28552
rect 6236 28500 6242 28552
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 6638 28500 6644 28552
rect 6696 28540 6702 28552
rect 6825 28543 6883 28549
rect 6825 28540 6837 28543
rect 6696 28512 6837 28540
rect 6696 28500 6702 28512
rect 6825 28509 6837 28512
rect 6871 28509 6883 28543
rect 6825 28503 6883 28509
rect 6914 28500 6920 28552
rect 6972 28540 6978 28552
rect 7101 28543 7159 28549
rect 7101 28540 7113 28543
rect 6972 28512 7113 28540
rect 6972 28500 6978 28512
rect 7101 28509 7113 28512
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 7466 28500 7472 28552
rect 7524 28500 7530 28552
rect 7760 28549 7788 28580
rect 8665 28577 8677 28611
rect 8711 28608 8723 28611
rect 8711 28580 9168 28608
rect 8711 28577 8723 28580
rect 8665 28571 8723 28577
rect 7745 28543 7803 28549
rect 7745 28509 7757 28543
rect 7791 28509 7803 28543
rect 7745 28503 7803 28509
rect 7929 28543 7987 28549
rect 7929 28509 7941 28543
rect 7975 28540 7987 28543
rect 8478 28540 8484 28552
rect 7975 28512 8484 28540
rect 7975 28509 7987 28512
rect 7929 28503 7987 28509
rect 8478 28500 8484 28512
rect 8536 28540 8542 28552
rect 8573 28543 8631 28549
rect 8573 28540 8585 28543
rect 8536 28512 8585 28540
rect 8536 28500 8542 28512
rect 8573 28509 8585 28512
rect 8619 28509 8631 28543
rect 8573 28503 8631 28509
rect 8757 28543 8815 28549
rect 8757 28509 8769 28543
rect 8803 28540 8815 28543
rect 8846 28540 8852 28552
rect 8803 28512 8852 28540
rect 8803 28509 8815 28512
rect 8757 28503 8815 28509
rect 6196 28472 6224 28500
rect 5460 28444 6224 28472
rect 7377 28475 7435 28481
rect 7377 28441 7389 28475
rect 7423 28472 7435 28475
rect 8294 28472 8300 28484
rect 7423 28444 8300 28472
rect 7423 28441 7435 28444
rect 7377 28435 7435 28441
rect 8294 28432 8300 28444
rect 8352 28432 8358 28484
rect 2593 28407 2651 28413
rect 2593 28373 2605 28407
rect 2639 28373 2651 28407
rect 2593 28367 2651 28373
rect 2958 28364 2964 28416
rect 3016 28364 3022 28416
rect 3053 28407 3111 28413
rect 3053 28373 3065 28407
rect 3099 28404 3111 28407
rect 3234 28404 3240 28416
rect 3099 28376 3240 28404
rect 3099 28373 3111 28376
rect 3053 28367 3111 28373
rect 3234 28364 3240 28376
rect 3292 28364 3298 28416
rect 3510 28364 3516 28416
rect 3568 28364 3574 28416
rect 3786 28364 3792 28416
rect 3844 28364 3850 28416
rect 6270 28364 6276 28416
rect 6328 28364 6334 28416
rect 6730 28364 6736 28416
rect 6788 28364 6794 28416
rect 7193 28407 7251 28413
rect 7193 28373 7205 28407
rect 7239 28404 7251 28407
rect 7282 28404 7288 28416
rect 7239 28376 7288 28404
rect 7239 28373 7251 28376
rect 7193 28367 7251 28373
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 8588 28404 8616 28503
rect 8846 28500 8852 28512
rect 8904 28500 8910 28552
rect 9140 28549 9168 28580
rect 8941 28543 8999 28549
rect 8941 28509 8953 28543
rect 8987 28509 8999 28543
rect 8941 28503 8999 28509
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 8956 28472 8984 28503
rect 9030 28472 9036 28484
rect 8956 28444 9036 28472
rect 9030 28432 9036 28444
rect 9088 28472 9094 28484
rect 9232 28472 9260 28648
rect 9493 28645 9505 28648
rect 9539 28645 9551 28679
rect 9493 28639 9551 28645
rect 9401 28611 9459 28617
rect 9401 28577 9413 28611
rect 9447 28608 9459 28611
rect 9858 28608 9864 28620
rect 9447 28580 9864 28608
rect 9447 28577 9459 28580
rect 9401 28571 9459 28577
rect 9858 28568 9864 28580
rect 9916 28568 9922 28620
rect 14200 28617 14228 28716
rect 14366 28704 14372 28716
rect 14424 28744 14430 28756
rect 14424 28716 14688 28744
rect 14424 28704 14430 28716
rect 14550 28636 14556 28688
rect 14608 28636 14614 28688
rect 14660 28676 14688 28716
rect 14734 28704 14740 28756
rect 14792 28744 14798 28756
rect 14921 28747 14979 28753
rect 14921 28744 14933 28747
rect 14792 28716 14933 28744
rect 14792 28704 14798 28716
rect 14921 28713 14933 28716
rect 14967 28713 14979 28747
rect 14921 28707 14979 28713
rect 17126 28704 17132 28756
rect 17184 28704 17190 28756
rect 17589 28747 17647 28753
rect 17589 28713 17601 28747
rect 17635 28744 17647 28747
rect 18046 28744 18052 28756
rect 17635 28716 18052 28744
rect 17635 28713 17647 28716
rect 17589 28707 17647 28713
rect 18046 28704 18052 28716
rect 18104 28704 18110 28756
rect 14660 28648 15332 28676
rect 14185 28611 14243 28617
rect 14185 28577 14197 28611
rect 14231 28577 14243 28611
rect 14185 28571 14243 28577
rect 14645 28611 14703 28617
rect 14645 28577 14657 28611
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 9677 28543 9735 28549
rect 9677 28540 9689 28543
rect 9088 28444 9260 28472
rect 9324 28512 9689 28540
rect 9088 28432 9094 28444
rect 9324 28416 9352 28512
rect 9677 28509 9689 28512
rect 9723 28509 9735 28543
rect 9677 28503 9735 28509
rect 9766 28500 9772 28552
rect 9824 28500 9830 28552
rect 10318 28500 10324 28552
rect 10376 28500 10382 28552
rect 10594 28500 10600 28552
rect 10652 28500 10658 28552
rect 13817 28543 13875 28549
rect 13817 28509 13829 28543
rect 13863 28540 13875 28543
rect 14090 28540 14096 28552
rect 13863 28512 14096 28540
rect 13863 28509 13875 28512
rect 13817 28503 13875 28509
rect 14090 28500 14096 28512
rect 14148 28500 14154 28552
rect 14660 28540 14688 28571
rect 15304 28552 15332 28648
rect 17144 28608 17172 28704
rect 17221 28679 17279 28685
rect 17221 28645 17233 28679
rect 17267 28676 17279 28679
rect 17954 28676 17960 28688
rect 17267 28648 17960 28676
rect 17267 28645 17279 28648
rect 17221 28639 17279 28645
rect 17954 28636 17960 28648
rect 18012 28636 18018 28688
rect 17144 28580 17448 28608
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14660 28512 14749 28540
rect 14737 28509 14749 28512
rect 14783 28509 14795 28543
rect 14737 28503 14795 28509
rect 15286 28500 15292 28552
rect 15344 28500 15350 28552
rect 15378 28500 15384 28552
rect 15436 28500 15442 28552
rect 17037 28543 17095 28549
rect 17037 28509 17049 28543
rect 17083 28540 17095 28543
rect 17218 28540 17224 28552
rect 17083 28512 17224 28540
rect 17083 28509 17095 28512
rect 17037 28503 17095 28509
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 17420 28549 17448 28580
rect 17405 28543 17463 28549
rect 17405 28509 17417 28543
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 17865 28543 17923 28549
rect 17865 28509 17877 28543
rect 17911 28540 17923 28543
rect 18138 28540 18144 28552
rect 17911 28512 18144 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18874 28500 18880 28552
rect 18932 28540 18938 28552
rect 19245 28543 19303 28549
rect 19245 28540 19257 28543
rect 18932 28512 19257 28540
rect 18932 28500 18938 28512
rect 19245 28509 19257 28512
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 21450 28500 21456 28552
rect 21508 28500 21514 28552
rect 14292 28444 18184 28472
rect 9306 28404 9312 28416
rect 8588 28376 9312 28404
rect 9306 28364 9312 28376
rect 9364 28364 9370 28416
rect 11698 28364 11704 28416
rect 11756 28404 11762 28416
rect 14292 28404 14320 28444
rect 11756 28376 14320 28404
rect 11756 28364 11762 28376
rect 15194 28364 15200 28416
rect 15252 28364 15258 28416
rect 18046 28364 18052 28416
rect 18104 28364 18110 28416
rect 18156 28404 18184 28444
rect 19150 28432 19156 28484
rect 19208 28472 19214 28484
rect 19490 28475 19548 28481
rect 19490 28472 19502 28475
rect 19208 28444 19502 28472
rect 19208 28432 19214 28444
rect 19490 28441 19502 28444
rect 19536 28441 19548 28475
rect 25866 28472 25872 28484
rect 19490 28435 19548 28441
rect 19628 28444 25872 28472
rect 19628 28404 19656 28444
rect 25866 28432 25872 28444
rect 25924 28432 25930 28484
rect 18156 28376 19656 28404
rect 20622 28364 20628 28416
rect 20680 28364 20686 28416
rect 21634 28364 21640 28416
rect 21692 28364 21698 28416
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 1762 28209 1768 28212
rect 1755 28203 1768 28209
rect 1755 28200 1767 28203
rect 1723 28172 1767 28200
rect 1755 28169 1767 28172
rect 1755 28163 1768 28169
rect 1762 28160 1768 28163
rect 1820 28160 1826 28212
rect 2130 28160 2136 28212
rect 2188 28200 2194 28212
rect 2188 28172 2774 28200
rect 2188 28160 2194 28172
rect 2225 28135 2283 28141
rect 2225 28101 2237 28135
rect 2271 28132 2283 28135
rect 2590 28132 2596 28144
rect 2271 28104 2596 28132
rect 2271 28101 2283 28104
rect 2225 28095 2283 28101
rect 2590 28092 2596 28104
rect 2648 28092 2654 28144
rect 2038 28024 2044 28076
rect 2096 28064 2102 28076
rect 2498 28064 2504 28076
rect 2096 28036 2504 28064
rect 2096 28024 2102 28036
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2746 28064 2774 28172
rect 3510 28160 3516 28212
rect 3568 28160 3574 28212
rect 5626 28160 5632 28212
rect 5684 28200 5690 28212
rect 5721 28203 5779 28209
rect 5721 28200 5733 28203
rect 5684 28172 5733 28200
rect 5684 28160 5690 28172
rect 5721 28169 5733 28172
rect 5767 28169 5779 28203
rect 6270 28200 6276 28212
rect 5721 28163 5779 28169
rect 5920 28172 6276 28200
rect 3528 28132 3556 28160
rect 5920 28141 5948 28172
rect 6270 28160 6276 28172
rect 6328 28160 6334 28212
rect 6730 28160 6736 28212
rect 6788 28200 6794 28212
rect 7377 28203 7435 28209
rect 7377 28200 7389 28203
rect 6788 28172 7389 28200
rect 6788 28160 6794 28172
rect 7377 28169 7389 28172
rect 7423 28169 7435 28203
rect 7377 28163 7435 28169
rect 7742 28160 7748 28212
rect 7800 28160 7806 28212
rect 9030 28160 9036 28212
rect 9088 28200 9094 28212
rect 9088 28172 9168 28200
rect 9088 28160 9094 28172
rect 3252 28104 3556 28132
rect 5905 28135 5963 28141
rect 3252 28073 3280 28104
rect 5905 28101 5917 28135
rect 5951 28101 5963 28135
rect 5905 28095 5963 28101
rect 6914 28092 6920 28144
rect 6972 28132 6978 28144
rect 6972 28104 7328 28132
rect 6972 28092 6978 28104
rect 3510 28073 3516 28076
rect 2869 28067 2927 28073
rect 2869 28064 2881 28067
rect 2746 28036 2881 28064
rect 2869 28033 2881 28036
rect 2915 28033 2927 28067
rect 2869 28027 2927 28033
rect 3237 28067 3295 28073
rect 3237 28033 3249 28067
rect 3283 28033 3295 28067
rect 3237 28027 3295 28033
rect 3478 28067 3516 28073
rect 3478 28033 3490 28067
rect 3478 28027 3516 28033
rect 3510 28024 3516 28027
rect 3568 28024 3574 28076
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28064 4215 28067
rect 4246 28064 4252 28076
rect 4203 28036 4252 28064
rect 4203 28033 4215 28036
rect 4157 28027 4215 28033
rect 4246 28024 4252 28036
rect 4304 28024 4310 28076
rect 4424 28067 4482 28073
rect 4424 28033 4436 28067
rect 4470 28064 4482 28067
rect 4798 28064 4804 28076
rect 4470 28036 4804 28064
rect 4470 28033 4482 28036
rect 4424 28027 4482 28033
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 5629 28067 5687 28073
rect 5629 28064 5641 28067
rect 5276 28036 5641 28064
rect 2317 27999 2375 28005
rect 2317 27965 2329 27999
rect 2363 27996 2375 27999
rect 3142 27996 3148 28008
rect 2363 27968 3148 27996
rect 2363 27965 2375 27968
rect 2317 27959 2375 27965
rect 3142 27956 3148 27968
rect 3200 27956 3206 28008
rect 5276 27940 5304 28036
rect 5629 28033 5641 28036
rect 5675 28033 5687 28067
rect 5629 28027 5687 28033
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 6822 28024 6828 28076
rect 6880 28024 6886 28076
rect 7300 28073 7328 28104
rect 7009 28067 7067 28073
rect 7009 28064 7021 28067
rect 6932 28036 7021 28064
rect 5258 27888 5264 27940
rect 5316 27888 5322 27940
rect 6932 27928 6960 28036
rect 7009 28033 7021 28036
rect 7055 28033 7067 28067
rect 7009 28027 7067 28033
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28033 7343 28067
rect 7285 28027 7343 28033
rect 7469 28067 7527 28073
rect 7469 28033 7481 28067
rect 7515 28064 7527 28067
rect 7760 28064 7788 28160
rect 8386 28092 8392 28144
rect 8444 28132 8450 28144
rect 9140 28141 9168 28172
rect 9306 28160 9312 28212
rect 9364 28160 9370 28212
rect 10045 28203 10103 28209
rect 10045 28169 10057 28203
rect 10091 28200 10103 28203
rect 10594 28200 10600 28212
rect 10091 28172 10600 28200
rect 10091 28169 10103 28172
rect 10045 28163 10103 28169
rect 10594 28160 10600 28172
rect 10652 28160 10658 28212
rect 15194 28160 15200 28212
rect 15252 28160 15258 28212
rect 18046 28160 18052 28212
rect 18104 28160 18110 28212
rect 19150 28160 19156 28212
rect 19208 28160 19214 28212
rect 19702 28160 19708 28212
rect 19760 28160 19766 28212
rect 21634 28160 21640 28212
rect 21692 28200 21698 28212
rect 21692 28172 22094 28200
rect 21692 28160 21698 28172
rect 9125 28135 9183 28141
rect 8444 28104 9076 28132
rect 8444 28092 8450 28104
rect 7515 28036 7788 28064
rect 8941 28067 8999 28073
rect 7515 28033 7527 28036
rect 7469 28027 7527 28033
rect 8941 28033 8953 28067
rect 8987 28033 8999 28067
rect 9048 28064 9076 28104
rect 9125 28101 9137 28135
rect 9171 28101 9183 28135
rect 9324 28132 9352 28160
rect 9585 28135 9643 28141
rect 9324 28104 9428 28132
rect 9125 28095 9183 28101
rect 9355 28101 9428 28104
rect 9355 28067 9367 28101
rect 9401 28070 9428 28101
rect 9585 28101 9597 28135
rect 9631 28132 9643 28135
rect 9766 28132 9772 28144
rect 9631 28104 9772 28132
rect 9631 28101 9643 28104
rect 9585 28095 9643 28101
rect 9401 28067 9413 28070
rect 9048 28036 9260 28064
rect 9355 28061 9413 28067
rect 8941 28027 8999 28033
rect 8956 27996 8984 28027
rect 9232 27996 9260 28036
rect 9600 27996 9628 28095
rect 9766 28092 9772 28104
rect 9824 28092 9830 28144
rect 14912 28135 14970 28141
rect 14912 28101 14924 28135
rect 14958 28132 14970 28135
rect 15212 28132 15240 28160
rect 14958 28104 15240 28132
rect 18064 28132 18092 28160
rect 18610 28135 18668 28141
rect 18610 28132 18622 28135
rect 18064 28104 18622 28132
rect 14958 28101 14970 28104
rect 14912 28095 14970 28101
rect 18610 28101 18622 28104
rect 18656 28101 18668 28135
rect 18610 28095 18668 28101
rect 20524 28135 20582 28141
rect 20524 28101 20536 28135
rect 20570 28132 20582 28135
rect 20714 28132 20720 28144
rect 20570 28104 20720 28132
rect 20570 28101 20582 28104
rect 20524 28095 20582 28101
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 22066 28141 22094 28172
rect 22066 28135 22124 28141
rect 22066 28101 22078 28135
rect 22112 28101 22124 28135
rect 22066 28095 22124 28101
rect 9858 28024 9864 28076
rect 9916 28024 9922 28076
rect 9950 28024 9956 28076
rect 10008 28024 10014 28076
rect 12802 28024 12808 28076
rect 12860 28024 12866 28076
rect 14093 28067 14151 28073
rect 14093 28033 14105 28067
rect 14139 28033 14151 28067
rect 14093 28027 14151 28033
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28064 14335 28067
rect 15654 28064 15660 28076
rect 14323 28036 15660 28064
rect 14323 28033 14335 28036
rect 14277 28027 14335 28033
rect 8956 27968 9168 27996
rect 9232 27968 9628 27996
rect 8757 27931 8815 27937
rect 8757 27928 8769 27931
rect 6564 27900 6960 27928
rect 7024 27900 8769 27928
rect 6564 27872 6592 27900
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 3050 27860 3056 27872
rect 2832 27832 3056 27860
rect 2832 27820 2838 27832
rect 3050 27820 3056 27832
rect 3108 27860 3114 27872
rect 3237 27863 3295 27869
rect 3237 27860 3249 27863
rect 3108 27832 3249 27860
rect 3108 27820 3114 27832
rect 3237 27829 3249 27832
rect 3283 27829 3295 27863
rect 3237 27823 3295 27829
rect 3326 27820 3332 27872
rect 3384 27869 3390 27872
rect 3384 27863 3433 27869
rect 3384 27829 3387 27863
rect 3421 27829 3433 27863
rect 3384 27823 3433 27829
rect 3384 27820 3390 27823
rect 5074 27820 5080 27872
rect 5132 27860 5138 27872
rect 5534 27860 5540 27872
rect 5132 27832 5540 27860
rect 5132 27820 5138 27832
rect 5534 27820 5540 27832
rect 5592 27820 5598 27872
rect 5902 27820 5908 27872
rect 5960 27820 5966 27872
rect 6546 27820 6552 27872
rect 6604 27820 6610 27872
rect 6730 27820 6736 27872
rect 6788 27860 6794 27872
rect 7024 27860 7052 27900
rect 8757 27897 8769 27900
rect 8803 27897 8815 27931
rect 8757 27891 8815 27897
rect 9140 27928 9168 27968
rect 9140 27900 9444 27928
rect 6788 27832 7052 27860
rect 6788 27820 6794 27832
rect 7190 27820 7196 27872
rect 7248 27820 7254 27872
rect 8478 27820 8484 27872
rect 8536 27860 8542 27872
rect 9140 27860 9168 27900
rect 8536 27832 9168 27860
rect 9217 27863 9275 27869
rect 8536 27820 8542 27832
rect 9217 27829 9229 27863
rect 9263 27860 9275 27863
rect 9306 27860 9312 27872
rect 9263 27832 9312 27860
rect 9263 27829 9275 27832
rect 9217 27823 9275 27829
rect 9306 27820 9312 27832
rect 9364 27820 9370 27872
rect 9416 27869 9444 27900
rect 9401 27863 9459 27869
rect 9401 27829 9413 27863
rect 9447 27829 9459 27863
rect 9401 27823 9459 27829
rect 12618 27820 12624 27872
rect 12676 27820 12682 27872
rect 13906 27820 13912 27872
rect 13964 27820 13970 27872
rect 14108 27860 14136 28027
rect 15654 28024 15660 28036
rect 15712 28024 15718 28076
rect 18966 28024 18972 28076
rect 19024 28024 19030 28076
rect 19886 28024 19892 28076
rect 19944 28024 19950 28076
rect 14642 27956 14648 28008
rect 14700 27956 14706 28008
rect 18874 27956 18880 28008
rect 18932 27996 18938 28008
rect 20257 27999 20315 28005
rect 20257 27996 20269 27999
rect 18932 27968 20269 27996
rect 18932 27956 18938 27968
rect 20257 27965 20269 27968
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 21634 27956 21640 28008
rect 21692 27996 21698 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21692 27968 21833 27996
rect 21692 27956 21698 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 15562 27860 15568 27872
rect 14108 27832 15568 27860
rect 15562 27820 15568 27832
rect 15620 27860 15626 27872
rect 16025 27863 16083 27869
rect 16025 27860 16037 27863
rect 15620 27832 16037 27860
rect 15620 27820 15626 27832
rect 16025 27829 16037 27832
rect 16071 27829 16083 27863
rect 16025 27823 16083 27829
rect 17494 27820 17500 27872
rect 17552 27820 17558 27872
rect 21174 27820 21180 27872
rect 21232 27860 21238 27872
rect 21637 27863 21695 27869
rect 21637 27860 21649 27863
rect 21232 27832 21649 27860
rect 21232 27820 21238 27832
rect 21637 27829 21649 27832
rect 21683 27829 21695 27863
rect 21637 27823 21695 27829
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 22244 27832 23213 27860
rect 22244 27820 22250 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 4246 27616 4252 27668
rect 4304 27656 4310 27668
rect 4304 27628 5396 27656
rect 4304 27616 4310 27628
rect 2866 27548 2872 27600
rect 2924 27548 2930 27600
rect 4798 27548 4804 27600
rect 4856 27588 4862 27600
rect 4893 27591 4951 27597
rect 4893 27588 4905 27591
rect 4856 27560 4905 27588
rect 4856 27548 4862 27560
rect 4893 27557 4905 27560
rect 4939 27557 4951 27591
rect 5368 27588 5396 27628
rect 7558 27616 7564 27668
rect 7616 27656 7622 27668
rect 9858 27656 9864 27668
rect 7616 27628 9864 27656
rect 7616 27616 7622 27628
rect 9858 27616 9864 27628
rect 9916 27656 9922 27668
rect 10410 27656 10416 27668
rect 9916 27628 10416 27656
rect 9916 27616 9922 27628
rect 10410 27616 10416 27628
rect 10468 27616 10474 27668
rect 14502 27628 15240 27656
rect 5368 27560 5580 27588
rect 4893 27551 4951 27557
rect 1670 27480 1676 27532
rect 1728 27520 1734 27532
rect 1765 27523 1823 27529
rect 1765 27520 1777 27523
rect 1728 27492 1777 27520
rect 1728 27480 1734 27492
rect 1765 27489 1777 27492
rect 1811 27520 1823 27523
rect 2317 27523 2375 27529
rect 2317 27520 2329 27523
rect 1811 27492 2329 27520
rect 1811 27489 1823 27492
rect 1765 27483 1823 27489
rect 2317 27489 2329 27492
rect 2363 27489 2375 27523
rect 2317 27483 2375 27489
rect 3326 27480 3332 27532
rect 3384 27480 3390 27532
rect 4433 27523 4491 27529
rect 4433 27489 4445 27523
rect 4479 27489 4491 27523
rect 4433 27483 4491 27489
rect 4617 27523 4675 27529
rect 4617 27489 4629 27523
rect 4663 27520 4675 27523
rect 4982 27520 4988 27532
rect 4663 27492 4988 27520
rect 4663 27489 4675 27492
rect 4617 27483 4675 27489
rect 2133 27455 2191 27461
rect 2133 27452 2145 27455
rect 2056 27424 2145 27452
rect 2056 27328 2084 27424
rect 2133 27421 2145 27424
rect 2179 27421 2191 27455
rect 2133 27415 2191 27421
rect 2222 27412 2228 27464
rect 2280 27412 2286 27464
rect 2409 27455 2467 27461
rect 2409 27421 2421 27455
rect 2455 27452 2467 27455
rect 2498 27452 2504 27464
rect 2455 27424 2504 27452
rect 2455 27421 2467 27424
rect 2409 27415 2467 27421
rect 2498 27412 2504 27424
rect 2556 27412 2562 27464
rect 3142 27412 3148 27464
rect 3200 27452 3206 27464
rect 3421 27455 3479 27461
rect 3421 27452 3433 27455
rect 3200 27424 3433 27452
rect 3200 27412 3206 27424
rect 3421 27421 3433 27424
rect 3467 27421 3479 27455
rect 4448 27452 4476 27483
rect 4982 27480 4988 27492
rect 5040 27520 5046 27532
rect 5350 27520 5356 27532
rect 5040 27492 5356 27520
rect 5040 27480 5046 27492
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 4798 27452 4804 27464
rect 4448 27424 4804 27452
rect 3421 27415 3479 27421
rect 3436 27384 3464 27415
rect 4798 27412 4804 27424
rect 4856 27412 4862 27464
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27421 4951 27455
rect 4893 27415 4951 27421
rect 5077 27455 5135 27461
rect 5077 27421 5089 27455
rect 5123 27452 5135 27455
rect 5166 27452 5172 27464
rect 5123 27424 5172 27452
rect 5123 27421 5135 27424
rect 5077 27415 5135 27421
rect 4908 27384 4936 27415
rect 5166 27412 5172 27424
rect 5224 27452 5230 27464
rect 5442 27452 5448 27464
rect 5224 27424 5448 27452
rect 5224 27412 5230 27424
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 5552 27452 5580 27560
rect 8938 27548 8944 27600
rect 8996 27588 9002 27600
rect 9125 27591 9183 27597
rect 9125 27588 9137 27591
rect 8996 27560 9137 27588
rect 8996 27548 9002 27560
rect 9125 27557 9137 27560
rect 9171 27557 9183 27591
rect 9125 27551 9183 27557
rect 10318 27520 10324 27532
rect 9232 27492 10324 27520
rect 6825 27455 6883 27461
rect 6825 27452 6837 27455
rect 5552 27424 6837 27452
rect 6825 27421 6837 27424
rect 6871 27452 6883 27455
rect 6914 27452 6920 27464
rect 6871 27424 6920 27452
rect 6871 27421 6883 27424
rect 6825 27415 6883 27421
rect 6914 27412 6920 27424
rect 6972 27452 6978 27464
rect 9232 27452 9260 27492
rect 10318 27480 10324 27492
rect 10376 27520 10382 27532
rect 10413 27523 10471 27529
rect 10413 27520 10425 27523
rect 10376 27492 10425 27520
rect 10376 27480 10382 27492
rect 10413 27489 10425 27492
rect 10459 27489 10471 27523
rect 14502 27520 14530 27628
rect 15212 27600 15240 27628
rect 15304 27628 17080 27656
rect 15304 27600 15332 27628
rect 14645 27591 14703 27597
rect 14645 27557 14657 27591
rect 14691 27557 14703 27591
rect 14645 27551 14703 27557
rect 10413 27483 10471 27489
rect 14476 27492 14530 27520
rect 14660 27520 14688 27551
rect 15194 27548 15200 27600
rect 15252 27548 15258 27600
rect 15286 27548 15292 27600
rect 15344 27548 15350 27600
rect 17052 27588 17080 27628
rect 18138 27616 18144 27668
rect 18196 27616 18202 27668
rect 18877 27659 18935 27665
rect 18877 27625 18889 27659
rect 18923 27656 18935 27659
rect 18966 27656 18972 27668
rect 18923 27628 18972 27656
rect 18923 27625 18935 27628
rect 18877 27619 18935 27625
rect 18966 27616 18972 27628
rect 19024 27616 19030 27668
rect 19886 27616 19892 27668
rect 19944 27656 19950 27668
rect 19981 27659 20039 27665
rect 19981 27656 19993 27659
rect 19944 27628 19993 27656
rect 19944 27616 19950 27628
rect 19981 27625 19993 27628
rect 20027 27625 20039 27659
rect 19981 27619 20039 27625
rect 20714 27616 20720 27668
rect 20772 27616 20778 27668
rect 21450 27616 21456 27668
rect 21508 27616 21514 27668
rect 22186 27616 22192 27668
rect 22244 27616 22250 27668
rect 17052 27560 17172 27588
rect 17144 27520 17172 27560
rect 17402 27548 17408 27600
rect 17460 27588 17466 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17460 27560 17509 27588
rect 17460 27548 17466 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27588 18107 27591
rect 20622 27588 20628 27600
rect 18095 27560 20628 27588
rect 18095 27557 18107 27560
rect 18049 27551 18107 27557
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 22005 27591 22063 27597
rect 22005 27557 22017 27591
rect 22051 27588 22063 27591
rect 22204 27588 22232 27616
rect 22051 27560 22232 27588
rect 22051 27557 22063 27560
rect 22005 27551 22063 27557
rect 21542 27520 21548 27532
rect 14660 27492 15424 27520
rect 6972 27424 9260 27452
rect 6972 27412 6978 27424
rect 9306 27412 9312 27464
rect 9364 27412 9370 27464
rect 10686 27412 10692 27464
rect 10744 27412 10750 27464
rect 12345 27455 12403 27461
rect 12345 27421 12357 27455
rect 12391 27452 12403 27455
rect 12434 27452 12440 27464
rect 12391 27424 12440 27452
rect 12391 27421 12403 27424
rect 12345 27415 12403 27421
rect 12434 27412 12440 27424
rect 12492 27412 12498 27464
rect 12618 27461 12624 27464
rect 12612 27452 12624 27461
rect 12579 27424 12624 27452
rect 12612 27415 12624 27424
rect 12618 27412 12624 27415
rect 12676 27412 12682 27464
rect 14476 27461 14504 27492
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13740 27424 14105 27452
rect 5902 27384 5908 27396
rect 3436 27356 4844 27384
rect 4908 27356 5908 27384
rect 2038 27276 2044 27328
rect 2096 27276 2102 27328
rect 2130 27276 2136 27328
rect 2188 27276 2194 27328
rect 3329 27319 3387 27325
rect 3329 27285 3341 27319
rect 3375 27316 3387 27319
rect 3789 27319 3847 27325
rect 3789 27316 3801 27319
rect 3375 27288 3801 27316
rect 3375 27285 3387 27288
rect 3329 27279 3387 27285
rect 3789 27285 3801 27288
rect 3835 27285 3847 27319
rect 3789 27279 3847 27285
rect 4154 27276 4160 27328
rect 4212 27276 4218 27328
rect 4246 27276 4252 27328
rect 4304 27276 4310 27328
rect 4816 27316 4844 27356
rect 5902 27344 5908 27356
rect 5960 27344 5966 27396
rect 6580 27387 6638 27393
rect 6580 27353 6592 27387
rect 6626 27384 6638 27387
rect 6730 27384 6736 27396
rect 6626 27356 6736 27384
rect 6626 27353 6638 27356
rect 6580 27347 6638 27353
rect 6730 27344 6736 27356
rect 6788 27344 6794 27396
rect 7190 27393 7196 27396
rect 7184 27384 7196 27393
rect 7151 27356 7196 27384
rect 7184 27347 7196 27356
rect 7190 27344 7196 27347
rect 7248 27344 7254 27396
rect 12069 27387 12127 27393
rect 12069 27353 12081 27387
rect 12115 27384 12127 27387
rect 13630 27384 13636 27396
rect 12115 27356 13636 27384
rect 12115 27353 12127 27356
rect 12069 27347 12127 27353
rect 13630 27344 13636 27356
rect 13688 27344 13694 27396
rect 4890 27316 4896 27328
rect 4816 27288 4896 27316
rect 4890 27276 4896 27288
rect 4948 27276 4954 27328
rect 5445 27319 5503 27325
rect 5445 27285 5457 27319
rect 5491 27316 5503 27319
rect 5534 27316 5540 27328
rect 5491 27288 5540 27316
rect 5491 27285 5503 27288
rect 5445 27279 5503 27285
rect 5534 27276 5540 27288
rect 5592 27276 5598 27328
rect 8297 27319 8355 27325
rect 8297 27285 8309 27319
rect 8343 27316 8355 27319
rect 8478 27316 8484 27328
rect 8343 27288 8484 27316
rect 8343 27285 8355 27288
rect 8297 27279 8355 27285
rect 8478 27276 8484 27288
rect 8536 27276 8542 27328
rect 9122 27276 9128 27328
rect 9180 27316 9186 27328
rect 11698 27316 11704 27328
rect 9180 27288 11704 27316
rect 9180 27276 9186 27288
rect 11698 27276 11704 27288
rect 11756 27276 11762 27328
rect 13170 27276 13176 27328
rect 13228 27316 13234 27328
rect 13740 27325 13768 27424
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 14734 27412 14740 27464
rect 14792 27412 14798 27464
rect 14918 27412 14924 27464
rect 14976 27412 14982 27464
rect 15010 27412 15016 27464
rect 15068 27412 15074 27464
rect 15105 27455 15163 27461
rect 15105 27421 15117 27455
rect 15151 27452 15163 27455
rect 15194 27452 15200 27464
rect 15151 27424 15200 27452
rect 15151 27421 15163 27424
rect 15105 27415 15163 27421
rect 15194 27412 15200 27424
rect 15252 27412 15258 27464
rect 15286 27412 15292 27464
rect 15344 27412 15350 27464
rect 15396 27461 15424 27492
rect 15672 27492 16252 27520
rect 17144 27492 21548 27520
rect 15562 27461 15568 27464
rect 15381 27455 15439 27461
rect 15381 27421 15393 27455
rect 15427 27421 15439 27455
rect 15381 27415 15439 27421
rect 15529 27455 15568 27461
rect 15529 27421 15541 27455
rect 15529 27415 15568 27421
rect 15562 27412 15568 27415
rect 15620 27412 15626 27464
rect 15672 27461 15700 27492
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 15746 27412 15752 27464
rect 15804 27412 15810 27464
rect 15887 27455 15945 27461
rect 15887 27421 15899 27455
rect 15933 27452 15945 27455
rect 15933 27424 16068 27452
rect 15933 27421 15945 27424
rect 15887 27415 15945 27421
rect 14277 27387 14335 27393
rect 14277 27353 14289 27387
rect 14323 27353 14335 27387
rect 14277 27347 14335 27353
rect 14369 27387 14427 27393
rect 14369 27353 14381 27387
rect 14415 27384 14427 27387
rect 14568 27384 14596 27412
rect 14415 27356 14596 27384
rect 14415 27353 14427 27356
rect 14369 27347 14427 27353
rect 13725 27319 13783 27325
rect 13725 27316 13737 27319
rect 13228 27288 13737 27316
rect 13228 27276 13234 27288
rect 13725 27285 13737 27288
rect 13771 27285 13783 27319
rect 14292 27316 14320 27347
rect 14936 27316 14964 27412
rect 15304 27384 15332 27412
rect 16040 27384 16068 27424
rect 16114 27412 16120 27464
rect 16172 27412 16178 27464
rect 16224 27452 16252 27492
rect 21542 27480 21548 27492
rect 21600 27520 21606 27532
rect 21729 27523 21787 27529
rect 21729 27520 21741 27523
rect 21600 27492 21741 27520
rect 21600 27480 21606 27492
rect 21729 27489 21741 27492
rect 21775 27489 21787 27523
rect 21729 27483 21787 27489
rect 22189 27523 22247 27529
rect 22189 27489 22201 27523
rect 22235 27489 22247 27523
rect 22189 27483 22247 27489
rect 23584 27492 23980 27520
rect 16224 27424 16896 27452
rect 16868 27396 16896 27424
rect 19610 27412 19616 27464
rect 19668 27452 19674 27464
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 19668 27424 20269 27452
rect 19668 27412 19674 27424
rect 20257 27421 20269 27424
rect 20303 27452 20315 27455
rect 20625 27455 20683 27461
rect 20303 27424 20576 27452
rect 20303 27421 20315 27424
rect 20257 27415 20315 27421
rect 20548 27396 20576 27424
rect 20625 27421 20637 27455
rect 20671 27452 20683 27455
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 20671 27424 20913 27452
rect 20671 27421 20683 27424
rect 20625 27415 20683 27421
rect 20901 27421 20913 27424
rect 20947 27421 20959 27455
rect 22204 27452 22232 27483
rect 23584 27452 23612 27492
rect 23952 27461 23980 27492
rect 22204 27424 23612 27452
rect 23661 27455 23719 27461
rect 20901 27415 20959 27421
rect 23661 27421 23673 27455
rect 23707 27452 23719 27455
rect 23937 27455 23995 27461
rect 23707 27424 23888 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 16384 27387 16442 27393
rect 15304 27356 15608 27384
rect 16040 27356 16160 27384
rect 15580 27328 15608 27356
rect 16132 27328 16160 27356
rect 16384 27353 16396 27387
rect 16430 27384 16442 27387
rect 16574 27384 16580 27396
rect 16430 27356 16580 27384
rect 16430 27353 16442 27356
rect 16384 27347 16442 27353
rect 16574 27344 16580 27356
rect 16632 27344 16638 27396
rect 16850 27344 16856 27396
rect 16908 27344 16914 27396
rect 17678 27344 17684 27396
rect 17736 27344 17742 27396
rect 18509 27387 18567 27393
rect 18509 27353 18521 27387
rect 18555 27353 18567 27387
rect 18509 27347 18567 27353
rect 18693 27387 18751 27393
rect 18693 27353 18705 27387
rect 18739 27384 18751 27387
rect 19426 27384 19432 27396
rect 18739 27356 19432 27384
rect 18739 27353 18751 27356
rect 18693 27347 18751 27353
rect 14292 27288 14964 27316
rect 13725 27279 13783 27285
rect 15286 27276 15292 27328
rect 15344 27276 15350 27328
rect 15562 27276 15568 27328
rect 15620 27276 15626 27328
rect 16022 27276 16028 27328
rect 16080 27276 16086 27328
rect 16114 27276 16120 27328
rect 16172 27276 16178 27328
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 18524 27316 18552 27347
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 19794 27344 19800 27396
rect 19852 27344 19858 27396
rect 20438 27344 20444 27396
rect 20496 27344 20502 27396
rect 20530 27344 20536 27396
rect 20588 27384 20594 27396
rect 21085 27387 21143 27393
rect 21085 27384 21097 27387
rect 20588 27356 21097 27384
rect 20588 27344 20594 27356
rect 21085 27353 21097 27356
rect 21131 27353 21143 27387
rect 21085 27347 21143 27353
rect 21174 27344 21180 27396
rect 21232 27384 21238 27396
rect 21269 27387 21327 27393
rect 21269 27384 21281 27387
rect 21232 27356 21281 27384
rect 21232 27344 21238 27356
rect 21269 27353 21281 27356
rect 21315 27353 21327 27387
rect 21269 27347 21327 27353
rect 23416 27387 23474 27393
rect 23416 27353 23428 27387
rect 23462 27384 23474 27387
rect 23860 27384 23888 27424
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 24394 27412 24400 27464
rect 24452 27412 24458 27464
rect 24412 27384 24440 27412
rect 23462 27356 23796 27384
rect 23860 27356 24440 27384
rect 23462 27353 23474 27356
rect 23416 27347 23474 27353
rect 20806 27316 20812 27328
rect 16540 27288 20812 27316
rect 16540 27276 16546 27288
rect 20806 27276 20812 27288
rect 20864 27276 20870 27328
rect 22281 27319 22339 27325
rect 22281 27285 22293 27319
rect 22327 27316 22339 27319
rect 22922 27316 22928 27328
rect 22327 27288 22928 27316
rect 22327 27285 22339 27288
rect 22281 27279 22339 27285
rect 22922 27276 22928 27288
rect 22980 27276 22986 27328
rect 23768 27325 23796 27356
rect 23753 27319 23811 27325
rect 23753 27285 23765 27319
rect 23799 27285 23811 27319
rect 23753 27279 23811 27285
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1670 27112 1676 27124
rect 1412 27084 1676 27112
rect 1412 26985 1440 27084
rect 1670 27072 1676 27084
rect 1728 27072 1734 27124
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 1857 27115 1915 27121
rect 1857 27112 1869 27115
rect 1811 27084 1869 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 1857 27081 1869 27084
rect 1903 27112 1915 27115
rect 2130 27112 2136 27124
rect 1903 27084 2136 27112
rect 1903 27081 1915 27084
rect 1857 27075 1915 27081
rect 1872 26985 1900 27075
rect 2130 27072 2136 27084
rect 2188 27112 2194 27124
rect 2685 27115 2743 27121
rect 2685 27112 2697 27115
rect 2188 27084 2697 27112
rect 2188 27072 2194 27084
rect 2685 27081 2697 27084
rect 2731 27081 2743 27115
rect 2685 27075 2743 27081
rect 5166 27072 5172 27124
rect 5224 27072 5230 27124
rect 6822 27112 6828 27124
rect 5276 27084 6828 27112
rect 2498 27004 2504 27056
rect 2556 27044 2562 27056
rect 2556 27016 4108 27044
rect 2556 27004 2562 27016
rect 1397 26979 1455 26985
rect 1397 26945 1409 26979
rect 1443 26945 1455 26979
rect 1857 26979 1915 26985
rect 1857 26976 1869 26979
rect 1397 26939 1455 26945
rect 1688 26948 1869 26976
rect 1688 26840 1716 26948
rect 1857 26945 1869 26948
rect 1903 26945 1915 26979
rect 1857 26939 1915 26945
rect 2038 26936 2044 26988
rect 2096 26976 2102 26988
rect 2961 26979 3019 26985
rect 2961 26976 2973 26979
rect 2096 26948 2452 26976
rect 2096 26936 2102 26948
rect 1765 26911 1823 26917
rect 1765 26877 1777 26911
rect 1811 26908 1823 26911
rect 2148 26908 2176 26948
rect 1811 26880 2176 26908
rect 1811 26877 1823 26880
rect 1765 26871 1823 26877
rect 2222 26868 2228 26920
rect 2280 26908 2286 26920
rect 2317 26911 2375 26917
rect 2317 26908 2329 26911
rect 2280 26880 2329 26908
rect 2280 26868 2286 26880
rect 2317 26877 2329 26880
rect 2363 26877 2375 26911
rect 2424 26908 2452 26948
rect 2700 26948 2973 26976
rect 2700 26908 2728 26948
rect 2961 26945 2973 26948
rect 3007 26945 3019 26979
rect 2961 26939 3019 26945
rect 3050 26936 3056 26988
rect 3108 26936 3114 26988
rect 3326 26936 3332 26988
rect 3384 26936 3390 26988
rect 3510 26936 3516 26988
rect 3568 26936 3574 26988
rect 4080 26985 4108 27016
rect 4154 27004 4160 27056
rect 4212 27044 4218 27056
rect 5276 27044 5304 27084
rect 6822 27072 6828 27084
rect 6880 27072 6886 27124
rect 7098 27072 7104 27124
rect 7156 27112 7162 27124
rect 9769 27115 9827 27121
rect 9769 27112 9781 27115
rect 7156 27084 9781 27112
rect 7156 27072 7162 27084
rect 9769 27081 9781 27084
rect 9815 27081 9827 27115
rect 9769 27075 9827 27081
rect 10686 27072 10692 27124
rect 10744 27072 10750 27124
rect 13449 27115 13507 27121
rect 13449 27081 13461 27115
rect 13495 27081 13507 27115
rect 13449 27075 13507 27081
rect 4212 27016 5304 27044
rect 5337 27047 5395 27053
rect 4212 27004 4218 27016
rect 5337 27013 5349 27047
rect 5383 27013 5395 27047
rect 5337 27007 5395 27013
rect 4065 26979 4123 26985
rect 4065 26976 4077 26979
rect 4023 26948 4077 26976
rect 4065 26945 4077 26948
rect 4111 26945 4123 26979
rect 4065 26939 4123 26945
rect 2424 26880 2728 26908
rect 2317 26871 2375 26877
rect 2685 26843 2743 26849
rect 2685 26840 2697 26843
rect 1688 26812 2697 26840
rect 2685 26809 2697 26812
rect 2731 26840 2743 26843
rect 2866 26840 2872 26852
rect 2731 26812 2872 26840
rect 2731 26809 2743 26812
rect 2685 26803 2743 26809
rect 2866 26800 2872 26812
rect 2924 26800 2930 26852
rect 2958 26800 2964 26852
rect 3016 26840 3022 26852
rect 3237 26843 3295 26849
rect 3237 26840 3249 26843
rect 3016 26812 3249 26840
rect 3016 26800 3022 26812
rect 3237 26809 3249 26812
rect 3283 26840 3295 26843
rect 3602 26840 3608 26852
rect 3283 26812 3608 26840
rect 3283 26809 3295 26812
rect 3237 26803 3295 26809
rect 3602 26800 3608 26812
rect 3660 26800 3666 26852
rect 4080 26840 4108 26939
rect 5258 26868 5264 26920
rect 5316 26908 5322 26920
rect 5352 26908 5380 27007
rect 5534 27004 5540 27056
rect 5592 27044 5598 27056
rect 5592 27016 6040 27044
rect 5592 27004 5598 27016
rect 6012 26985 6040 27016
rect 6086 27004 6092 27056
rect 6144 27044 6150 27056
rect 8938 27044 8944 27056
rect 6144 27016 8944 27044
rect 6144 27004 6150 27016
rect 8938 27004 8944 27016
rect 8996 27004 9002 27056
rect 12434 27044 12440 27056
rect 11716 27016 12440 27044
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26976 6055 26979
rect 6043 26948 6500 26976
rect 6043 26945 6055 26948
rect 5997 26939 6055 26945
rect 5828 26908 5856 26939
rect 6270 26908 6276 26920
rect 5316 26880 6276 26908
rect 5316 26868 5322 26880
rect 6270 26868 6276 26880
rect 6328 26868 6334 26920
rect 6472 26917 6500 26948
rect 7374 26936 7380 26988
rect 7432 26976 7438 26988
rect 7745 26979 7803 26985
rect 7745 26976 7757 26979
rect 7432 26948 7757 26976
rect 7432 26936 7438 26948
rect 7745 26945 7757 26948
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26976 8079 26979
rect 8478 26976 8484 26988
rect 8067 26948 8484 26976
rect 8067 26945 8079 26948
rect 8021 26939 8079 26945
rect 8478 26936 8484 26948
rect 8536 26936 8542 26988
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 6457 26911 6515 26917
rect 6457 26877 6469 26911
rect 6503 26908 6515 26911
rect 7929 26911 7987 26917
rect 6503 26880 7696 26908
rect 6503 26877 6515 26880
rect 6457 26871 6515 26877
rect 5994 26840 6000 26852
rect 4080 26812 6000 26840
rect 5994 26800 6000 26812
rect 6052 26800 6058 26852
rect 6086 26800 6092 26852
rect 6144 26840 6150 26852
rect 7561 26843 7619 26849
rect 7561 26840 7573 26843
rect 6144 26812 7573 26840
rect 6144 26800 6150 26812
rect 7561 26809 7573 26812
rect 7607 26809 7619 26843
rect 7668 26840 7696 26880
rect 7929 26877 7941 26911
rect 7975 26908 7987 26911
rect 8294 26908 8300 26920
rect 7975 26880 8300 26908
rect 7975 26877 7987 26880
rect 7929 26871 7987 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 9324 26908 9352 26939
rect 10410 26936 10416 26988
rect 10468 26936 10474 26988
rect 11716 26985 11744 27016
rect 12434 27004 12440 27016
rect 12492 27004 12498 27056
rect 13464 27044 13492 27075
rect 13906 27072 13912 27124
rect 13964 27072 13970 27124
rect 14734 27072 14740 27124
rect 14792 27072 14798 27124
rect 15286 27072 15292 27124
rect 15344 27072 15350 27124
rect 15378 27072 15384 27124
rect 15436 27072 15442 27124
rect 17494 27112 17500 27124
rect 16832 27084 17500 27112
rect 13786 27047 13844 27053
rect 13786 27044 13798 27047
rect 13464 27016 13798 27044
rect 13786 27013 13798 27016
rect 13832 27013 13844 27047
rect 13786 27007 13844 27013
rect 11974 26985 11980 26988
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 11968 26939 11980 26985
rect 9180 26880 9352 26908
rect 9180 26868 9186 26880
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 9677 26911 9735 26917
rect 9677 26908 9689 26911
rect 9456 26880 9689 26908
rect 9456 26868 9462 26880
rect 9677 26877 9689 26880
rect 9723 26877 9735 26911
rect 9677 26871 9735 26877
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26877 9919 26911
rect 10612 26908 10640 26939
rect 11974 26936 11980 26939
rect 12032 26936 12038 26988
rect 13265 26979 13323 26985
rect 13265 26945 13277 26979
rect 13311 26976 13323 26979
rect 13924 26976 13952 27072
rect 13311 26948 13952 26976
rect 13311 26945 13323 26948
rect 13265 26939 13323 26945
rect 9861 26871 9919 26877
rect 10244 26880 10640 26908
rect 7668 26812 9536 26840
rect 7561 26803 7619 26809
rect 2884 26772 2912 26800
rect 9508 26784 9536 26812
rect 3694 26772 3700 26784
rect 2884 26744 3700 26772
rect 3694 26732 3700 26744
rect 3752 26732 3758 26784
rect 5074 26732 5080 26784
rect 5132 26772 5138 26784
rect 5353 26775 5411 26781
rect 5353 26772 5365 26775
rect 5132 26744 5365 26772
rect 5132 26732 5138 26744
rect 5353 26741 5365 26744
rect 5399 26741 5411 26775
rect 5353 26735 5411 26741
rect 6181 26775 6239 26781
rect 6181 26741 6193 26775
rect 6227 26772 6239 26775
rect 6362 26772 6368 26784
rect 6227 26744 6368 26772
rect 6227 26741 6239 26744
rect 6181 26735 6239 26741
rect 6362 26732 6368 26744
rect 6420 26732 6426 26784
rect 7006 26732 7012 26784
rect 7064 26732 7070 26784
rect 7650 26732 7656 26784
rect 7708 26772 7714 26784
rect 7745 26775 7803 26781
rect 7745 26772 7757 26775
rect 7708 26744 7757 26772
rect 7708 26732 7714 26744
rect 7745 26741 7757 26744
rect 7791 26741 7803 26775
rect 7745 26735 7803 26741
rect 9214 26732 9220 26784
rect 9272 26772 9278 26784
rect 9401 26775 9459 26781
rect 9401 26772 9413 26775
rect 9272 26744 9413 26772
rect 9272 26732 9278 26744
rect 9401 26741 9413 26744
rect 9447 26741 9459 26775
rect 9401 26735 9459 26741
rect 9490 26732 9496 26784
rect 9548 26732 9554 26784
rect 9876 26772 9904 26871
rect 10244 26849 10272 26880
rect 12894 26868 12900 26920
rect 12952 26908 12958 26920
rect 13541 26911 13599 26917
rect 13541 26908 13553 26911
rect 12952 26880 13553 26908
rect 12952 26868 12958 26880
rect 13541 26877 13553 26880
rect 13587 26877 13599 26911
rect 13541 26871 13599 26877
rect 10229 26843 10287 26849
rect 10229 26809 10241 26843
rect 10275 26809 10287 26843
rect 10229 26803 10287 26809
rect 11054 26772 11060 26784
rect 9876 26744 11060 26772
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 14752 26772 14780 27072
rect 15304 27044 15332 27072
rect 15304 27016 16712 27044
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26945 15623 26979
rect 15565 26939 15623 26945
rect 15580 26908 15608 26939
rect 15654 26936 15660 26988
rect 15712 26976 15718 26988
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15712 26948 15761 26976
rect 15712 26936 15718 26948
rect 15749 26945 15761 26948
rect 15795 26976 15807 26979
rect 16482 26976 16488 26988
rect 15795 26948 16488 26976
rect 15795 26945 15807 26948
rect 15749 26939 15807 26945
rect 16482 26936 16488 26948
rect 16540 26936 16546 26988
rect 16684 26985 16712 27016
rect 16832 26985 16860 27084
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 21600 27084 22600 27112
rect 21600 27072 21606 27084
rect 17037 27047 17095 27053
rect 17037 27013 17049 27047
rect 17083 27044 17095 27047
rect 17402 27044 17408 27056
rect 17083 27016 17408 27044
rect 17083 27013 17095 27016
rect 17037 27007 17095 27013
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 19337 27047 19395 27053
rect 19337 27013 19349 27047
rect 19383 27044 19395 27047
rect 19610 27044 19616 27056
rect 19383 27016 19616 27044
rect 19383 27013 19395 27016
rect 19337 27007 19395 27013
rect 19610 27004 19616 27016
rect 19668 27004 19674 27056
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16817 26979 16875 26985
rect 16817 26945 16829 26979
rect 16863 26945 16875 26979
rect 16817 26939 16875 26945
rect 16832 26908 16860 26939
rect 16942 26936 16948 26988
rect 17000 26936 17006 26988
rect 17134 26979 17192 26985
rect 17134 26976 17146 26979
rect 17052 26948 17146 26976
rect 15580 26880 16860 26908
rect 17052 26840 17080 26948
rect 17134 26945 17146 26948
rect 17180 26945 17192 26979
rect 17134 26939 17192 26945
rect 19150 26936 19156 26988
rect 19208 26936 19214 26988
rect 19702 26985 19708 26988
rect 19696 26939 19708 26985
rect 19702 26936 19708 26939
rect 19760 26936 19766 26988
rect 18046 26868 18052 26920
rect 18104 26908 18110 26920
rect 18874 26908 18880 26920
rect 18104 26880 18880 26908
rect 18104 26868 18110 26880
rect 18874 26868 18880 26880
rect 18932 26908 18938 26920
rect 22572 26917 22600 27084
rect 23934 26936 23940 26988
rect 23992 26976 23998 26988
rect 24222 26979 24280 26985
rect 24222 26976 24234 26979
rect 23992 26948 24234 26976
rect 23992 26936 23998 26948
rect 24222 26945 24234 26948
rect 24268 26945 24280 26979
rect 24222 26939 24280 26945
rect 24394 26936 24400 26988
rect 24452 26976 24458 26988
rect 24489 26979 24547 26985
rect 24489 26976 24501 26979
rect 24452 26948 24501 26976
rect 24452 26936 24458 26948
rect 24489 26945 24501 26948
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 19429 26911 19487 26917
rect 19429 26908 19441 26911
rect 18932 26880 19441 26908
rect 18932 26868 18938 26880
rect 19429 26877 19441 26880
rect 19475 26877 19487 26911
rect 19429 26871 19487 26877
rect 22557 26911 22615 26917
rect 22557 26877 22569 26911
rect 22603 26908 22615 26911
rect 23290 26908 23296 26920
rect 22603 26880 23296 26908
rect 22603 26877 22615 26880
rect 22557 26871 22615 26877
rect 23290 26868 23296 26880
rect 23348 26868 23354 26920
rect 16132 26812 17080 26840
rect 16132 26784 16160 26812
rect 22922 26800 22928 26852
rect 22980 26800 22986 26852
rect 13136 26744 14780 26772
rect 13136 26732 13142 26744
rect 14826 26732 14832 26784
rect 14884 26772 14890 26784
rect 14921 26775 14979 26781
rect 14921 26772 14933 26775
rect 14884 26744 14933 26772
rect 14884 26732 14890 26744
rect 14921 26741 14933 26744
rect 14967 26741 14979 26775
rect 14921 26735 14979 26741
rect 16114 26732 16120 26784
rect 16172 26732 16178 26784
rect 17034 26732 17040 26784
rect 17092 26772 17098 26784
rect 17313 26775 17371 26781
rect 17313 26772 17325 26775
rect 17092 26744 17325 26772
rect 17092 26732 17098 26744
rect 17313 26741 17325 26744
rect 17359 26741 17371 26775
rect 17313 26735 17371 26741
rect 18966 26732 18972 26784
rect 19024 26732 19030 26784
rect 20070 26732 20076 26784
rect 20128 26772 20134 26784
rect 20438 26772 20444 26784
rect 20128 26744 20444 26772
rect 20128 26732 20134 26744
rect 20438 26732 20444 26744
rect 20496 26772 20502 26784
rect 20809 26775 20867 26781
rect 20809 26772 20821 26775
rect 20496 26744 20821 26772
rect 20496 26732 20502 26744
rect 20809 26741 20821 26744
rect 20855 26741 20867 26775
rect 20809 26735 20867 26741
rect 23014 26732 23020 26784
rect 23072 26732 23078 26784
rect 23106 26732 23112 26784
rect 23164 26732 23170 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 2866 26528 2872 26580
rect 2924 26568 2930 26580
rect 3326 26568 3332 26580
rect 2924 26540 3332 26568
rect 2924 26528 2930 26540
rect 3326 26528 3332 26540
rect 3384 26568 3390 26580
rect 4709 26571 4767 26577
rect 4709 26568 4721 26571
rect 3384 26540 4721 26568
rect 3384 26528 3390 26540
rect 4709 26537 4721 26540
rect 4755 26537 4767 26571
rect 4709 26531 4767 26537
rect 4893 26571 4951 26577
rect 4893 26537 4905 26571
rect 4939 26568 4951 26571
rect 4982 26568 4988 26580
rect 4939 26540 4988 26568
rect 4939 26537 4951 26540
rect 4893 26531 4951 26537
rect 4982 26528 4988 26540
rect 5040 26568 5046 26580
rect 5534 26568 5540 26580
rect 5040 26540 5540 26568
rect 5040 26528 5046 26540
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 5994 26528 6000 26580
rect 6052 26528 6058 26580
rect 6086 26528 6092 26580
rect 6144 26528 6150 26580
rect 6730 26528 6736 26580
rect 6788 26568 6794 26580
rect 6825 26571 6883 26577
rect 6825 26568 6837 26571
rect 6788 26540 6837 26568
rect 6788 26528 6794 26540
rect 6825 26537 6837 26540
rect 6871 26537 6883 26571
rect 6825 26531 6883 26537
rect 7006 26528 7012 26580
rect 7064 26528 7070 26580
rect 9950 26528 9956 26580
rect 10008 26528 10014 26580
rect 11974 26528 11980 26580
rect 12032 26528 12038 26580
rect 12713 26571 12771 26577
rect 12713 26537 12725 26571
rect 12759 26568 12771 26571
rect 12802 26568 12808 26580
rect 12759 26540 12808 26568
rect 12759 26537 12771 26540
rect 12713 26531 12771 26537
rect 12802 26528 12808 26540
rect 12860 26528 12866 26580
rect 13078 26528 13084 26580
rect 13136 26528 13142 26580
rect 16574 26528 16580 26580
rect 16632 26528 16638 26580
rect 17310 26528 17316 26580
rect 17368 26568 17374 26580
rect 17368 26540 18460 26568
rect 17368 26528 17374 26540
rect 4065 26503 4123 26509
rect 4065 26500 4077 26503
rect 2746 26472 4077 26500
rect 2746 26444 2774 26472
rect 4065 26469 4077 26472
rect 4111 26500 4123 26503
rect 4338 26500 4344 26512
rect 4111 26472 4344 26500
rect 4111 26469 4123 26472
rect 4065 26463 4123 26469
rect 4338 26460 4344 26472
rect 4396 26460 4402 26512
rect 6012 26500 6040 26528
rect 4908 26472 6040 26500
rect 2682 26392 2688 26444
rect 2740 26404 2774 26444
rect 4356 26404 4844 26432
rect 2740 26392 2746 26404
rect 2958 26324 2964 26376
rect 3016 26364 3022 26376
rect 3510 26364 3516 26376
rect 3016 26336 3516 26364
rect 3016 26324 3022 26336
rect 3510 26324 3516 26336
rect 3568 26364 3574 26376
rect 4356 26373 4384 26404
rect 4816 26376 4844 26404
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3568 26336 3985 26364
rect 3568 26324 3574 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26333 4399 26367
rect 4341 26327 4399 26333
rect 4522 26324 4528 26376
rect 4580 26324 4586 26376
rect 4798 26324 4804 26376
rect 4856 26324 4862 26376
rect 3418 26256 3424 26308
rect 3476 26256 3482 26308
rect 4908 26305 4936 26472
rect 5074 26392 5080 26444
rect 5132 26392 5138 26444
rect 5997 26435 6055 26441
rect 5997 26401 6009 26435
rect 6043 26432 6055 26435
rect 6104 26432 6132 26528
rect 6043 26404 6132 26432
rect 6043 26401 6055 26404
rect 5997 26395 6055 26401
rect 6270 26392 6276 26444
rect 6328 26432 6334 26444
rect 6328 26404 6960 26432
rect 6328 26392 6334 26404
rect 5092 26364 5120 26392
rect 5537 26367 5595 26373
rect 5537 26364 5549 26367
rect 5092 26336 5549 26364
rect 5537 26333 5549 26336
rect 5583 26333 5595 26367
rect 5537 26327 5595 26333
rect 5902 26324 5908 26376
rect 5960 26324 5966 26376
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 6362 26324 6368 26376
rect 6420 26324 6426 26376
rect 6546 26324 6552 26376
rect 6604 26364 6610 26376
rect 6932 26373 6960 26404
rect 6641 26367 6699 26373
rect 6641 26364 6653 26367
rect 6604 26336 6653 26364
rect 6604 26324 6610 26336
rect 6641 26333 6653 26336
rect 6687 26333 6699 26367
rect 6641 26327 6699 26333
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26333 6975 26367
rect 7024 26364 7052 26528
rect 12621 26503 12679 26509
rect 12621 26469 12633 26503
rect 12667 26500 12679 26503
rect 13096 26500 13124 26528
rect 12667 26472 13124 26500
rect 12667 26469 12679 26472
rect 12621 26463 12679 26469
rect 13170 26460 13176 26512
rect 13228 26460 13234 26512
rect 13630 26460 13636 26512
rect 13688 26500 13694 26512
rect 16758 26500 16764 26512
rect 13688 26472 16764 26500
rect 13688 26460 13694 26472
rect 16758 26460 16764 26472
rect 16816 26460 16822 26512
rect 17405 26503 17463 26509
rect 17405 26469 17417 26503
rect 17451 26469 17463 26503
rect 18432 26500 18460 26540
rect 19702 26528 19708 26580
rect 19760 26528 19766 26580
rect 23014 26528 23020 26580
rect 23072 26528 23078 26580
rect 23569 26571 23627 26577
rect 23569 26537 23581 26571
rect 23615 26568 23627 26571
rect 23934 26568 23940 26580
rect 23615 26540 23940 26568
rect 23615 26537 23627 26540
rect 23569 26531 23627 26537
rect 23934 26528 23940 26540
rect 23992 26528 23998 26580
rect 20717 26503 20775 26509
rect 20717 26500 20729 26503
rect 18432 26472 20729 26500
rect 17405 26463 17463 26469
rect 20717 26469 20729 26472
rect 20763 26469 20775 26503
rect 20717 26463 20775 26469
rect 9493 26435 9551 26441
rect 9493 26432 9505 26435
rect 9232 26404 9505 26432
rect 7101 26367 7159 26373
rect 7101 26364 7113 26367
rect 7024 26336 7113 26364
rect 6917 26327 6975 26333
rect 7101 26333 7113 26336
rect 7147 26333 7159 26367
rect 7101 26327 7159 26333
rect 9232 26308 9260 26404
rect 9493 26401 9505 26404
rect 9539 26401 9551 26435
rect 9493 26395 9551 26401
rect 11054 26392 11060 26444
rect 11112 26432 11118 26444
rect 14458 26432 14464 26444
rect 11112 26404 14464 26432
rect 11112 26392 11118 26404
rect 14458 26392 14464 26404
rect 14516 26392 14522 26444
rect 17420 26432 17448 26463
rect 17420 26404 17632 26432
rect 12158 26324 12164 26376
rect 12216 26324 12222 26376
rect 15746 26324 15752 26376
rect 15804 26324 15810 26376
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26364 16819 26367
rect 17126 26364 17132 26376
rect 16807 26336 17132 26364
rect 16807 26333 16819 26336
rect 16761 26327 16819 26333
rect 17126 26324 17132 26336
rect 17184 26324 17190 26376
rect 17218 26324 17224 26376
rect 17276 26324 17282 26376
rect 17497 26367 17555 26373
rect 17497 26333 17509 26367
rect 17543 26333 17555 26367
rect 17604 26364 17632 26404
rect 18966 26392 18972 26444
rect 19024 26392 19030 26444
rect 17753 26367 17811 26373
rect 17753 26364 17765 26367
rect 17604 26336 17765 26364
rect 17497 26327 17555 26333
rect 17753 26333 17765 26336
rect 17799 26333 17811 26367
rect 17753 26327 17811 26333
rect 4893 26299 4951 26305
rect 4893 26265 4905 26299
rect 4939 26265 4951 26299
rect 4893 26259 4951 26265
rect 5077 26299 5135 26305
rect 5077 26265 5089 26299
rect 5123 26265 5135 26299
rect 7009 26299 7067 26305
rect 7009 26296 7021 26299
rect 5077 26259 5135 26265
rect 6472 26268 7021 26296
rect 2130 26188 2136 26240
rect 2188 26188 2194 26240
rect 4338 26188 4344 26240
rect 4396 26228 4402 26240
rect 5092 26228 5120 26259
rect 6472 26237 6500 26268
rect 7009 26265 7021 26268
rect 7055 26265 7067 26299
rect 7009 26259 7067 26265
rect 9214 26256 9220 26308
rect 9272 26256 9278 26308
rect 9398 26256 9404 26308
rect 9456 26256 9462 26308
rect 9490 26256 9496 26308
rect 9548 26256 9554 26308
rect 12253 26299 12311 26305
rect 12253 26265 12265 26299
rect 12299 26296 12311 26299
rect 12805 26299 12863 26305
rect 12805 26296 12817 26299
rect 12299 26268 12817 26296
rect 12299 26265 12311 26268
rect 12253 26259 12311 26265
rect 12805 26265 12817 26268
rect 12851 26296 12863 26299
rect 13078 26296 13084 26308
rect 12851 26268 13084 26296
rect 12851 26265 12863 26268
rect 12805 26259 12863 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 17512 26296 17540 26327
rect 18046 26324 18052 26376
rect 18104 26324 18110 26376
rect 18984 26364 19012 26392
rect 19521 26367 19579 26373
rect 19521 26364 19533 26367
rect 18984 26336 19533 26364
rect 19521 26333 19533 26336
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 21358 26324 21364 26376
rect 21416 26364 21422 26376
rect 22097 26367 22155 26373
rect 22097 26364 22109 26367
rect 21416 26336 22109 26364
rect 21416 26324 21422 26336
rect 22097 26333 22109 26336
rect 22143 26333 22155 26367
rect 23032 26364 23060 26528
rect 23385 26367 23443 26373
rect 23385 26364 23397 26367
rect 23032 26336 23397 26364
rect 22097 26327 22155 26333
rect 23385 26333 23397 26336
rect 23431 26333 23443 26367
rect 23385 26327 23443 26333
rect 18064 26296 18092 26324
rect 19426 26296 19432 26308
rect 17512 26268 18092 26296
rect 18892 26268 19432 26296
rect 4396 26200 5120 26228
rect 6457 26231 6515 26237
rect 4396 26188 4402 26200
rect 6457 26197 6469 26231
rect 6503 26197 6515 26231
rect 6457 26191 6515 26197
rect 6546 26188 6552 26240
rect 6604 26228 6610 26240
rect 9122 26228 9128 26240
rect 6604 26200 9128 26228
rect 6604 26188 6610 26200
rect 9122 26188 9128 26200
rect 9180 26228 9186 26240
rect 10594 26228 10600 26240
rect 9180 26200 10600 26228
rect 9180 26188 9186 26200
rect 10594 26188 10600 26200
rect 10652 26188 10658 26240
rect 13262 26188 13268 26240
rect 13320 26188 13326 26240
rect 15565 26231 15623 26237
rect 15565 26197 15577 26231
rect 15611 26228 15623 26231
rect 15654 26228 15660 26240
rect 15611 26200 15660 26228
rect 15611 26197 15623 26200
rect 15565 26191 15623 26197
rect 15654 26188 15660 26200
rect 15712 26188 15718 26240
rect 18892 26237 18920 26268
rect 19426 26256 19432 26268
rect 19484 26256 19490 26308
rect 21450 26256 21456 26308
rect 21508 26296 21514 26308
rect 21830 26299 21888 26305
rect 21830 26296 21842 26299
rect 21508 26268 21842 26296
rect 21508 26256 21514 26268
rect 21830 26265 21842 26268
rect 21876 26265 21888 26299
rect 21830 26259 21888 26265
rect 18877 26231 18935 26237
rect 18877 26197 18889 26231
rect 18923 26197 18935 26231
rect 18877 26191 18935 26197
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 2130 25984 2136 26036
rect 2188 26024 2194 26036
rect 3973 26027 4031 26033
rect 2188 25996 3556 26024
rect 2188 25984 2194 25996
rect 2639 25959 2697 25965
rect 2639 25925 2651 25959
rect 2685 25956 2697 25959
rect 2866 25956 2872 25968
rect 2685 25928 2872 25956
rect 2685 25925 2697 25928
rect 2639 25919 2697 25925
rect 2866 25916 2872 25928
rect 2924 25916 2930 25968
rect 2961 25959 3019 25965
rect 2961 25925 2973 25959
rect 3007 25956 3019 25959
rect 3050 25956 3056 25968
rect 3007 25928 3056 25956
rect 3007 25925 3019 25928
rect 2961 25919 3019 25925
rect 3050 25916 3056 25928
rect 3108 25916 3114 25968
rect 2133 25891 2191 25897
rect 2133 25857 2145 25891
rect 2179 25888 2191 25891
rect 2222 25888 2228 25900
rect 2179 25860 2228 25888
rect 2179 25857 2191 25860
rect 2133 25851 2191 25857
rect 2222 25848 2228 25860
rect 2280 25848 2286 25900
rect 2314 25848 2320 25900
rect 2372 25848 2378 25900
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 2501 25891 2559 25897
rect 2501 25857 2513 25891
rect 2547 25888 2559 25891
rect 3142 25888 3148 25900
rect 2547 25860 3148 25888
rect 2547 25857 2559 25860
rect 2501 25851 2559 25857
rect 2424 25820 2452 25851
rect 3142 25848 3148 25860
rect 3200 25888 3206 25900
rect 3528 25897 3556 25996
rect 3973 25993 3985 26027
rect 4019 26024 4031 26027
rect 4246 26024 4252 26036
rect 4019 25996 4252 26024
rect 4019 25993 4031 25996
rect 3973 25987 4031 25993
rect 4246 25984 4252 25996
rect 4304 25984 4310 26036
rect 4338 25984 4344 26036
rect 4396 25984 4402 26036
rect 5350 25984 5356 26036
rect 5408 26024 5414 26036
rect 6454 26024 6460 26036
rect 5408 25996 6460 26024
rect 5408 25984 5414 25996
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 7466 25984 7472 26036
rect 7524 26024 7530 26036
rect 7653 26027 7711 26033
rect 7653 26024 7665 26027
rect 7524 25996 7665 26024
rect 7524 25984 7530 25996
rect 7653 25993 7665 25996
rect 7699 25993 7711 26027
rect 10318 26024 10324 26036
rect 7653 25987 7711 25993
rect 9685 25996 10324 26024
rect 4522 25956 4528 25968
rect 3620 25928 4528 25956
rect 3237 25891 3295 25897
rect 3237 25888 3249 25891
rect 3200 25860 3249 25888
rect 3200 25848 3206 25860
rect 3237 25857 3249 25860
rect 3283 25857 3295 25891
rect 3237 25851 3295 25857
rect 3513 25891 3571 25897
rect 3513 25857 3525 25891
rect 3559 25857 3571 25891
rect 3513 25851 3571 25857
rect 2332 25792 2452 25820
rect 2777 25823 2835 25829
rect 2332 25684 2360 25792
rect 2777 25789 2789 25823
rect 2823 25789 2835 25823
rect 2777 25783 2835 25789
rect 2406 25712 2412 25764
rect 2464 25752 2470 25764
rect 2792 25752 2820 25783
rect 2866 25780 2872 25832
rect 2924 25780 2930 25832
rect 3050 25780 3056 25832
rect 3108 25780 3114 25832
rect 3421 25823 3479 25829
rect 3421 25789 3433 25823
rect 3467 25820 3479 25823
rect 3620 25820 3648 25928
rect 4522 25916 4528 25928
rect 4580 25916 4586 25968
rect 4890 25916 4896 25968
rect 4948 25956 4954 25968
rect 4948 25928 5120 25956
rect 4948 25916 4954 25928
rect 3694 25848 3700 25900
rect 3752 25888 3758 25900
rect 3881 25891 3939 25897
rect 3881 25888 3893 25891
rect 3752 25860 3893 25888
rect 3752 25848 3758 25860
rect 3881 25857 3893 25860
rect 3927 25857 3939 25891
rect 3881 25851 3939 25857
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4706 25888 4712 25900
rect 4028 25860 4712 25888
rect 4028 25848 4034 25860
rect 4706 25848 4712 25860
rect 4764 25888 4770 25900
rect 5092 25897 5120 25928
rect 6730 25916 6736 25968
rect 6788 25956 6794 25968
rect 8849 25959 8907 25965
rect 8849 25956 8861 25959
rect 6788 25928 8861 25956
rect 6788 25916 6794 25928
rect 8849 25925 8861 25928
rect 8895 25925 8907 25959
rect 8849 25919 8907 25925
rect 4801 25891 4859 25897
rect 4801 25888 4813 25891
rect 4764 25860 4813 25888
rect 4764 25848 4770 25860
rect 4801 25857 4813 25860
rect 4847 25857 4859 25891
rect 4801 25851 4859 25857
rect 5077 25891 5135 25897
rect 5077 25857 5089 25891
rect 5123 25857 5135 25891
rect 5077 25851 5135 25857
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 3467 25792 3648 25820
rect 4433 25823 4491 25829
rect 3467 25789 3479 25792
rect 3421 25783 3479 25789
rect 4433 25789 4445 25823
rect 4479 25789 4491 25823
rect 4433 25783 4491 25789
rect 4617 25823 4675 25829
rect 4617 25789 4629 25823
rect 4663 25820 4675 25823
rect 4890 25820 4896 25832
rect 4663 25792 4896 25820
rect 4663 25789 4675 25792
rect 4617 25783 4675 25789
rect 3068 25752 3096 25780
rect 2464 25724 3096 25752
rect 2464 25712 2470 25724
rect 3050 25684 3056 25696
rect 2332 25656 3056 25684
rect 3050 25644 3056 25656
rect 3108 25684 3114 25696
rect 3436 25684 3464 25783
rect 4338 25712 4344 25764
rect 4396 25752 4402 25764
rect 4448 25752 4476 25783
rect 4890 25780 4896 25792
rect 4948 25780 4954 25832
rect 7208 25820 7236 25851
rect 7374 25848 7380 25900
rect 7432 25848 7438 25900
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7742 25888 7748 25900
rect 7515 25860 7748 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 7837 25891 7895 25897
rect 7837 25857 7849 25891
rect 7883 25857 7895 25891
rect 7837 25851 7895 25857
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25888 7987 25891
rect 8018 25888 8024 25900
rect 7975 25860 8024 25888
rect 7975 25857 7987 25860
rect 7929 25851 7987 25857
rect 7852 25820 7880 25851
rect 8018 25848 8024 25860
rect 8076 25848 8082 25900
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 7208 25792 7604 25820
rect 4396 25724 4476 25752
rect 4396 25712 4402 25724
rect 4522 25712 4528 25764
rect 4580 25752 4586 25764
rect 6086 25752 6092 25764
rect 4580 25724 6092 25752
rect 4580 25712 4586 25724
rect 6086 25712 6092 25724
rect 6144 25712 6150 25764
rect 7576 25696 7604 25792
rect 7668 25792 7880 25820
rect 7668 25696 7696 25792
rect 8128 25752 8156 25851
rect 8202 25848 8208 25900
rect 8260 25848 8266 25900
rect 8757 25891 8815 25897
rect 8757 25857 8769 25891
rect 8803 25857 8815 25891
rect 8864 25888 8892 25919
rect 9685 25897 9713 25996
rect 10318 25984 10324 25996
rect 10376 26024 10382 26036
rect 11238 26024 11244 26036
rect 10376 25996 11244 26024
rect 10376 25984 10382 25996
rect 11238 25984 11244 25996
rect 11296 25984 11302 26036
rect 13262 25984 13268 26036
rect 13320 25984 13326 26036
rect 15746 25984 15752 26036
rect 15804 25984 15810 26036
rect 15930 25984 15936 26036
rect 15988 26024 15994 26036
rect 15988 25996 16988 26024
rect 15988 25984 15994 25996
rect 10244 25928 10640 25956
rect 10244 25897 10272 25928
rect 9677 25891 9735 25897
rect 9677 25888 9689 25891
rect 8864 25860 9689 25888
rect 8757 25851 8815 25857
rect 9677 25857 9689 25860
rect 9723 25888 9735 25891
rect 10229 25891 10287 25897
rect 9723 25860 9818 25888
rect 9723 25857 9735 25860
rect 9677 25851 9735 25857
rect 10229 25857 10241 25891
rect 10275 25857 10287 25891
rect 10229 25851 10287 25857
rect 10321 25891 10379 25897
rect 10321 25857 10333 25891
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 8478 25780 8484 25832
rect 8536 25820 8542 25832
rect 8772 25820 8800 25851
rect 8536 25792 8800 25820
rect 8536 25780 8542 25792
rect 9766 25780 9772 25832
rect 9824 25820 9830 25832
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9824 25792 9965 25820
rect 9824 25780 9830 25792
rect 9953 25789 9965 25792
rect 9999 25820 10011 25823
rect 10336 25820 10364 25851
rect 10410 25848 10416 25900
rect 10468 25888 10474 25900
rect 10505 25891 10563 25897
rect 10505 25888 10517 25891
rect 10468 25860 10517 25888
rect 10468 25848 10474 25860
rect 10505 25857 10517 25860
rect 10551 25857 10563 25891
rect 10505 25851 10563 25857
rect 10612 25832 10640 25928
rect 12894 25848 12900 25900
rect 12952 25848 12958 25900
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25888 13139 25891
rect 13280 25888 13308 25984
rect 16960 25965 16988 25996
rect 17218 25984 17224 26036
rect 17276 26024 17282 26036
rect 17405 26027 17463 26033
rect 17405 26024 17417 26027
rect 17276 25996 17417 26024
rect 17276 25984 17282 25996
rect 17405 25993 17417 25996
rect 17451 25993 17463 26027
rect 17405 25987 17463 25993
rect 18693 26027 18751 26033
rect 18693 25993 18705 26027
rect 18739 25993 18751 26027
rect 18693 25987 18751 25993
rect 16945 25959 17003 25965
rect 13127 25860 13308 25888
rect 13832 25928 16252 25956
rect 13127 25857 13139 25860
rect 13081 25851 13139 25857
rect 9999 25792 10364 25820
rect 9999 25789 10011 25792
rect 9953 25783 10011 25789
rect 10594 25780 10600 25832
rect 10652 25780 10658 25832
rect 12912 25820 12940 25848
rect 13832 25820 13860 25928
rect 16224 25897 16252 25928
rect 16945 25925 16957 25959
rect 16991 25956 17003 25959
rect 17678 25956 17684 25968
rect 16991 25928 17684 25956
rect 16991 25925 17003 25928
rect 16945 25919 17003 25925
rect 17678 25916 17684 25928
rect 17736 25916 17742 25968
rect 18046 25916 18052 25968
rect 18104 25916 18110 25968
rect 18708 25956 18736 25987
rect 21450 25984 21456 26036
rect 21508 25984 21514 26036
rect 19030 25959 19088 25965
rect 19030 25956 19042 25959
rect 18708 25928 19042 25956
rect 19030 25925 19042 25928
rect 19076 25925 19088 25959
rect 21821 25959 21879 25965
rect 21821 25956 21833 25959
rect 19030 25919 19088 25925
rect 20824 25928 21833 25956
rect 20824 25900 20852 25928
rect 21821 25925 21833 25928
rect 21867 25925 21879 25959
rect 21821 25919 21879 25925
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16209 25891 16267 25897
rect 16209 25857 16221 25891
rect 16255 25857 16267 25891
rect 16209 25851 16267 25857
rect 18233 25891 18291 25897
rect 18233 25857 18245 25891
rect 18279 25857 18291 25891
rect 18233 25851 18291 25857
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 18874 25888 18880 25900
rect 18555 25860 18880 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 12912 25792 13860 25820
rect 15289 25823 15347 25829
rect 15289 25789 15301 25823
rect 15335 25820 15347 25823
rect 15562 25820 15568 25832
rect 15335 25792 15568 25820
rect 15335 25789 15347 25792
rect 15289 25783 15347 25789
rect 15562 25780 15568 25792
rect 15620 25780 15626 25832
rect 16132 25820 16160 25851
rect 16132 25792 16436 25820
rect 15657 25755 15715 25761
rect 8128 25724 11008 25752
rect 10980 25696 11008 25724
rect 15657 25721 15669 25755
rect 15703 25752 15715 25755
rect 15746 25752 15752 25764
rect 15703 25724 15752 25752
rect 15703 25721 15715 25724
rect 15657 25715 15715 25721
rect 15746 25712 15752 25724
rect 15804 25752 15810 25764
rect 16298 25752 16304 25764
rect 15804 25724 16304 25752
rect 15804 25712 15810 25724
rect 16298 25712 16304 25724
rect 16356 25712 16362 25764
rect 3108 25656 3464 25684
rect 3108 25644 3114 25656
rect 3510 25644 3516 25696
rect 3568 25644 3574 25696
rect 3602 25644 3608 25696
rect 3660 25684 3666 25696
rect 4893 25687 4951 25693
rect 4893 25684 4905 25687
rect 3660 25656 4905 25684
rect 3660 25644 3666 25656
rect 4893 25653 4905 25656
rect 4939 25653 4951 25687
rect 4893 25647 4951 25653
rect 5258 25644 5264 25696
rect 5316 25644 5322 25696
rect 6638 25644 6644 25696
rect 6696 25684 6702 25696
rect 7009 25687 7067 25693
rect 7009 25684 7021 25687
rect 6696 25656 7021 25684
rect 6696 25644 6702 25656
rect 7009 25653 7021 25656
rect 7055 25653 7067 25687
rect 7009 25647 7067 25653
rect 7558 25644 7564 25696
rect 7616 25644 7622 25696
rect 7650 25644 7656 25696
rect 7708 25644 7714 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 9493 25687 9551 25693
rect 9493 25684 9505 25687
rect 9088 25656 9505 25684
rect 9088 25644 9094 25656
rect 9493 25653 9505 25656
rect 9539 25653 9551 25687
rect 9493 25647 9551 25653
rect 9861 25687 9919 25693
rect 9861 25653 9873 25687
rect 9907 25684 9919 25687
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 9907 25656 10149 25684
rect 9907 25653 9919 25656
rect 9861 25647 9919 25653
rect 10137 25653 10149 25656
rect 10183 25653 10195 25687
rect 10137 25647 10195 25653
rect 10410 25644 10416 25696
rect 10468 25644 10474 25696
rect 10962 25644 10968 25696
rect 11020 25644 11026 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 12897 25687 12955 25693
rect 12897 25684 12909 25687
rect 12860 25656 12909 25684
rect 12860 25644 12866 25656
rect 12897 25653 12909 25656
rect 12943 25653 12955 25687
rect 12897 25647 12955 25653
rect 15470 25644 15476 25696
rect 15528 25684 15534 25696
rect 15933 25687 15991 25693
rect 15933 25684 15945 25687
rect 15528 25656 15945 25684
rect 15528 25644 15534 25656
rect 15933 25653 15945 25656
rect 15979 25684 15991 25687
rect 16206 25684 16212 25696
rect 15979 25656 16212 25684
rect 15979 25653 15991 25656
rect 15933 25647 15991 25653
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 16408 25693 16436 25792
rect 17310 25712 17316 25764
rect 17368 25712 17374 25764
rect 16393 25687 16451 25693
rect 16393 25653 16405 25687
rect 16439 25684 16451 25687
rect 18248 25684 18276 25851
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 20806 25848 20812 25900
rect 20864 25848 20870 25900
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25888 22063 25891
rect 22554 25888 22560 25900
rect 22051 25860 22560 25888
rect 22051 25857 22063 25860
rect 22005 25851 22063 25857
rect 18782 25780 18788 25832
rect 18840 25780 18846 25832
rect 21284 25820 21312 25851
rect 22554 25848 22560 25860
rect 22612 25888 22618 25900
rect 22612 25860 25820 25888
rect 22612 25848 22618 25860
rect 22189 25823 22247 25829
rect 22189 25820 22201 25823
rect 21284 25792 22201 25820
rect 22189 25789 22201 25792
rect 22235 25789 22247 25823
rect 22189 25783 22247 25789
rect 25792 25764 25820 25860
rect 21634 25752 21640 25764
rect 19720 25724 21640 25752
rect 19720 25684 19748 25724
rect 21634 25712 21640 25724
rect 21692 25712 21698 25764
rect 25774 25712 25780 25764
rect 25832 25712 25838 25764
rect 16439 25656 19748 25684
rect 16439 25653 16451 25656
rect 16393 25647 16451 25653
rect 19794 25644 19800 25696
rect 19852 25684 19858 25696
rect 20165 25687 20223 25693
rect 20165 25684 20177 25687
rect 19852 25656 20177 25684
rect 19852 25644 19858 25656
rect 20165 25653 20177 25656
rect 20211 25653 20223 25687
rect 20165 25647 20223 25653
rect 20254 25644 20260 25696
rect 20312 25684 20318 25696
rect 25866 25684 25872 25696
rect 20312 25656 25872 25684
rect 20312 25644 20318 25656
rect 25866 25644 25872 25656
rect 25924 25644 25930 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 2314 25440 2320 25492
rect 2372 25480 2378 25492
rect 3602 25480 3608 25492
rect 2372 25452 3608 25480
rect 2372 25440 2378 25452
rect 3602 25440 3608 25452
rect 3660 25440 3666 25492
rect 4338 25440 4344 25492
rect 4396 25480 4402 25492
rect 4617 25483 4675 25489
rect 4617 25480 4629 25483
rect 4396 25452 4629 25480
rect 4396 25440 4402 25452
rect 4617 25449 4629 25452
rect 4663 25449 4675 25483
rect 4617 25443 4675 25449
rect 5258 25440 5264 25492
rect 5316 25440 5322 25492
rect 5350 25440 5356 25492
rect 5408 25480 5414 25492
rect 5408 25452 6776 25480
rect 5408 25440 5414 25452
rect 5276 25412 5304 25440
rect 3988 25384 5304 25412
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 2774 25344 2780 25356
rect 2547 25316 2780 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 3053 25279 3111 25285
rect 3053 25245 3065 25279
rect 3099 25245 3111 25279
rect 3053 25239 3111 25245
rect 3068 25208 3096 25239
rect 3326 25236 3332 25288
rect 3384 25236 3390 25288
rect 3988 25285 4016 25384
rect 6638 25372 6644 25424
rect 6696 25372 6702 25424
rect 4798 25304 4804 25356
rect 4856 25344 4862 25356
rect 5169 25347 5227 25353
rect 5169 25344 5181 25347
rect 4856 25316 5181 25344
rect 4856 25304 4862 25316
rect 5169 25313 5181 25316
rect 5215 25313 5227 25347
rect 5718 25344 5724 25356
rect 5169 25307 5227 25313
rect 5368 25316 5724 25344
rect 3513 25279 3571 25285
rect 3513 25245 3525 25279
rect 3559 25276 3571 25279
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3559 25248 3801 25276
rect 3559 25245 3571 25248
rect 3513 25239 3571 25245
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25245 4031 25279
rect 3973 25239 4031 25245
rect 4154 25236 4160 25288
rect 4212 25236 4218 25288
rect 4246 25236 4252 25288
rect 4304 25236 4310 25288
rect 4982 25236 4988 25288
rect 5040 25236 5046 25288
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25276 5135 25279
rect 5368 25276 5396 25316
rect 5718 25304 5724 25316
rect 5776 25304 5782 25356
rect 6656 25344 6684 25372
rect 6380 25316 6684 25344
rect 5123 25248 5396 25276
rect 5445 25279 5503 25285
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 5445 25245 5457 25279
rect 5491 25276 5503 25279
rect 5534 25276 5540 25288
rect 5491 25248 5540 25276
rect 5491 25245 5503 25248
rect 5445 25239 5503 25245
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 6380 25285 6408 25316
rect 6748 25285 6776 25452
rect 8202 25440 8208 25492
rect 8260 25440 8266 25492
rect 10410 25440 10416 25492
rect 10468 25440 10474 25492
rect 10962 25440 10968 25492
rect 11020 25440 11026 25492
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 16816 25452 18828 25480
rect 16816 25440 16822 25452
rect 7282 25372 7288 25424
rect 7340 25412 7346 25424
rect 7742 25412 7748 25424
rect 7340 25384 7748 25412
rect 7340 25372 7346 25384
rect 7742 25372 7748 25384
rect 7800 25372 7806 25424
rect 7837 25415 7895 25421
rect 7837 25381 7849 25415
rect 7883 25412 7895 25415
rect 8220 25412 8248 25440
rect 7883 25384 8248 25412
rect 7883 25381 7895 25384
rect 7837 25375 7895 25381
rect 7193 25347 7251 25353
rect 7193 25313 7205 25347
rect 7239 25344 7251 25347
rect 7852 25344 7880 25375
rect 8386 25372 8392 25424
rect 8444 25412 8450 25424
rect 10137 25415 10195 25421
rect 10137 25412 10149 25415
rect 8444 25384 10149 25412
rect 8444 25372 8450 25384
rect 10137 25381 10149 25384
rect 10183 25381 10195 25415
rect 10137 25375 10195 25381
rect 8941 25347 8999 25353
rect 8941 25344 8953 25347
rect 7239 25316 7880 25344
rect 8128 25316 8953 25344
rect 7239 25313 7251 25316
rect 7193 25307 7251 25313
rect 6365 25279 6423 25285
rect 6365 25245 6377 25279
rect 6411 25245 6423 25279
rect 6365 25239 6423 25245
rect 6457 25279 6515 25285
rect 6457 25245 6469 25279
rect 6503 25245 6515 25279
rect 6457 25239 6515 25245
rect 6641 25279 6699 25285
rect 6641 25245 6653 25279
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25245 6791 25279
rect 6733 25239 6791 25245
rect 7285 25279 7343 25285
rect 7285 25245 7297 25279
rect 7331 25276 7343 25279
rect 7374 25276 7380 25288
rect 7331 25248 7380 25276
rect 7331 25245 7343 25248
rect 7285 25239 7343 25245
rect 6181 25211 6239 25217
rect 6181 25208 6193 25211
rect 3068 25180 6193 25208
rect 6181 25177 6193 25180
rect 6227 25177 6239 25211
rect 6181 25171 6239 25177
rect 3694 25100 3700 25152
rect 3752 25140 3758 25152
rect 5350 25140 5356 25152
rect 3752 25112 5356 25140
rect 3752 25100 3758 25112
rect 5350 25100 5356 25112
rect 5408 25100 5414 25152
rect 5537 25143 5595 25149
rect 5537 25109 5549 25143
rect 5583 25140 5595 25143
rect 5810 25140 5816 25152
rect 5583 25112 5816 25140
rect 5583 25109 5595 25112
rect 5537 25103 5595 25109
rect 5810 25100 5816 25112
rect 5868 25100 5874 25152
rect 6472 25140 6500 25239
rect 6656 25208 6684 25239
rect 7374 25236 7380 25248
rect 7432 25236 7438 25288
rect 7466 25236 7472 25288
rect 7524 25236 7530 25288
rect 7558 25236 7564 25288
rect 7616 25276 7622 25288
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 7616 25248 7665 25276
rect 7616 25236 7622 25248
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 6822 25208 6828 25220
rect 6656 25180 6828 25208
rect 6822 25168 6828 25180
rect 6880 25168 6886 25220
rect 7484 25208 7512 25236
rect 6932 25180 7512 25208
rect 7668 25208 7696 25239
rect 7742 25236 7748 25288
rect 7800 25236 7806 25288
rect 8128 25285 8156 25316
rect 8941 25313 8953 25316
rect 8987 25344 8999 25347
rect 9030 25344 9036 25356
rect 8987 25316 9036 25344
rect 8987 25313 8999 25316
rect 8941 25307 8999 25313
rect 9030 25304 9036 25316
rect 9088 25304 9094 25356
rect 10428 25344 10456 25440
rect 10594 25372 10600 25424
rect 10652 25412 10658 25424
rect 11241 25415 11299 25421
rect 10652 25384 11100 25412
rect 10652 25372 10658 25384
rect 11072 25353 11100 25384
rect 11241 25381 11253 25415
rect 11287 25412 11299 25415
rect 12069 25415 12127 25421
rect 12069 25412 12081 25415
rect 11287 25384 12081 25412
rect 11287 25381 11299 25384
rect 11241 25375 11299 25381
rect 11057 25347 11115 25353
rect 9140 25316 9812 25344
rect 10428 25316 10824 25344
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 8297 25279 8355 25285
rect 8297 25245 8309 25279
rect 8343 25276 8355 25279
rect 8478 25276 8484 25288
rect 8343 25248 8484 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 8757 25279 8815 25285
rect 8628 25248 8708 25276
rect 8628 25236 8634 25248
rect 8386 25208 8392 25220
rect 7668 25180 8392 25208
rect 6932 25140 6960 25180
rect 8386 25168 8392 25180
rect 8444 25168 8450 25220
rect 8680 25208 8708 25248
rect 8757 25245 8769 25279
rect 8803 25276 8815 25279
rect 9140 25276 9168 25316
rect 8803 25248 9168 25276
rect 8803 25245 8815 25248
rect 8757 25239 8815 25245
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 9582 25236 9588 25288
rect 9640 25236 9646 25288
rect 9784 25285 9812 25316
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25276 9827 25279
rect 9858 25276 9864 25288
rect 9815 25248 9864 25276
rect 9815 25245 9827 25248
rect 9769 25239 9827 25245
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 10318 25236 10324 25288
rect 10376 25236 10382 25288
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25245 10471 25279
rect 10413 25239 10471 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 9600 25208 9628 25236
rect 8680 25180 9628 25208
rect 6472 25112 6960 25140
rect 7006 25100 7012 25152
rect 7064 25100 7070 25152
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 7377 25143 7435 25149
rect 7377 25140 7389 25143
rect 7340 25112 7389 25140
rect 7340 25100 7346 25112
rect 7377 25109 7389 25112
rect 7423 25109 7435 25143
rect 7377 25103 7435 25109
rect 7558 25100 7564 25152
rect 7616 25100 7622 25152
rect 7742 25100 7748 25152
rect 7800 25140 7806 25152
rect 8018 25140 8024 25152
rect 7800 25112 8024 25140
rect 7800 25100 7806 25112
rect 8018 25100 8024 25112
rect 8076 25140 8082 25152
rect 8941 25143 8999 25149
rect 8941 25140 8953 25143
rect 8076 25112 8953 25140
rect 8076 25100 8082 25112
rect 8941 25109 8953 25112
rect 8987 25109 8999 25143
rect 10428 25140 10456 25239
rect 10520 25208 10548 25239
rect 10594 25236 10600 25288
rect 10652 25236 10658 25288
rect 10796 25285 10824 25316
rect 11057 25313 11069 25347
rect 11103 25313 11115 25347
rect 11057 25307 11115 25313
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 11517 25347 11575 25353
rect 11517 25344 11529 25347
rect 11195 25316 11529 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 11517 25313 11529 25316
rect 11563 25313 11575 25347
rect 11517 25307 11575 25313
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25276 10839 25279
rect 10873 25279 10931 25285
rect 10873 25276 10885 25279
rect 10827 25248 10885 25276
rect 10827 25245 10839 25248
rect 10781 25239 10839 25245
rect 10873 25245 10885 25248
rect 10919 25245 10931 25279
rect 10873 25239 10931 25245
rect 11238 25236 11244 25288
rect 11296 25276 11302 25288
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11296 25248 11437 25276
rect 11296 25236 11302 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11532 25208 11560 25307
rect 10520 25180 11560 25208
rect 11624 25140 11652 25384
rect 12069 25381 12081 25384
rect 12115 25381 12127 25415
rect 12069 25375 12127 25381
rect 14461 25415 14519 25421
rect 14461 25381 14473 25415
rect 14507 25412 14519 25415
rect 14734 25412 14740 25424
rect 14507 25384 14740 25412
rect 14507 25381 14519 25384
rect 14461 25375 14519 25381
rect 14734 25372 14740 25384
rect 14792 25372 14798 25424
rect 18800 25412 18828 25452
rect 18874 25440 18880 25492
rect 18932 25480 18938 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 18932 25452 19257 25480
rect 18932 25440 18938 25452
rect 19245 25449 19257 25452
rect 19291 25449 19303 25483
rect 19245 25443 19303 25449
rect 21634 25440 21640 25492
rect 21692 25480 21698 25492
rect 21692 25452 24440 25480
rect 21692 25440 21698 25452
rect 20254 25412 20260 25424
rect 18800 25384 20260 25412
rect 20254 25372 20260 25384
rect 20312 25372 20318 25424
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12023 25316 12296 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25276 11759 25279
rect 11790 25276 11796 25288
rect 11747 25248 11796 25276
rect 11747 25245 11759 25248
rect 11701 25239 11759 25245
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 11882 25236 11888 25288
rect 11940 25236 11946 25288
rect 12268 25285 12296 25316
rect 12434 25304 12440 25356
rect 12492 25344 12498 25356
rect 12529 25347 12587 25353
rect 12529 25344 12541 25347
rect 12492 25316 12541 25344
rect 12492 25304 12498 25316
rect 12529 25313 12541 25316
rect 12575 25313 12587 25347
rect 12529 25307 12587 25313
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25313 14611 25347
rect 14553 25307 14611 25313
rect 16868 25316 17448 25344
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 12253 25279 12311 25285
rect 12253 25245 12265 25279
rect 12299 25276 12311 25279
rect 12342 25276 12348 25288
rect 12299 25248 12348 25276
rect 12299 25245 12311 25248
rect 12253 25239 12311 25245
rect 11808 25208 11836 25236
rect 12084 25208 12112 25239
rect 12342 25236 12348 25248
rect 12400 25236 12406 25288
rect 12802 25285 12808 25288
rect 12796 25276 12808 25285
rect 12763 25248 12808 25276
rect 12796 25239 12808 25248
rect 12802 25236 12808 25239
rect 12860 25236 12866 25288
rect 14568 25276 14596 25307
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 14568 25248 14841 25276
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 15381 25279 15439 25285
rect 15381 25245 15393 25279
rect 15427 25276 15439 25279
rect 15470 25276 15476 25288
rect 15427 25248 15476 25276
rect 15427 25245 15439 25248
rect 15381 25239 15439 25245
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 15654 25285 15660 25288
rect 15648 25276 15660 25285
rect 15615 25248 15660 25276
rect 15648 25239 15660 25248
rect 15654 25236 15660 25239
rect 15712 25236 15718 25288
rect 16868 25285 16896 25316
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25245 16911 25279
rect 17313 25279 17371 25285
rect 17313 25276 17325 25279
rect 16853 25239 16911 25245
rect 16960 25248 17325 25276
rect 14093 25211 14151 25217
rect 14093 25208 14105 25211
rect 11808 25180 12112 25208
rect 13832 25180 14105 25208
rect 10428 25112 11652 25140
rect 8941 25103 8999 25109
rect 13630 25100 13636 25152
rect 13688 25140 13694 25152
rect 13832 25140 13860 25180
rect 14093 25177 14105 25180
rect 14139 25208 14151 25211
rect 15930 25208 15936 25220
rect 14139 25180 15936 25208
rect 14139 25177 14151 25180
rect 14093 25171 14151 25177
rect 15930 25168 15936 25180
rect 15988 25168 15994 25220
rect 16206 25168 16212 25220
rect 16264 25208 16270 25220
rect 16960 25208 16988 25248
rect 17313 25245 17325 25248
rect 17359 25245 17371 25279
rect 17420 25276 17448 25316
rect 18782 25304 18788 25356
rect 18840 25344 18846 25356
rect 19242 25344 19248 25356
rect 18840 25316 19248 25344
rect 18840 25304 18846 25316
rect 19242 25304 19248 25316
rect 19300 25344 19306 25356
rect 22204 25353 22232 25452
rect 23753 25415 23811 25421
rect 23753 25381 23765 25415
rect 23799 25381 23811 25415
rect 23753 25375 23811 25381
rect 22189 25347 22247 25353
rect 19300 25316 20760 25344
rect 19300 25304 19306 25316
rect 20732 25285 20760 25316
rect 22189 25313 22201 25347
rect 22235 25313 22247 25347
rect 22189 25307 22247 25313
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 17420 25248 19625 25276
rect 17313 25239 17371 25245
rect 16264 25180 16988 25208
rect 17037 25211 17095 25217
rect 16264 25168 16270 25180
rect 17037 25177 17049 25211
rect 17083 25177 17095 25211
rect 17328 25208 17356 25239
rect 17880 25220 17908 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25276 20775 25279
rect 21358 25276 21364 25288
rect 20763 25248 21364 25276
rect 20763 25245 20775 25248
rect 20717 25239 20775 25245
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 17402 25208 17408 25220
rect 17328 25180 17408 25208
rect 17037 25171 17095 25177
rect 13688 25112 13860 25140
rect 13688 25100 13694 25112
rect 13906 25100 13912 25152
rect 13964 25100 13970 25152
rect 14642 25100 14648 25152
rect 14700 25100 14706 25152
rect 16761 25143 16819 25149
rect 16761 25109 16773 25143
rect 16807 25140 16819 25143
rect 16942 25140 16948 25152
rect 16807 25112 16948 25140
rect 16807 25109 16819 25112
rect 16761 25103 16819 25109
rect 16942 25100 16948 25112
rect 17000 25140 17006 25152
rect 17052 25140 17080 25171
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 17580 25211 17638 25217
rect 17580 25177 17592 25211
rect 17626 25208 17638 25211
rect 17770 25208 17776 25220
rect 17626 25180 17776 25208
rect 17626 25177 17638 25180
rect 17580 25171 17638 25177
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 17862 25168 17868 25220
rect 17920 25168 17926 25220
rect 19429 25211 19487 25217
rect 19429 25177 19441 25211
rect 19475 25177 19487 25211
rect 19429 25171 19487 25177
rect 20984 25211 21042 25217
rect 20984 25177 20996 25211
rect 21030 25208 21042 25211
rect 21266 25208 21272 25220
rect 21030 25180 21272 25208
rect 21030 25177 21042 25180
rect 20984 25171 21042 25177
rect 17000 25112 17080 25140
rect 17221 25143 17279 25149
rect 17000 25100 17006 25112
rect 17221 25109 17233 25143
rect 17267 25140 17279 25143
rect 17954 25140 17960 25152
rect 17267 25112 17960 25140
rect 17267 25109 17279 25112
rect 17221 25103 17279 25109
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 18693 25143 18751 25149
rect 18693 25109 18705 25143
rect 18739 25140 18751 25143
rect 18874 25140 18880 25152
rect 18739 25112 18880 25140
rect 18739 25109 18751 25112
rect 18693 25103 18751 25109
rect 18874 25100 18880 25112
rect 18932 25140 18938 25152
rect 19444 25140 19472 25171
rect 21266 25168 21272 25180
rect 21324 25168 21330 25220
rect 22462 25217 22468 25220
rect 22456 25171 22468 25217
rect 22462 25168 22468 25171
rect 22520 25168 22526 25220
rect 23768 25208 23796 25375
rect 24412 25288 24440 25452
rect 25774 25440 25780 25492
rect 25832 25440 25838 25492
rect 24394 25236 24400 25288
rect 24452 25236 24458 25288
rect 23584 25180 23796 25208
rect 18932 25112 19472 25140
rect 22097 25143 22155 25149
rect 18932 25100 18938 25112
rect 22097 25109 22109 25143
rect 22143 25140 22155 25143
rect 22370 25140 22376 25152
rect 22143 25112 22376 25140
rect 22143 25109 22155 25112
rect 22097 25103 22155 25109
rect 22370 25100 22376 25112
rect 22428 25100 22434 25152
rect 23584 25149 23612 25180
rect 23768 25152 23796 25180
rect 24118 25168 24124 25220
rect 24176 25168 24182 25220
rect 24302 25168 24308 25220
rect 24360 25208 24366 25220
rect 24642 25211 24700 25217
rect 24642 25208 24654 25211
rect 24360 25180 24654 25208
rect 24360 25168 24366 25180
rect 24642 25177 24654 25180
rect 24688 25177 24700 25211
rect 24642 25171 24700 25177
rect 23569 25143 23627 25149
rect 23569 25109 23581 25143
rect 23615 25109 23627 25143
rect 23569 25103 23627 25109
rect 23658 25100 23664 25152
rect 23716 25100 23722 25152
rect 23750 25100 23756 25152
rect 23808 25100 23814 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4525 24939 4583 24945
rect 4525 24936 4537 24939
rect 4212 24908 4537 24936
rect 4212 24896 4218 24908
rect 4525 24905 4537 24908
rect 4571 24905 4583 24939
rect 4525 24899 4583 24905
rect 4893 24939 4951 24945
rect 4893 24905 4905 24939
rect 4939 24936 4951 24939
rect 6546 24936 6552 24948
rect 4939 24908 6552 24936
rect 4939 24905 4951 24908
rect 4893 24899 4951 24905
rect 6546 24896 6552 24908
rect 6604 24896 6610 24948
rect 6638 24896 6644 24948
rect 6696 24896 6702 24948
rect 7374 24896 7380 24948
rect 7432 24936 7438 24948
rect 8205 24939 8263 24945
rect 8205 24936 8217 24939
rect 7432 24908 8217 24936
rect 7432 24896 7438 24908
rect 8205 24905 8217 24908
rect 8251 24905 8263 24939
rect 9858 24936 9864 24948
rect 8205 24899 8263 24905
rect 8404 24908 9864 24936
rect 2222 24828 2228 24880
rect 2280 24828 2286 24880
rect 2409 24871 2467 24877
rect 2409 24837 2421 24871
rect 2455 24837 2467 24871
rect 2409 24831 2467 24837
rect 4816 24840 5028 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 1949 24803 2007 24809
rect 1949 24800 1961 24803
rect 1719 24772 1961 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 1949 24769 1961 24772
rect 1995 24769 2007 24803
rect 2424 24800 2452 24831
rect 2498 24800 2504 24812
rect 2424 24772 2504 24800
rect 1949 24763 2007 24769
rect 2498 24760 2504 24772
rect 2556 24760 2562 24812
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 2700 24732 2728 24763
rect 1872 24704 2728 24732
rect 1872 24673 1900 24704
rect 1857 24667 1915 24673
rect 1857 24633 1869 24667
rect 1903 24633 1915 24667
rect 1857 24627 1915 24633
rect 2314 24624 2320 24676
rect 2372 24664 2378 24676
rect 2866 24664 2872 24676
rect 2372 24636 2872 24664
rect 2372 24624 2378 24636
rect 2866 24624 2872 24636
rect 2924 24664 2930 24676
rect 4816 24664 4844 24840
rect 5000 24800 5028 24840
rect 5258 24828 5264 24880
rect 5316 24868 5322 24880
rect 6454 24868 6460 24880
rect 5316 24840 6460 24868
rect 5316 24828 5322 24840
rect 6454 24828 6460 24840
rect 6512 24828 6518 24880
rect 6656 24868 6684 24896
rect 7282 24868 7288 24880
rect 6564 24840 6684 24868
rect 6748 24840 7288 24868
rect 5629 24803 5687 24809
rect 5000 24772 5580 24800
rect 4982 24692 4988 24744
rect 5040 24692 5046 24744
rect 5169 24735 5227 24741
rect 5169 24701 5181 24735
rect 5215 24701 5227 24735
rect 5169 24695 5227 24701
rect 2924 24636 4844 24664
rect 2924 24624 2930 24636
rect 1486 24556 1492 24608
rect 1544 24596 1550 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 1544 24568 2237 24596
rect 1544 24556 1550 24568
rect 2225 24565 2237 24568
rect 2271 24596 2283 24599
rect 2774 24596 2780 24608
rect 2271 24568 2780 24596
rect 2271 24565 2283 24568
rect 2225 24559 2283 24565
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 3973 24599 4031 24605
rect 3973 24596 3985 24599
rect 3476 24568 3985 24596
rect 3476 24556 3482 24568
rect 3973 24565 3985 24568
rect 4019 24565 4031 24599
rect 3973 24559 4031 24565
rect 4062 24556 4068 24608
rect 4120 24596 4126 24608
rect 4706 24596 4712 24608
rect 4120 24568 4712 24596
rect 4120 24556 4126 24568
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 4890 24556 4896 24608
rect 4948 24596 4954 24608
rect 5184 24596 5212 24695
rect 5552 24608 5580 24772
rect 5629 24769 5641 24803
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 5721 24803 5779 24809
rect 5721 24769 5733 24803
rect 5767 24769 5779 24803
rect 5721 24763 5779 24769
rect 4948 24568 5212 24596
rect 4948 24556 4954 24568
rect 5442 24556 5448 24608
rect 5500 24556 5506 24608
rect 5534 24556 5540 24608
rect 5592 24556 5598 24608
rect 5644 24596 5672 24763
rect 5736 24732 5764 24763
rect 5810 24760 5816 24812
rect 5868 24800 5874 24812
rect 5905 24803 5963 24809
rect 5905 24800 5917 24803
rect 5868 24772 5917 24800
rect 5868 24760 5874 24772
rect 5905 24769 5917 24772
rect 5951 24769 5963 24803
rect 5905 24763 5963 24769
rect 5997 24803 6055 24809
rect 5997 24769 6009 24803
rect 6043 24800 6055 24803
rect 6270 24800 6276 24812
rect 6043 24772 6276 24800
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 6564 24809 6592 24840
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 6748 24800 6776 24840
rect 7282 24828 7288 24840
rect 7340 24868 7346 24880
rect 7340 24840 7512 24868
rect 7340 24828 7346 24840
rect 7484 24812 7512 24840
rect 6687 24772 6776 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 6822 24760 6828 24812
rect 6880 24760 6886 24812
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24800 6975 24803
rect 7006 24800 7012 24812
rect 6963 24772 7012 24800
rect 6963 24769 6975 24772
rect 6917 24763 6975 24769
rect 7006 24760 7012 24772
rect 7064 24760 7070 24812
rect 7190 24760 7196 24812
rect 7248 24800 7254 24812
rect 7248 24772 7420 24800
rect 7248 24760 7254 24772
rect 6365 24735 6423 24741
rect 6365 24732 6377 24735
rect 5736 24704 6377 24732
rect 6365 24701 6377 24704
rect 6411 24701 6423 24735
rect 6840 24732 6868 24760
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 6840 24704 7297 24732
rect 6365 24695 6423 24701
rect 7285 24701 7297 24704
rect 7331 24701 7343 24735
rect 7392 24732 7420 24772
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 8404 24809 8432 24908
rect 9858 24896 9864 24908
rect 9916 24936 9922 24948
rect 9916 24908 10732 24936
rect 9916 24896 9922 24908
rect 8570 24828 8576 24880
rect 8628 24828 8634 24880
rect 8846 24828 8852 24880
rect 8904 24868 8910 24880
rect 9306 24868 9312 24880
rect 8904 24840 9312 24868
rect 8904 24828 8910 24840
rect 9306 24828 9312 24840
rect 9364 24828 9370 24880
rect 10318 24828 10324 24880
rect 10376 24868 10382 24880
rect 10597 24871 10655 24877
rect 10597 24868 10609 24871
rect 10376 24840 10609 24868
rect 10376 24828 10382 24840
rect 10597 24837 10609 24840
rect 10643 24837 10655 24871
rect 10597 24831 10655 24837
rect 8389 24803 8447 24809
rect 8389 24769 8401 24803
rect 8435 24769 8447 24803
rect 8389 24763 8447 24769
rect 8481 24803 8539 24809
rect 8481 24769 8493 24803
rect 8527 24800 8539 24803
rect 8588 24800 8616 24828
rect 8527 24772 8616 24800
rect 8665 24803 8723 24809
rect 8527 24769 8539 24772
rect 8481 24763 8539 24769
rect 8665 24769 8677 24803
rect 8711 24800 8723 24803
rect 9030 24800 9036 24812
rect 8711 24772 9036 24800
rect 8711 24769 8723 24772
rect 8665 24763 8723 24769
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 9490 24800 9496 24812
rect 9447 24772 9496 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 7745 24735 7803 24741
rect 7745 24732 7757 24735
rect 7392 24704 7757 24732
rect 7285 24695 7343 24701
rect 7745 24701 7757 24704
rect 7791 24701 7803 24735
rect 7745 24695 7803 24701
rect 8570 24692 8576 24744
rect 8628 24732 8634 24744
rect 8846 24732 8852 24744
rect 8628 24704 8852 24732
rect 8628 24692 8634 24704
rect 8846 24692 8852 24704
rect 8904 24692 8910 24744
rect 9140 24732 9168 24763
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 10045 24803 10103 24809
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10137 24763 10195 24769
rect 9769 24735 9827 24741
rect 9769 24732 9781 24735
rect 9140 24704 9781 24732
rect 9769 24701 9781 24704
rect 9815 24701 9827 24735
rect 9769 24695 9827 24701
rect 7469 24667 7527 24673
rect 7469 24633 7481 24667
rect 7515 24664 7527 24667
rect 7558 24664 7564 24676
rect 7515 24636 7564 24664
rect 7515 24633 7527 24636
rect 7469 24627 7527 24633
rect 7558 24624 7564 24636
rect 7616 24664 7622 24676
rect 8941 24667 8999 24673
rect 8941 24664 8953 24667
rect 7616 24636 8953 24664
rect 7616 24624 7622 24636
rect 8941 24633 8953 24636
rect 8987 24633 8999 24667
rect 10060 24664 10088 24763
rect 10152 24732 10180 24763
rect 10226 24760 10232 24812
rect 10284 24760 10290 24812
rect 10410 24760 10416 24812
rect 10468 24760 10474 24812
rect 10502 24760 10508 24812
rect 10560 24760 10566 24812
rect 10704 24800 10732 24908
rect 11882 24896 11888 24948
rect 11940 24936 11946 24948
rect 12161 24939 12219 24945
rect 12161 24936 12173 24939
rect 11940 24908 12173 24936
rect 11940 24896 11946 24908
rect 12161 24905 12173 24908
rect 12207 24905 12219 24939
rect 12161 24899 12219 24905
rect 17770 24896 17776 24948
rect 17828 24896 17834 24948
rect 17954 24896 17960 24948
rect 18012 24896 18018 24948
rect 21266 24896 21272 24948
rect 21324 24896 21330 24948
rect 22462 24896 22468 24948
rect 22520 24896 22526 24948
rect 23658 24896 23664 24948
rect 23716 24896 23722 24948
rect 23937 24939 23995 24945
rect 23937 24905 23949 24939
rect 23983 24936 23995 24939
rect 24302 24936 24308 24948
rect 23983 24908 24308 24936
rect 23983 24905 23995 24908
rect 23937 24899 23995 24905
rect 24302 24896 24308 24908
rect 24360 24896 24366 24948
rect 10778 24828 10784 24880
rect 10836 24877 10842 24880
rect 10836 24871 10855 24877
rect 10843 24837 10855 24871
rect 10836 24831 10855 24837
rect 14268 24871 14326 24877
rect 14268 24837 14280 24871
rect 14314 24868 14326 24871
rect 14642 24868 14648 24880
rect 14314 24840 14648 24868
rect 14314 24837 14326 24840
rect 14268 24831 14326 24837
rect 10836 24828 10842 24831
rect 14642 24828 14648 24840
rect 14700 24828 14706 24880
rect 16592 24840 16804 24868
rect 16592 24812 16620 24840
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 10704 24772 11529 24800
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 10520 24732 10548 24760
rect 11716 24732 11744 24763
rect 11882 24760 11888 24812
rect 11940 24800 11946 24812
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11940 24772 12081 24800
rect 11940 24760 11946 24772
rect 12069 24769 12081 24772
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 12342 24760 12348 24812
rect 12400 24760 12406 24812
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 12986 24800 12992 24812
rect 12492 24772 12992 24800
rect 12492 24760 12498 24772
rect 12986 24760 12992 24772
rect 13044 24800 13050 24812
rect 14001 24803 14059 24809
rect 14001 24800 14013 24803
rect 13044 24772 14013 24800
rect 13044 24760 13050 24772
rect 14001 24769 14013 24772
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 16574 24760 16580 24812
rect 16632 24760 16638 24812
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16776 24800 16804 24840
rect 16942 24828 16948 24880
rect 17000 24828 17006 24880
rect 16850 24800 16856 24812
rect 16776 24772 16856 24800
rect 16669 24763 16727 24769
rect 12360 24732 12388 24760
rect 10152 24704 10548 24732
rect 10980 24704 12388 24732
rect 10980 24673 11008 24704
rect 15930 24692 15936 24744
rect 15988 24692 15994 24744
rect 8941 24627 8999 24633
rect 9784 24636 10088 24664
rect 10965 24667 11023 24673
rect 9784 24608 9812 24636
rect 10965 24633 10977 24667
rect 11011 24633 11023 24667
rect 10965 24627 11023 24633
rect 15381 24667 15439 24673
rect 15381 24633 15393 24667
rect 15427 24664 15439 24667
rect 15657 24667 15715 24673
rect 15657 24664 15669 24667
rect 15427 24636 15669 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 15657 24633 15669 24636
rect 15703 24664 15715 24667
rect 16684 24664 16712 24763
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 15703 24636 16712 24664
rect 15703 24633 15715 24636
rect 15657 24627 15715 24633
rect 7650 24596 7656 24608
rect 5644 24568 7656 24596
rect 7650 24556 7656 24568
rect 7708 24556 7714 24608
rect 9766 24556 9772 24608
rect 9824 24556 9830 24608
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10008 24568 10793 24596
rect 10008 24556 10014 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 15470 24556 15476 24608
rect 15528 24556 15534 24608
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 17052 24596 17080 24763
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 17184 24772 17325 24800
rect 17184 24760 17190 24772
rect 17313 24769 17325 24772
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 17494 24760 17500 24812
rect 17552 24760 17558 24812
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24800 17739 24803
rect 17862 24800 17868 24812
rect 17727 24772 17868 24800
rect 17727 24769 17739 24772
rect 17681 24763 17739 24769
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 17972 24809 18000 24896
rect 19076 24840 19656 24868
rect 17957 24803 18015 24809
rect 17957 24769 17969 24803
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 18966 24760 18972 24812
rect 19024 24760 19030 24812
rect 19076 24732 19104 24840
rect 19501 24803 19559 24809
rect 19501 24800 19513 24803
rect 17144 24704 19104 24732
rect 19168 24772 19513 24800
rect 17144 24608 17172 24704
rect 19168 24673 19196 24772
rect 19501 24769 19513 24772
rect 19547 24769 19559 24803
rect 19628 24800 19656 24840
rect 20806 24828 20812 24880
rect 20864 24868 20870 24880
rect 21821 24871 21879 24877
rect 21821 24868 21833 24871
rect 20864 24840 21833 24868
rect 20864 24828 20870 24840
rect 21821 24837 21833 24840
rect 21867 24837 21879 24871
rect 21821 24831 21879 24837
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 19628 24772 20729 24800
rect 19501 24763 19559 24769
rect 20717 24769 20729 24772
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 21453 24803 21511 24809
rect 21453 24769 21465 24803
rect 21499 24769 21511 24803
rect 21453 24763 21511 24769
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22189 24803 22247 24809
rect 22189 24769 22201 24803
rect 22235 24800 22247 24803
rect 22281 24803 22339 24809
rect 22281 24800 22293 24803
rect 22235 24772 22293 24800
rect 22235 24769 22247 24772
rect 22189 24763 22247 24769
rect 22281 24769 22293 24772
rect 22327 24769 22339 24803
rect 23676 24800 23704 24896
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 23676 24772 23765 24800
rect 22281 24763 22339 24769
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 23753 24763 23811 24769
rect 19242 24692 19248 24744
rect 19300 24692 19306 24744
rect 20732 24732 20760 24763
rect 21177 24735 21235 24741
rect 20732 24704 21128 24732
rect 19153 24667 19211 24673
rect 19153 24633 19165 24667
rect 19199 24633 19211 24667
rect 19153 24627 19211 24633
rect 20993 24667 21051 24673
rect 20993 24633 21005 24667
rect 21039 24633 21051 24667
rect 21100 24664 21128 24704
rect 21177 24701 21189 24735
rect 21223 24732 21235 24735
rect 21468 24732 21496 24763
rect 21223 24704 21496 24732
rect 22020 24732 22048 24763
rect 22370 24732 22376 24744
rect 22020 24704 22376 24732
rect 21223 24701 21235 24704
rect 21177 24695 21235 24701
rect 22370 24692 22376 24704
rect 22428 24692 22434 24744
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 25130 24732 25136 24744
rect 24176 24704 25136 24732
rect 24176 24692 24182 24704
rect 25130 24692 25136 24704
rect 25188 24732 25194 24744
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 25188 24704 25237 24732
rect 25188 24692 25194 24704
rect 25225 24701 25237 24704
rect 25271 24701 25283 24735
rect 25225 24695 25283 24701
rect 24136 24664 24164 24692
rect 21100 24636 24164 24664
rect 20993 24627 21051 24633
rect 16172 24568 17080 24596
rect 16172 24556 16178 24568
rect 17126 24556 17132 24608
rect 17184 24556 17190 24608
rect 17218 24556 17224 24608
rect 17276 24556 17282 24608
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 20625 24599 20683 24605
rect 20625 24596 20637 24599
rect 19576 24568 20637 24596
rect 19576 24556 19582 24568
rect 20625 24565 20637 24568
rect 20671 24596 20683 24599
rect 21008 24596 21036 24627
rect 24946 24624 24952 24676
rect 25004 24624 25010 24676
rect 20671 24568 21036 24596
rect 20671 24565 20683 24568
rect 20625 24559 20683 24565
rect 24762 24556 24768 24608
rect 24820 24556 24826 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 2590 24352 2596 24404
rect 2648 24352 2654 24404
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3513 24395 3571 24401
rect 3513 24392 3525 24395
rect 3384 24364 3525 24392
rect 3384 24352 3390 24364
rect 3513 24361 3525 24364
rect 3559 24361 3571 24395
rect 3513 24355 3571 24361
rect 4893 24395 4951 24401
rect 4893 24361 4905 24395
rect 4939 24392 4951 24395
rect 4982 24392 4988 24404
rect 4939 24364 4988 24392
rect 4939 24361 4951 24364
rect 4893 24355 4951 24361
rect 4982 24352 4988 24364
rect 5040 24352 5046 24404
rect 5184 24364 6040 24392
rect 2314 24284 2320 24336
rect 2372 24284 2378 24336
rect 3160 24296 3924 24324
rect 1394 24216 1400 24268
rect 1452 24216 1458 24268
rect 2332 24256 2360 24284
rect 2240 24228 2360 24256
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 1857 24151 1915 24157
rect 1872 24120 1900 24151
rect 1946 24148 1952 24200
rect 2004 24188 2010 24200
rect 2240 24197 2268 24228
rect 2774 24216 2780 24268
rect 2832 24216 2838 24268
rect 3160 24265 3188 24296
rect 3896 24268 3924 24296
rect 3145 24259 3203 24265
rect 3145 24225 3157 24259
rect 3191 24225 3203 24259
rect 3145 24219 3203 24225
rect 3234 24216 3240 24268
rect 3292 24256 3298 24268
rect 3605 24259 3663 24265
rect 3292 24228 3556 24256
rect 3292 24216 3298 24228
rect 2225 24191 2283 24197
rect 2225 24188 2237 24191
rect 2004 24160 2237 24188
rect 2004 24148 2010 24160
rect 2225 24157 2237 24160
rect 2271 24157 2283 24191
rect 2225 24151 2283 24157
rect 2314 24148 2320 24200
rect 2372 24148 2378 24200
rect 2792 24188 2820 24216
rect 3329 24191 3387 24197
rect 3329 24188 3341 24191
rect 2792 24160 3341 24188
rect 3329 24157 3341 24160
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24157 3479 24191
rect 3528 24188 3556 24228
rect 3605 24225 3617 24259
rect 3651 24256 3663 24259
rect 3694 24256 3700 24268
rect 3651 24228 3700 24256
rect 3651 24225 3663 24228
rect 3605 24219 3663 24225
rect 3694 24216 3700 24228
rect 3752 24216 3758 24268
rect 3878 24216 3884 24268
rect 3936 24216 3942 24268
rect 4433 24259 4491 24265
rect 4433 24225 4445 24259
rect 4479 24256 4491 24259
rect 4890 24256 4896 24268
rect 4479 24228 4896 24256
rect 4479 24225 4491 24228
rect 4433 24219 4491 24225
rect 4890 24216 4896 24228
rect 4948 24216 4954 24268
rect 5077 24191 5135 24197
rect 3528 24160 4476 24188
rect 3421 24151 3479 24157
rect 2774 24120 2780 24132
rect 1872 24092 2780 24120
rect 2774 24080 2780 24092
rect 2832 24080 2838 24132
rect 2869 24123 2927 24129
rect 2869 24089 2881 24123
rect 2915 24120 2927 24123
rect 2958 24120 2964 24132
rect 2915 24092 2964 24120
rect 2915 24089 2927 24092
rect 2869 24083 2927 24089
rect 2958 24080 2964 24092
rect 3016 24080 3022 24132
rect 3142 24080 3148 24132
rect 3200 24120 3206 24132
rect 3436 24120 3464 24151
rect 4338 24120 4344 24132
rect 3200 24092 3464 24120
rect 4172 24092 4344 24120
rect 3200 24080 3206 24092
rect 4172 24061 4200 24092
rect 4338 24080 4344 24092
rect 4396 24080 4402 24132
rect 3053 24055 3111 24061
rect 3053 24021 3065 24055
rect 3099 24052 3111 24055
rect 3789 24055 3847 24061
rect 3789 24052 3801 24055
rect 3099 24024 3801 24052
rect 3099 24021 3111 24024
rect 3053 24015 3111 24021
rect 3789 24021 3801 24024
rect 3835 24021 3847 24055
rect 3789 24015 3847 24021
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24021 4215 24055
rect 4157 24015 4215 24021
rect 4246 24012 4252 24064
rect 4304 24012 4310 24064
rect 4448 24052 4476 24160
rect 5077 24157 5089 24191
rect 5123 24188 5135 24191
rect 5184 24188 5212 24364
rect 6012 24336 6040 24364
rect 9582 24352 9588 24404
rect 9640 24392 9646 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 9640 24364 10057 24392
rect 9640 24352 9646 24364
rect 10045 24361 10057 24364
rect 10091 24361 10103 24395
rect 10045 24355 10103 24361
rect 15470 24352 15476 24404
rect 15528 24352 15534 24404
rect 15657 24395 15715 24401
rect 15657 24361 15669 24395
rect 15703 24392 15715 24395
rect 15746 24392 15752 24404
rect 15703 24364 15752 24392
rect 15703 24361 15715 24364
rect 15657 24355 15715 24361
rect 15746 24352 15752 24364
rect 15804 24352 15810 24404
rect 16132 24364 18276 24392
rect 5442 24324 5448 24336
rect 5276 24296 5448 24324
rect 5276 24197 5304 24296
rect 5442 24284 5448 24296
rect 5500 24284 5506 24336
rect 5994 24284 6000 24336
rect 6052 24284 6058 24336
rect 6181 24327 6239 24333
rect 6181 24293 6193 24327
rect 6227 24293 6239 24327
rect 6181 24287 6239 24293
rect 6917 24327 6975 24333
rect 6917 24293 6929 24327
rect 6963 24293 6975 24327
rect 6917 24287 6975 24293
rect 6196 24256 6224 24287
rect 5460 24228 6224 24256
rect 5123 24160 5212 24188
rect 5261 24191 5319 24197
rect 5123 24157 5135 24160
rect 5077 24151 5135 24157
rect 5261 24157 5273 24191
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 5350 24148 5356 24200
rect 5408 24188 5414 24200
rect 5460 24197 5488 24228
rect 6822 24216 6828 24268
rect 6880 24216 6886 24268
rect 6932 24256 6960 24287
rect 10778 24284 10784 24336
rect 10836 24284 10842 24336
rect 13541 24327 13599 24333
rect 13541 24293 13553 24327
rect 13587 24324 13599 24327
rect 13906 24324 13912 24336
rect 13587 24296 13912 24324
rect 13587 24293 13599 24296
rect 13541 24287 13599 24293
rect 13906 24284 13912 24296
rect 13964 24284 13970 24336
rect 6932 24228 7512 24256
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5408 24160 5457 24188
rect 5408 24148 5414 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 5445 24151 5503 24157
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24157 5963 24191
rect 5905 24151 5963 24157
rect 5169 24123 5227 24129
rect 5169 24089 5181 24123
rect 5215 24120 5227 24123
rect 5920 24120 5948 24151
rect 6086 24148 6092 24200
rect 6144 24148 6150 24200
rect 6362 24148 6368 24200
rect 6420 24188 6426 24200
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 6420 24160 6469 24188
rect 6420 24148 6426 24160
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 6840 24188 6868 24216
rect 7484 24200 7512 24228
rect 9306 24216 9312 24268
rect 9364 24256 9370 24268
rect 10796 24256 10824 24284
rect 9364 24228 10824 24256
rect 10965 24259 11023 24265
rect 9364 24216 9370 24228
rect 6917 24191 6975 24197
rect 6917 24188 6929 24191
rect 6840 24160 6929 24188
rect 6457 24151 6515 24157
rect 6917 24157 6929 24160
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 7006 24148 7012 24200
rect 7064 24148 7070 24200
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24188 7251 24191
rect 7374 24188 7380 24200
rect 7239 24160 7380 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 7466 24148 7472 24200
rect 7524 24148 7530 24200
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24157 7711 24191
rect 7653 24151 7711 24157
rect 5215 24092 5948 24120
rect 5215 24089 5227 24092
rect 5169 24083 5227 24089
rect 5629 24055 5687 24061
rect 5629 24052 5641 24055
rect 4448 24024 5641 24052
rect 5629 24021 5641 24024
rect 5675 24021 5687 24055
rect 5920 24052 5948 24092
rect 5994 24080 6000 24132
rect 6052 24120 6058 24132
rect 6181 24123 6239 24129
rect 6181 24120 6193 24123
rect 6052 24092 6193 24120
rect 6052 24080 6058 24092
rect 6181 24089 6193 24092
rect 6227 24089 6239 24123
rect 6181 24083 6239 24089
rect 7285 24123 7343 24129
rect 7285 24089 7297 24123
rect 7331 24089 7343 24123
rect 7392 24120 7420 24148
rect 7668 24120 7696 24151
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9585 24191 9643 24197
rect 9585 24188 9597 24191
rect 8812 24160 9597 24188
rect 8812 24148 8818 24160
rect 9585 24157 9597 24160
rect 9631 24157 9643 24191
rect 9585 24151 9643 24157
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 10229 24191 10287 24197
rect 10229 24188 10241 24191
rect 10008 24160 10241 24188
rect 10008 24148 10014 24160
rect 10229 24157 10241 24160
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 10318 24148 10324 24200
rect 10376 24148 10382 24200
rect 10428 24197 10456 24228
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11698 24256 11704 24268
rect 11011 24228 11704 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11698 24216 11704 24228
rect 11756 24216 11762 24268
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 13633 24259 13691 24265
rect 11848 24228 12296 24256
rect 11848 24216 11854 24228
rect 10876 24200 10928 24206
rect 10413 24191 10471 24197
rect 10413 24157 10425 24191
rect 10459 24157 10471 24191
rect 10413 24151 10471 24157
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 10643 24160 10732 24188
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 7392 24092 7696 24120
rect 7285 24083 7343 24089
rect 6270 24052 6276 24064
rect 5920 24024 6276 24052
rect 5629 24015 5687 24021
rect 6270 24012 6276 24024
rect 6328 24012 6334 24064
rect 6365 24055 6423 24061
rect 6365 24021 6377 24055
rect 6411 24052 6423 24055
rect 6730 24052 6736 24064
rect 6411 24024 6736 24052
rect 6411 24021 6423 24024
rect 6365 24015 6423 24021
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 7300 24052 7328 24083
rect 9030 24080 9036 24132
rect 9088 24120 9094 24132
rect 9401 24123 9459 24129
rect 9401 24120 9413 24123
rect 9088 24092 9413 24120
rect 9088 24080 9094 24092
rect 9401 24089 9413 24092
rect 9447 24089 9459 24123
rect 9401 24083 9459 24089
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10704 24120 10732 24160
rect 11882 24188 11888 24200
rect 10876 24142 10928 24148
rect 11716 24160 11888 24188
rect 9916 24092 10732 24120
rect 9916 24080 9922 24092
rect 7248 24024 7328 24052
rect 7653 24055 7711 24061
rect 7248 24012 7254 24024
rect 7653 24021 7665 24055
rect 7699 24052 7711 24055
rect 8570 24052 8576 24064
rect 7699 24024 8576 24052
rect 7699 24021 7711 24024
rect 7653 24015 7711 24021
rect 8570 24012 8576 24024
rect 8628 24012 8634 24064
rect 9769 24055 9827 24061
rect 9769 24021 9781 24055
rect 9815 24052 9827 24055
rect 10410 24052 10416 24064
rect 9815 24024 10416 24052
rect 9815 24021 9827 24024
rect 9769 24015 9827 24021
rect 10410 24012 10416 24024
rect 10468 24012 10474 24064
rect 10704 24052 10732 24092
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 11716 24120 11744 24160
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 12268 24197 12296 24228
rect 13633 24225 13645 24259
rect 13679 24256 13691 24259
rect 13679 24228 13952 24256
rect 13679 24225 13691 24228
rect 13633 24219 13691 24225
rect 12253 24191 12311 24197
rect 12253 24157 12265 24191
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 13924 24197 13952 24228
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12400 24160 12541 24188
rect 12400 24148 12406 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 13909 24191 13967 24197
rect 13909 24157 13921 24191
rect 13955 24157 13967 24191
rect 13909 24151 13967 24157
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15488 24188 15516 24352
rect 15562 24216 15568 24268
rect 15620 24256 15626 24268
rect 15620 24228 15684 24256
rect 15620 24216 15626 24228
rect 15151 24160 15516 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 11296 24092 11744 24120
rect 12161 24123 12219 24129
rect 11296 24080 11302 24092
rect 12161 24089 12173 24123
rect 12207 24089 12219 24123
rect 12161 24083 12219 24089
rect 12176 24052 12204 24083
rect 13078 24080 13084 24132
rect 13136 24120 13142 24132
rect 13173 24123 13231 24129
rect 13173 24120 13185 24123
rect 13136 24092 13185 24120
rect 13136 24080 13142 24092
rect 13173 24089 13185 24092
rect 13219 24089 13231 24123
rect 13173 24083 13231 24089
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 14642 24120 14648 24132
rect 14516 24092 14648 24120
rect 14516 24080 14522 24092
rect 14642 24080 14648 24092
rect 14700 24120 14706 24132
rect 15656 24129 15684 24228
rect 15641 24123 15699 24129
rect 14700 24092 15608 24120
rect 14700 24080 14706 24092
rect 10704 24024 12204 24052
rect 13722 24012 13728 24064
rect 13780 24012 13786 24064
rect 14921 24055 14979 24061
rect 14921 24021 14933 24055
rect 14967 24052 14979 24055
rect 15286 24052 15292 24064
rect 14967 24024 15292 24052
rect 14967 24021 14979 24024
rect 14921 24015 14979 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 15470 24012 15476 24064
rect 15528 24012 15534 24064
rect 15580 24052 15608 24092
rect 15641 24089 15653 24123
rect 15687 24089 15699 24123
rect 15641 24083 15699 24089
rect 15841 24123 15899 24129
rect 15841 24089 15853 24123
rect 15887 24120 15899 24123
rect 16132 24120 16160 24364
rect 18248 24324 18276 24364
rect 18966 24352 18972 24404
rect 19024 24392 19030 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 19024 24364 19257 24392
rect 19024 24352 19030 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 21082 24324 21088 24336
rect 18248 24296 21088 24324
rect 21082 24284 21088 24296
rect 21140 24284 21146 24336
rect 23385 24327 23443 24333
rect 23385 24293 23397 24327
rect 23431 24293 23443 24327
rect 23385 24287 23443 24293
rect 19242 24216 19248 24268
rect 19300 24216 19306 24268
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 17402 24188 17408 24200
rect 17359 24160 17408 24188
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 17402 24148 17408 24160
rect 17460 24188 17466 24200
rect 19260 24188 19288 24216
rect 17460 24160 19288 24188
rect 19613 24191 19671 24197
rect 17460 24148 17466 24160
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 20806 24188 20812 24200
rect 19659 24160 20812 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 20806 24148 20812 24160
rect 20864 24148 20870 24200
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24188 22707 24191
rect 23017 24191 23075 24197
rect 22695 24160 22968 24188
rect 22695 24157 22707 24160
rect 22649 24151 22707 24157
rect 17586 24129 17592 24132
rect 15887 24092 16160 24120
rect 15887 24089 15899 24092
rect 15841 24083 15899 24089
rect 17580 24083 17592 24129
rect 15856 24052 15884 24083
rect 17586 24080 17592 24083
rect 17644 24080 17650 24132
rect 18782 24120 18788 24132
rect 18708 24092 18788 24120
rect 18708 24061 18736 24092
rect 18782 24080 18788 24092
rect 18840 24120 18846 24132
rect 19429 24123 19487 24129
rect 19429 24120 19441 24123
rect 18840 24092 19441 24120
rect 18840 24080 18846 24092
rect 19429 24089 19441 24092
rect 19475 24089 19487 24123
rect 19429 24083 19487 24089
rect 22738 24080 22744 24132
rect 22796 24080 22802 24132
rect 22830 24080 22836 24132
rect 22888 24080 22894 24132
rect 15580 24024 15884 24052
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24021 18751 24055
rect 18693 24015 18751 24021
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 22465 24055 22523 24061
rect 22465 24052 22477 24055
rect 22336 24024 22477 24052
rect 22336 24012 22342 24024
rect 22465 24021 22477 24024
rect 22511 24021 22523 24055
rect 22940 24052 22968 24160
rect 23017 24157 23029 24191
rect 23063 24188 23075 24191
rect 23198 24188 23204 24200
rect 23063 24160 23204 24188
rect 23063 24157 23075 24160
rect 23017 24151 23075 24157
rect 23198 24148 23204 24160
rect 23256 24188 23262 24200
rect 23400 24188 23428 24287
rect 23569 24259 23627 24265
rect 23569 24225 23581 24259
rect 23615 24256 23627 24259
rect 23615 24228 23704 24256
rect 23615 24225 23627 24228
rect 23569 24219 23627 24225
rect 23676 24197 23704 24228
rect 23256 24160 23428 24188
rect 23661 24191 23719 24197
rect 23256 24148 23262 24160
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 24394 24148 24400 24200
rect 24452 24148 24458 24200
rect 23109 24123 23167 24129
rect 23109 24089 23121 24123
rect 23155 24120 23167 24123
rect 23290 24120 23296 24132
rect 23155 24092 23296 24120
rect 23155 24089 23167 24092
rect 23109 24083 23167 24089
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 24642 24123 24700 24129
rect 24642 24120 24654 24123
rect 23860 24092 24654 24120
rect 23014 24052 23020 24064
rect 22940 24024 23020 24052
rect 22465 24015 22523 24021
rect 23014 24012 23020 24024
rect 23072 24012 23078 24064
rect 23860 24061 23888 24092
rect 24642 24089 24654 24092
rect 24688 24089 24700 24123
rect 24642 24083 24700 24089
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24021 23903 24055
rect 23845 24015 23903 24021
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25777 24055 25835 24061
rect 25777 24052 25789 24055
rect 25004 24024 25789 24052
rect 25004 24012 25010 24024
rect 25777 24021 25789 24024
rect 25823 24021 25835 24055
rect 25777 24015 25835 24021
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 2222 23808 2228 23860
rect 2280 23808 2286 23860
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 2832 23820 3617 23848
rect 2832 23808 2838 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 3605 23811 3663 23817
rect 4246 23808 4252 23860
rect 4304 23848 4310 23860
rect 4525 23851 4583 23857
rect 4525 23848 4537 23851
rect 4304 23820 4537 23848
rect 4304 23808 4310 23820
rect 4525 23817 4537 23820
rect 4571 23817 4583 23851
rect 4525 23811 4583 23817
rect 4709 23851 4767 23857
rect 4709 23817 4721 23851
rect 4755 23848 4767 23851
rect 5353 23851 5411 23857
rect 5353 23848 5365 23851
rect 4755 23820 5365 23848
rect 4755 23817 4767 23820
rect 4709 23811 4767 23817
rect 5353 23817 5365 23820
rect 5399 23817 5411 23851
rect 5353 23811 5411 23817
rect 5810 23808 5816 23860
rect 5868 23848 5874 23860
rect 5994 23848 6000 23860
rect 5868 23820 6000 23848
rect 5868 23808 5874 23820
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6730 23808 6736 23860
rect 6788 23808 6794 23860
rect 7392 23820 9352 23848
rect 1946 23672 1952 23724
rect 2004 23672 2010 23724
rect 2130 23672 2136 23724
rect 2188 23672 2194 23724
rect 2240 23721 2268 23808
rect 2682 23740 2688 23792
rect 2740 23780 2746 23792
rect 2740 23752 4016 23780
rect 2740 23740 2746 23752
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2314 23672 2320 23724
rect 2372 23672 2378 23724
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23681 2559 23715
rect 3142 23712 3148 23724
rect 2501 23675 2559 23681
rect 2746 23684 3148 23712
rect 2332 23644 2360 23672
rect 2240 23616 2360 23644
rect 2240 23520 2268 23616
rect 2516 23588 2544 23675
rect 2498 23536 2504 23588
rect 2556 23536 2562 23588
rect 2222 23468 2228 23520
rect 2280 23468 2286 23520
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2746 23508 2774 23684
rect 3142 23672 3148 23684
rect 3200 23672 3206 23724
rect 3789 23715 3847 23721
rect 3789 23681 3801 23715
rect 3835 23712 3847 23715
rect 3878 23712 3884 23724
rect 3835 23684 3884 23712
rect 3835 23681 3847 23684
rect 3789 23675 3847 23681
rect 3142 23536 3148 23588
rect 3200 23576 3206 23588
rect 3804 23576 3832 23675
rect 3878 23672 3884 23684
rect 3936 23672 3942 23724
rect 3988 23721 4016 23752
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 4120 23752 4384 23780
rect 4120 23740 4126 23752
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23681 4031 23715
rect 3973 23675 4031 23681
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23712 4215 23715
rect 4246 23712 4252 23724
rect 4203 23684 4252 23712
rect 4203 23681 4215 23684
rect 4157 23675 4215 23681
rect 4246 23672 4252 23684
rect 4304 23672 4310 23724
rect 4356 23721 4384 23752
rect 5626 23740 5632 23792
rect 5684 23740 5690 23792
rect 5718 23740 5724 23792
rect 5776 23780 5782 23792
rect 6365 23783 6423 23789
rect 6365 23780 6377 23783
rect 5776 23752 6377 23780
rect 5776 23740 5782 23752
rect 6365 23749 6377 23752
rect 6411 23749 6423 23783
rect 6365 23743 6423 23749
rect 6638 23740 6644 23792
rect 6696 23780 6702 23792
rect 7282 23780 7288 23792
rect 6696 23752 7288 23780
rect 6696 23740 6702 23752
rect 7282 23740 7288 23752
rect 7340 23740 7346 23792
rect 4341 23715 4399 23721
rect 4341 23681 4353 23715
rect 4387 23681 4399 23715
rect 4341 23675 4399 23681
rect 4706 23715 4764 23721
rect 4706 23681 4718 23715
rect 4752 23712 4764 23715
rect 5350 23712 5356 23724
rect 4752 23684 5356 23712
rect 4752 23681 4764 23684
rect 4706 23675 4764 23681
rect 5350 23672 5356 23684
rect 5408 23672 5414 23724
rect 5644 23712 5672 23740
rect 5644 23684 5764 23712
rect 5736 23656 5764 23684
rect 6822 23672 6828 23724
rect 6880 23672 6886 23724
rect 7006 23672 7012 23724
rect 7064 23712 7070 23724
rect 7101 23715 7159 23721
rect 7101 23712 7113 23715
rect 7064 23684 7113 23712
rect 7064 23672 7070 23684
rect 7101 23681 7113 23684
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23712 7251 23715
rect 7392 23712 7420 23820
rect 9324 23792 9352 23820
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 10870 23848 10876 23860
rect 10376 23820 10876 23848
rect 10376 23808 10382 23820
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 12897 23851 12955 23857
rect 12897 23817 12909 23851
rect 12943 23848 12955 23851
rect 12986 23848 12992 23860
rect 12943 23820 12992 23848
rect 12943 23817 12955 23820
rect 12897 23811 12955 23817
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 13722 23808 13728 23860
rect 13780 23808 13786 23860
rect 16114 23808 16120 23860
rect 16172 23808 16178 23860
rect 17497 23851 17555 23857
rect 17497 23817 17509 23851
rect 17543 23848 17555 23851
rect 17586 23848 17592 23860
rect 17543 23820 17592 23848
rect 17543 23817 17555 23820
rect 17497 23811 17555 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 19813 23851 19871 23857
rect 19813 23848 19825 23851
rect 18860 23820 19825 23848
rect 9306 23740 9312 23792
rect 9364 23740 9370 23792
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 10689 23783 10747 23789
rect 10689 23780 10701 23783
rect 10192 23752 10701 23780
rect 10192 23740 10198 23752
rect 10689 23749 10701 23752
rect 10735 23780 10747 23783
rect 10962 23780 10968 23792
rect 10735 23752 10968 23780
rect 10735 23749 10747 23752
rect 10689 23743 10747 23749
rect 10962 23740 10968 23752
rect 11020 23780 11026 23792
rect 11020 23752 11192 23780
rect 11020 23740 11026 23752
rect 7239 23684 7420 23712
rect 7239 23681 7251 23684
rect 7193 23675 7251 23681
rect 4062 23604 4068 23656
rect 4120 23604 4126 23656
rect 4430 23604 4436 23656
rect 4488 23644 4494 23656
rect 4982 23644 4988 23656
rect 4488 23616 4988 23644
rect 4488 23604 4494 23616
rect 4982 23604 4988 23616
rect 5040 23604 5046 23656
rect 5166 23604 5172 23656
rect 5224 23644 5230 23656
rect 5442 23644 5448 23656
rect 5224 23616 5448 23644
rect 5224 23604 5230 23616
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 5534 23604 5540 23656
rect 5592 23604 5598 23656
rect 5626 23604 5632 23656
rect 5684 23604 5690 23656
rect 5718 23604 5724 23656
rect 5776 23604 5782 23656
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 6178 23644 6184 23656
rect 5859 23616 6184 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 6178 23604 6184 23616
rect 6236 23604 6242 23656
rect 6457 23647 6515 23653
rect 6457 23613 6469 23647
rect 6503 23644 6515 23647
rect 6730 23644 6736 23656
rect 6503 23616 6736 23644
rect 6503 23613 6515 23616
rect 6457 23607 6515 23613
rect 6730 23604 6736 23616
rect 6788 23604 6794 23656
rect 7116 23644 7144 23675
rect 7466 23672 7472 23724
rect 7524 23672 7530 23724
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 7742 23672 7748 23724
rect 7800 23672 7806 23724
rect 8297 23715 8355 23721
rect 8297 23681 8309 23715
rect 8343 23712 8355 23715
rect 8386 23712 8392 23724
rect 8343 23684 8392 23712
rect 8343 23681 8355 23684
rect 8297 23675 8355 23681
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 10042 23672 10048 23724
rect 10100 23712 10106 23724
rect 11164 23721 11192 23752
rect 10505 23715 10563 23721
rect 10505 23712 10517 23715
rect 10100 23684 10517 23712
rect 10100 23672 10106 23684
rect 10505 23681 10517 23684
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 11057 23715 11115 23721
rect 11057 23712 11069 23715
rect 10827 23684 11069 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 11057 23681 11069 23684
rect 11103 23681 11115 23715
rect 11057 23675 11115 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 7116 23616 7328 23644
rect 6917 23579 6975 23585
rect 6917 23576 6929 23579
rect 3200 23548 3832 23576
rect 3988 23548 6929 23576
rect 3200 23536 3206 23548
rect 3988 23520 4016 23548
rect 6917 23545 6929 23548
rect 6963 23545 6975 23579
rect 6917 23539 6975 23545
rect 7300 23520 7328 23616
rect 10318 23604 10324 23656
rect 10376 23644 10382 23656
rect 10796 23644 10824 23675
rect 10376 23616 10824 23644
rect 11072 23644 11100 23675
rect 12802 23672 12808 23724
rect 12860 23672 12866 23724
rect 13004 23712 13032 23808
rect 13348 23783 13406 23789
rect 13348 23749 13360 23783
rect 13394 23780 13406 23783
rect 13740 23780 13768 23808
rect 13394 23752 13768 23780
rect 14912 23783 14970 23789
rect 13394 23749 13406 23752
rect 13348 23743 13406 23749
rect 14912 23749 14924 23783
rect 14958 23780 14970 23783
rect 15286 23780 15292 23792
rect 14958 23752 15292 23780
rect 14958 23749 14970 23752
rect 14912 23743 14970 23749
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 15562 23740 15568 23792
rect 15620 23780 15626 23792
rect 18860 23789 18888 23820
rect 19813 23817 19825 23820
rect 19859 23817 19871 23851
rect 19813 23811 19871 23817
rect 21453 23851 21511 23857
rect 21453 23817 21465 23851
rect 21499 23848 21511 23851
rect 21499 23820 22094 23848
rect 21499 23817 21511 23820
rect 21453 23811 21511 23817
rect 18845 23783 18903 23789
rect 18845 23780 18857 23783
rect 15620 23752 18857 23780
rect 15620 23740 15626 23752
rect 16316 23721 16344 23752
rect 18845 23749 18857 23752
rect 18891 23749 18903 23783
rect 18845 23743 18903 23749
rect 19061 23783 19119 23789
rect 19061 23749 19073 23783
rect 19107 23780 19119 23783
rect 19613 23783 19671 23789
rect 19613 23780 19625 23783
rect 19107 23752 19625 23780
rect 19107 23749 19119 23752
rect 19061 23743 19119 23749
rect 19613 23749 19625 23752
rect 19659 23780 19671 23783
rect 19702 23780 19708 23792
rect 19659 23752 19708 23780
rect 19659 23749 19671 23752
rect 19613 23743 19671 23749
rect 19702 23740 19708 23752
rect 19760 23780 19766 23792
rect 22066 23789 22094 23820
rect 23198 23808 23204 23860
rect 23256 23808 23262 23860
rect 24762 23808 24768 23860
rect 24820 23808 24826 23860
rect 24857 23851 24915 23857
rect 24857 23817 24869 23851
rect 24903 23817 24915 23851
rect 24857 23811 24915 23817
rect 20533 23783 20591 23789
rect 20533 23780 20545 23783
rect 19760 23752 20545 23780
rect 19760 23740 19766 23752
rect 20533 23749 20545 23752
rect 20579 23749 20591 23783
rect 20533 23743 20591 23749
rect 22066 23783 22124 23789
rect 22066 23749 22078 23783
rect 22112 23749 22124 23783
rect 22066 23743 22124 23749
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 23569 23783 23627 23789
rect 23569 23780 23581 23783
rect 22980 23752 23581 23780
rect 22980 23740 22986 23752
rect 23569 23749 23581 23752
rect 23615 23749 23627 23783
rect 23569 23743 23627 23749
rect 23661 23783 23719 23789
rect 23661 23749 23673 23783
rect 23707 23749 23719 23783
rect 23661 23743 23719 23749
rect 13081 23715 13139 23721
rect 13081 23712 13093 23715
rect 13004 23684 13093 23712
rect 13081 23681 13093 23684
rect 13127 23712 13139 23715
rect 14645 23715 14703 23721
rect 14645 23712 14657 23715
rect 13127 23684 14657 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 14645 23681 14657 23684
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23681 16359 23715
rect 16301 23675 16359 23681
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 11072 23616 12112 23644
rect 10376 23604 10382 23616
rect 7466 23536 7472 23588
rect 7524 23576 7530 23588
rect 8202 23576 8208 23588
rect 7524 23548 8208 23576
rect 7524 23536 7530 23548
rect 8202 23536 8208 23548
rect 8260 23536 8266 23588
rect 12084 23520 12112 23616
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 16485 23647 16543 23653
rect 16485 23644 16497 23647
rect 16172 23616 16497 23644
rect 16172 23604 16178 23616
rect 16485 23613 16497 23616
rect 16531 23613 16543 23647
rect 16485 23607 16543 23613
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16724 23616 16773 23644
rect 16724 23604 16730 23616
rect 16761 23613 16773 23616
rect 16807 23644 16819 23647
rect 17126 23644 17132 23656
rect 16807 23616 17132 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 17221 23647 17279 23653
rect 17221 23613 17233 23647
rect 17267 23644 17279 23647
rect 17328 23644 17356 23675
rect 21266 23672 21272 23724
rect 21324 23672 21330 23724
rect 21358 23672 21364 23724
rect 21416 23712 21422 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21416 23684 21833 23712
rect 21416 23672 21422 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 23474 23721 23480 23724
rect 22704 23684 23428 23712
rect 22704 23672 22710 23684
rect 17267 23616 17356 23644
rect 23400 23644 23428 23684
rect 23472 23675 23480 23721
rect 23474 23672 23480 23675
rect 23532 23672 23538 23724
rect 23676 23644 23704 23743
rect 23750 23672 23756 23724
rect 23808 23721 23814 23724
rect 23808 23715 23847 23721
rect 23835 23681 23847 23715
rect 23808 23675 23847 23681
rect 23808 23672 23814 23675
rect 23934 23672 23940 23724
rect 23992 23672 23998 23724
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 24780 23712 24808 23808
rect 24872 23780 24900 23811
rect 25194 23783 25252 23789
rect 25194 23780 25206 23783
rect 24872 23752 25206 23780
rect 25194 23749 25206 23752
rect 25240 23749 25252 23783
rect 25194 23743 25252 23749
rect 24719 23684 24808 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 23400 23616 23704 23644
rect 17267 23613 17279 23616
rect 17221 23607 17279 23613
rect 24394 23604 24400 23656
rect 24452 23644 24458 23656
rect 24949 23647 25007 23653
rect 24949 23644 24961 23647
rect 24452 23616 24961 23644
rect 24452 23604 24458 23616
rect 24949 23613 24961 23616
rect 24995 23613 25007 23647
rect 24949 23607 25007 23613
rect 16850 23536 16856 23588
rect 16908 23576 16914 23588
rect 17037 23579 17095 23585
rect 17037 23576 17049 23579
rect 16908 23548 17049 23576
rect 16908 23536 16914 23548
rect 17037 23545 17049 23548
rect 17083 23545 17095 23579
rect 17037 23539 17095 23545
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 19392 23548 21680 23576
rect 19392 23536 19398 23548
rect 21652 23520 21680 23548
rect 2455 23480 2774 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 3970 23468 3976 23520
rect 4028 23468 4034 23520
rect 4798 23468 4804 23520
rect 4856 23508 4862 23520
rect 5077 23511 5135 23517
rect 5077 23508 5089 23511
rect 4856 23480 5089 23508
rect 4856 23468 4862 23480
rect 5077 23477 5089 23480
rect 5123 23477 5135 23511
rect 5077 23471 5135 23477
rect 6546 23468 6552 23520
rect 6604 23468 6610 23520
rect 7282 23468 7288 23520
rect 7340 23468 7346 23520
rect 7561 23511 7619 23517
rect 7561 23477 7573 23511
rect 7607 23508 7619 23511
rect 7742 23508 7748 23520
rect 7607 23480 7748 23508
rect 7607 23477 7619 23480
rect 7561 23471 7619 23477
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 7834 23468 7840 23520
rect 7892 23508 7898 23520
rect 8662 23508 8668 23520
rect 7892 23480 8668 23508
rect 7892 23468 7898 23480
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9398 23508 9404 23520
rect 8996 23480 9404 23508
rect 8996 23468 9002 23480
rect 9398 23468 9404 23480
rect 9456 23508 9462 23520
rect 9585 23511 9643 23517
rect 9585 23508 9597 23511
rect 9456 23480 9597 23508
rect 9456 23468 9462 23480
rect 9585 23477 9597 23480
rect 9631 23477 9643 23511
rect 9585 23471 9643 23477
rect 10870 23468 10876 23520
rect 10928 23468 10934 23520
rect 12066 23468 12072 23520
rect 12124 23468 12130 23520
rect 14458 23468 14464 23520
rect 14516 23468 14522 23520
rect 16022 23468 16028 23520
rect 16080 23468 16086 23520
rect 18690 23468 18696 23520
rect 18748 23468 18754 23520
rect 18874 23468 18880 23520
rect 18932 23468 18938 23520
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 19978 23468 19984 23520
rect 20036 23468 20042 23520
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 21082 23508 21088 23520
rect 20855 23480 21088 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 21634 23468 21640 23520
rect 21692 23468 21698 23520
rect 22462 23468 22468 23520
rect 22520 23508 22526 23520
rect 23293 23511 23351 23517
rect 23293 23508 23305 23511
rect 22520 23480 23305 23508
rect 22520 23468 22526 23480
rect 23293 23477 23305 23480
rect 23339 23477 23351 23511
rect 23293 23471 23351 23477
rect 26326 23468 26332 23520
rect 26384 23468 26390 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 2958 23264 2964 23316
rect 3016 23304 3022 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 3016 23276 5089 23304
rect 3016 23264 3022 23276
rect 5077 23273 5089 23276
rect 5123 23273 5135 23307
rect 5077 23267 5135 23273
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 5813 23307 5871 23313
rect 5813 23304 5825 23307
rect 5684 23276 5825 23304
rect 5684 23264 5690 23276
rect 5813 23273 5825 23276
rect 5859 23273 5871 23307
rect 5813 23267 5871 23273
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 8113 23307 8171 23313
rect 8113 23304 8125 23307
rect 7248 23276 8125 23304
rect 7248 23264 7254 23276
rect 8113 23273 8125 23276
rect 8159 23273 8171 23307
rect 8113 23267 8171 23273
rect 8297 23307 8355 23313
rect 8297 23273 8309 23307
rect 8343 23304 8355 23307
rect 8478 23304 8484 23316
rect 8343 23276 8484 23304
rect 8343 23273 8355 23276
rect 8297 23267 8355 23273
rect 2130 23196 2136 23248
rect 2188 23236 2194 23248
rect 2590 23236 2596 23248
rect 2188 23208 2596 23236
rect 2188 23196 2194 23208
rect 2590 23196 2596 23208
rect 2648 23236 2654 23248
rect 6914 23236 6920 23248
rect 2648 23208 6920 23236
rect 2648 23196 2654 23208
rect 6914 23196 6920 23208
rect 6972 23236 6978 23248
rect 7377 23239 7435 23245
rect 7377 23236 7389 23239
rect 6972 23208 7389 23236
rect 6972 23196 6978 23208
rect 7377 23205 7389 23208
rect 7423 23205 7435 23239
rect 7377 23199 7435 23205
rect 1578 23128 1584 23180
rect 1636 23168 1642 23180
rect 5721 23171 5779 23177
rect 1636 23140 3280 23168
rect 1636 23128 1642 23140
rect 1854 23060 1860 23112
rect 1912 23100 1918 23112
rect 2317 23103 2375 23109
rect 2317 23100 2329 23103
rect 1912 23072 2329 23100
rect 1912 23060 1918 23072
rect 2317 23069 2329 23072
rect 2363 23100 2375 23103
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2363 23072 2881 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 2958 23060 2964 23112
rect 3016 23060 3022 23112
rect 3252 23109 3280 23140
rect 5721 23137 5733 23171
rect 5767 23137 5779 23171
rect 5721 23131 5779 23137
rect 5905 23171 5963 23177
rect 5905 23137 5917 23171
rect 5951 23168 5963 23171
rect 8128 23168 8156 23267
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 9401 23307 9459 23313
rect 9401 23273 9413 23307
rect 9447 23304 9459 23307
rect 9490 23304 9496 23316
rect 9447 23276 9496 23304
rect 9447 23273 9459 23276
rect 9401 23267 9459 23273
rect 9490 23264 9496 23276
rect 9548 23264 9554 23316
rect 9585 23307 9643 23313
rect 9585 23273 9597 23307
rect 9631 23304 9643 23307
rect 10226 23304 10232 23316
rect 9631 23276 10232 23304
rect 9631 23273 9643 23276
rect 9585 23267 9643 23273
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 10502 23264 10508 23316
rect 10560 23264 10566 23316
rect 11238 23264 11244 23316
rect 11296 23264 11302 23316
rect 13906 23264 13912 23316
rect 13964 23304 13970 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 13964 23276 14473 23304
rect 13964 23264 13970 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 15470 23264 15476 23316
rect 15528 23304 15534 23316
rect 15565 23307 15623 23313
rect 15565 23304 15577 23307
rect 15528 23276 15577 23304
rect 15528 23264 15534 23276
rect 15565 23273 15577 23276
rect 15611 23273 15623 23307
rect 15565 23267 15623 23273
rect 18782 23264 18788 23316
rect 18840 23264 18846 23316
rect 19334 23304 19340 23316
rect 18892 23276 19340 23304
rect 8386 23196 8392 23248
rect 8444 23196 8450 23248
rect 9950 23196 9956 23248
rect 10008 23236 10014 23248
rect 10045 23239 10103 23245
rect 10045 23236 10057 23239
rect 10008 23208 10057 23236
rect 10008 23196 10014 23208
rect 10045 23205 10057 23208
rect 10091 23205 10103 23239
rect 10045 23199 10103 23205
rect 10870 23196 10876 23248
rect 10928 23196 10934 23248
rect 14645 23239 14703 23245
rect 14645 23205 14657 23239
rect 14691 23236 14703 23239
rect 15657 23239 15715 23245
rect 15657 23236 15669 23239
rect 14691 23208 15669 23236
rect 14691 23205 14703 23208
rect 14645 23199 14703 23205
rect 15657 23205 15669 23208
rect 15703 23205 15715 23239
rect 15657 23199 15715 23205
rect 15933 23239 15991 23245
rect 15933 23205 15945 23239
rect 15979 23236 15991 23239
rect 18892 23236 18920 23276
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 19426 23264 19432 23316
rect 19484 23264 19490 23316
rect 19981 23307 20039 23313
rect 19981 23273 19993 23307
rect 20027 23304 20039 23307
rect 20622 23304 20628 23316
rect 20027 23276 20628 23304
rect 20027 23273 20039 23276
rect 19981 23267 20039 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 21266 23264 21272 23316
rect 21324 23304 21330 23316
rect 21453 23307 21511 23313
rect 21453 23304 21465 23307
rect 21324 23276 21465 23304
rect 21324 23264 21330 23276
rect 21453 23273 21465 23276
rect 21499 23273 21511 23307
rect 21453 23267 21511 23273
rect 23017 23307 23075 23313
rect 23017 23273 23029 23307
rect 23063 23304 23075 23307
rect 23934 23304 23940 23316
rect 23063 23276 23940 23304
rect 23063 23273 23075 23276
rect 23017 23267 23075 23273
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 15979 23208 18920 23236
rect 15979 23205 15991 23208
rect 15933 23199 15991 23205
rect 18966 23196 18972 23248
rect 19024 23236 19030 23248
rect 19245 23239 19303 23245
rect 19245 23236 19257 23239
rect 19024 23208 19257 23236
rect 19024 23196 19030 23208
rect 19245 23205 19257 23208
rect 19291 23205 19303 23239
rect 19245 23199 19303 23205
rect 20162 23196 20168 23248
rect 20220 23196 20226 23248
rect 22830 23196 22836 23248
rect 22888 23236 22894 23248
rect 23382 23236 23388 23248
rect 22888 23208 23388 23236
rect 22888 23196 22894 23208
rect 23382 23196 23388 23208
rect 23440 23196 23446 23248
rect 9030 23168 9036 23180
rect 5951 23140 7788 23168
rect 8128 23140 9036 23168
rect 5951 23137 5963 23140
rect 5905 23131 5963 23137
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23069 3295 23103
rect 3237 23063 3295 23069
rect 1946 22992 1952 23044
rect 2004 22992 2010 23044
rect 2593 23035 2651 23041
rect 2593 23001 2605 23035
rect 2639 23032 2651 23035
rect 2682 23032 2688 23044
rect 2639 23004 2688 23032
rect 2639 23001 2651 23004
rect 2593 22995 2651 23001
rect 2682 22992 2688 23004
rect 2740 23032 2746 23044
rect 2976 23032 3004 23060
rect 2740 23004 3004 23032
rect 2740 22992 2746 23004
rect 1964 22964 1992 22992
rect 2498 22964 2504 22976
rect 1964 22936 2504 22964
rect 2498 22924 2504 22936
rect 2556 22964 2562 22976
rect 3068 22964 3096 23063
rect 3252 23032 3280 23063
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 3789 23103 3847 23109
rect 3789 23100 3801 23103
rect 3476 23072 3801 23100
rect 3476 23060 3482 23072
rect 3789 23069 3801 23072
rect 3835 23069 3847 23103
rect 3789 23063 3847 23069
rect 4982 23060 4988 23112
rect 5040 23060 5046 23112
rect 5000 23032 5028 23060
rect 3252 23004 5028 23032
rect 5534 22964 5540 22976
rect 2556 22936 5540 22964
rect 2556 22924 2562 22936
rect 5534 22924 5540 22936
rect 5592 22924 5598 22976
rect 5736 22964 5764 23131
rect 7760 23112 7788 23140
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23100 6055 23103
rect 6638 23100 6644 23112
rect 6043 23072 6644 23100
rect 6043 23069 6055 23072
rect 5997 23063 6055 23069
rect 6638 23060 6644 23072
rect 6696 23060 6702 23112
rect 7742 23060 7748 23112
rect 7800 23060 7806 23112
rect 7834 23060 7840 23112
rect 7892 23060 7898 23112
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23094 8447 23103
rect 8588 23094 8616 23140
rect 9030 23128 9036 23140
rect 9088 23128 9094 23180
rect 9217 23171 9275 23177
rect 9217 23137 9229 23171
rect 9263 23168 9275 23171
rect 9858 23168 9864 23180
rect 9263 23140 9864 23168
rect 9263 23137 9275 23140
rect 9217 23131 9275 23137
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 10888 23168 10916 23196
rect 9968 23140 10916 23168
rect 9968 23109 9996 23140
rect 8435 23069 8616 23094
rect 8389 23066 8616 23069
rect 8665 23103 8723 23109
rect 8665 23069 8677 23103
rect 8711 23069 8723 23103
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8389 23063 8447 23066
rect 8665 23063 8723 23069
rect 9048 23072 9137 23100
rect 6086 22992 6092 23044
rect 6144 22992 6150 23044
rect 7852 23032 7880 23060
rect 7929 23035 7987 23041
rect 7929 23032 7941 23035
rect 7852 23004 7941 23032
rect 7929 23001 7941 23004
rect 7975 23001 7987 23035
rect 8680 23032 8708 23063
rect 7929 22995 7987 23001
rect 8404 23004 8708 23032
rect 6822 22964 6828 22976
rect 5736 22936 6828 22964
rect 6822 22924 6828 22936
rect 6880 22924 6886 22976
rect 7558 22924 7564 22976
rect 7616 22964 7622 22976
rect 8139 22967 8197 22973
rect 8139 22964 8151 22967
rect 7616 22936 8151 22964
rect 7616 22924 7622 22936
rect 8139 22933 8151 22936
rect 8185 22964 8197 22967
rect 8404 22964 8432 23004
rect 9048 22976 9076 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10042 23060 10048 23112
rect 10100 23060 10106 23112
rect 10134 23060 10140 23112
rect 10192 23060 10198 23112
rect 10318 23060 10324 23112
rect 10376 23060 10382 23112
rect 10612 23109 10640 23140
rect 10962 23128 10968 23180
rect 11020 23128 11026 23180
rect 16850 23168 16856 23180
rect 15120 23140 16856 23168
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23069 10471 23103
rect 10413 23063 10471 23069
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 10873 23103 10931 23109
rect 10873 23069 10885 23103
rect 10919 23100 10931 23103
rect 10980 23100 11008 23128
rect 10919 23072 11008 23100
rect 11057 23103 11115 23109
rect 10919 23069 10931 23072
rect 10873 23063 10931 23069
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 12529 23103 12587 23109
rect 11103 23072 11560 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 9674 22992 9680 23044
rect 9732 23032 9738 23044
rect 9769 23035 9827 23041
rect 9769 23032 9781 23035
rect 9732 23004 9781 23032
rect 9732 22992 9738 23004
rect 9769 23001 9781 23004
rect 9815 23032 9827 23035
rect 9815 23004 10180 23032
rect 9815 23001 9827 23004
rect 9769 22995 9827 23001
rect 8185 22936 8432 22964
rect 8573 22967 8631 22973
rect 8185 22933 8197 22936
rect 8139 22927 8197 22933
rect 8573 22933 8585 22967
rect 8619 22964 8631 22967
rect 8662 22964 8668 22976
rect 8619 22936 8668 22964
rect 8619 22933 8631 22936
rect 8573 22927 8631 22933
rect 8662 22924 8668 22936
rect 8720 22924 8726 22976
rect 9030 22924 9036 22976
rect 9088 22924 9094 22976
rect 10152 22964 10180 23004
rect 10428 22964 10456 23063
rect 11532 22976 11560 23072
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 14642 23100 14648 23112
rect 12575 23072 13032 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 13004 23044 13032 23072
rect 14292 23072 14648 23100
rect 12796 23035 12854 23041
rect 12796 23001 12808 23035
rect 12842 23032 12854 23035
rect 12894 23032 12900 23044
rect 12842 23004 12900 23032
rect 12842 23001 12854 23004
rect 12796 22995 12854 23001
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 12986 22992 12992 23044
rect 13044 22992 13050 23044
rect 14292 23041 14320 23072
rect 14642 23060 14648 23072
rect 14700 23060 14706 23112
rect 14277 23035 14335 23041
rect 14277 23032 14289 23035
rect 13096 23004 14289 23032
rect 10152 22936 10456 22964
rect 11514 22924 11520 22976
rect 11572 22924 11578 22976
rect 11606 22924 11612 22976
rect 11664 22964 11670 22976
rect 13096 22964 13124 23004
rect 14277 23001 14289 23004
rect 14323 23001 14335 23035
rect 15120 23032 15148 23140
rect 16850 23128 16856 23140
rect 16908 23168 16914 23180
rect 18325 23171 18383 23177
rect 18325 23168 18337 23171
rect 16908 23140 17264 23168
rect 16908 23128 16914 23140
rect 15197 23103 15255 23109
rect 15197 23069 15209 23103
rect 15243 23100 15255 23103
rect 15286 23100 15292 23112
rect 15243 23072 15292 23100
rect 15243 23069 15255 23072
rect 15197 23063 15255 23069
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 15378 23060 15384 23112
rect 15436 23060 15442 23112
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 16114 23060 16120 23112
rect 16172 23060 16178 23112
rect 16209 23103 16267 23109
rect 16209 23069 16221 23103
rect 16255 23100 16267 23103
rect 16255 23072 16344 23100
rect 16255 23069 16267 23072
rect 16209 23063 16267 23069
rect 14277 22995 14335 23001
rect 14384 23004 15148 23032
rect 11664 22936 13124 22964
rect 13909 22967 13967 22973
rect 11664 22924 11670 22936
rect 13909 22933 13921 22967
rect 13955 22964 13967 22967
rect 14384 22964 14412 23004
rect 13955 22936 14412 22964
rect 14487 22967 14545 22973
rect 13955 22933 13967 22936
rect 13909 22927 13967 22933
rect 14487 22933 14499 22967
rect 14533 22964 14545 22967
rect 15194 22964 15200 22976
rect 14533 22936 15200 22964
rect 14533 22933 14545 22936
rect 14487 22927 14545 22933
rect 15194 22924 15200 22936
rect 15252 22964 15258 22976
rect 16316 22964 16344 23072
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17092 23072 17141 23100
rect 17092 23060 17098 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 17236 23041 17264 23140
rect 17328 23140 18337 23168
rect 17328 23109 17356 23140
rect 18325 23137 18337 23140
rect 18371 23168 18383 23171
rect 22646 23168 22652 23180
rect 18371 23140 19564 23168
rect 18371 23137 18383 23140
rect 18325 23131 18383 23137
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 17460 23072 17509 23100
rect 17460 23060 17466 23072
rect 17497 23069 17509 23072
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 19334 23100 19340 23112
rect 18187 23072 19340 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 17221 23035 17279 23041
rect 17221 23001 17233 23035
rect 17267 23001 17279 23035
rect 18064 23032 18092 23063
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 19536 23100 19564 23140
rect 19711 23140 20208 23168
rect 19711 23100 19739 23140
rect 19536 23072 19739 23100
rect 20180 23100 20208 23140
rect 22112 23140 22652 23168
rect 22112 23100 22140 23140
rect 20180 23072 22140 23100
rect 22186 23060 22192 23112
rect 22244 23060 22250 23112
rect 22278 23060 22284 23112
rect 22336 23060 22342 23112
rect 22370 23060 22376 23112
rect 22428 23060 22434 23112
rect 22572 23109 22600 23140
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 22802 23140 23520 23168
rect 22802 23112 22830 23140
rect 23492 23112 23520 23140
rect 23584 23140 24532 23168
rect 22802 23109 22836 23112
rect 22557 23103 22615 23109
rect 22557 23069 22569 23103
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 22787 23103 22836 23109
rect 22787 23069 22799 23103
rect 22833 23069 22836 23103
rect 22787 23063 22836 23069
rect 22830 23060 22836 23063
rect 22888 23060 22894 23112
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23069 23259 23103
rect 23201 23063 23259 23069
rect 18064 23004 18184 23032
rect 17221 22995 17279 23001
rect 18156 22976 18184 23004
rect 18598 22992 18604 23044
rect 18656 22992 18662 23044
rect 19810 23041 19816 23044
rect 19567 23035 19625 23041
rect 19567 23032 19579 23035
rect 18708 23004 19579 23032
rect 15252 22936 16344 22964
rect 15252 22924 15258 22936
rect 16390 22924 16396 22976
rect 16448 22924 16454 22976
rect 16945 22967 17003 22973
rect 16945 22933 16957 22967
rect 16991 22964 17003 22967
rect 17402 22964 17408 22976
rect 16991 22936 17408 22964
rect 16991 22933 17003 22936
rect 16945 22927 17003 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 18138 22924 18144 22976
rect 18196 22924 18202 22976
rect 18625 22964 18653 22992
rect 18708 22964 18736 23004
rect 19567 23001 19579 23004
rect 19613 23001 19625 23035
rect 19567 22995 19625 23001
rect 19797 23035 19816 23041
rect 19797 23001 19809 23035
rect 19797 22995 19816 23001
rect 19810 22992 19816 22995
rect 19868 22992 19874 23044
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 21085 23035 21143 23041
rect 21085 23032 21097 23035
rect 20588 23004 21097 23032
rect 20588 22992 20594 23004
rect 21085 23001 21097 23004
rect 21131 23001 21143 23035
rect 21085 22995 21143 23001
rect 21266 22992 21272 23044
rect 21324 22992 21330 23044
rect 22204 23032 22232 23060
rect 22649 23035 22707 23041
rect 22649 23032 22661 23035
rect 22204 23004 22661 23032
rect 22649 23001 22661 23004
rect 22695 23001 22707 23035
rect 22649 22995 22707 23001
rect 23014 22992 23020 23044
rect 23072 23032 23078 23044
rect 23216 23032 23244 23063
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 23474 23060 23480 23112
rect 23532 23060 23538 23112
rect 23584 23109 23612 23140
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 24394 23060 24400 23112
rect 24452 23060 24458 23112
rect 24504 23100 24532 23140
rect 24946 23100 24952 23112
rect 24504 23072 24952 23100
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 23072 23004 23244 23032
rect 23293 23035 23351 23041
rect 23072 22992 23078 23004
rect 23293 23001 23305 23035
rect 23339 23001 23351 23035
rect 23293 22995 23351 23001
rect 18625 22936 18736 22964
rect 18782 22924 18788 22976
rect 18840 22973 18846 22976
rect 18840 22967 18859 22973
rect 18847 22933 18859 22967
rect 18840 22927 18859 22933
rect 18840 22924 18846 22927
rect 18966 22924 18972 22976
rect 19024 22924 19030 22976
rect 19426 22973 19432 22976
rect 19413 22967 19432 22973
rect 19413 22933 19425 22967
rect 19484 22964 19490 22976
rect 20007 22967 20065 22973
rect 20007 22964 20019 22967
rect 19484 22936 20019 22964
rect 19413 22927 19432 22933
rect 19426 22924 19432 22927
rect 19484 22924 19490 22936
rect 20007 22933 20019 22936
rect 20053 22964 20065 22967
rect 20714 22964 20720 22976
rect 20053 22936 20720 22964
rect 20053 22933 20065 22936
rect 20007 22927 20065 22933
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 22925 22967 22983 22973
rect 22925 22964 22937 22967
rect 22244 22936 22937 22964
rect 22244 22924 22250 22936
rect 22925 22933 22937 22936
rect 22971 22933 22983 22967
rect 23308 22964 23336 22995
rect 23934 22992 23940 23044
rect 23992 23032 23998 23044
rect 24642 23035 24700 23041
rect 24642 23032 24654 23035
rect 23992 23004 24654 23032
rect 23992 22992 23998 23004
rect 24642 23001 24654 23004
rect 24688 23001 24700 23035
rect 24642 22995 24700 23001
rect 25774 22964 25780 22976
rect 23308 22936 25780 22964
rect 22925 22927 22983 22933
rect 25774 22924 25780 22936
rect 25832 22924 25838 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2314 22760 2320 22772
rect 1820 22732 2320 22760
rect 1820 22720 1826 22732
rect 2314 22720 2320 22732
rect 2372 22760 2378 22772
rect 2501 22763 2559 22769
rect 2501 22760 2513 22763
rect 2372 22732 2513 22760
rect 2372 22720 2378 22732
rect 2501 22729 2513 22732
rect 2547 22729 2559 22763
rect 2501 22723 2559 22729
rect 2590 22720 2596 22772
rect 2648 22720 2654 22772
rect 2774 22760 2780 22772
rect 2746 22720 2780 22760
rect 2832 22720 2838 22772
rect 3694 22720 3700 22772
rect 3752 22760 3758 22772
rect 3881 22763 3939 22769
rect 3881 22760 3893 22763
rect 3752 22732 3893 22760
rect 3752 22720 3758 22732
rect 3881 22729 3893 22732
rect 3927 22729 3939 22763
rect 3881 22723 3939 22729
rect 4246 22720 4252 22772
rect 4304 22760 4310 22772
rect 5445 22763 5503 22769
rect 5445 22760 5457 22763
rect 4304 22732 5457 22760
rect 4304 22720 4310 22732
rect 5445 22729 5457 22732
rect 5491 22729 5503 22763
rect 5445 22723 5503 22729
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5994 22760 6000 22772
rect 5592 22732 6000 22760
rect 5592 22720 5598 22732
rect 5994 22720 6000 22732
rect 6052 22760 6058 22772
rect 6362 22760 6368 22772
rect 6052 22732 6368 22760
rect 6052 22720 6058 22732
rect 6362 22720 6368 22732
rect 6420 22720 6426 22772
rect 7466 22760 7472 22772
rect 6840 22732 7472 22760
rect 1949 22695 2007 22701
rect 1949 22661 1961 22695
rect 1995 22661 2007 22695
rect 1949 22655 2007 22661
rect 2225 22695 2283 22701
rect 2225 22661 2237 22695
rect 2271 22692 2283 22695
rect 2746 22692 2774 22720
rect 2271 22664 2774 22692
rect 2271 22661 2283 22664
rect 2225 22655 2283 22661
rect 1578 22584 1584 22636
rect 1636 22584 1642 22636
rect 1964 22488 1992 22655
rect 2866 22652 2872 22704
rect 2924 22692 2930 22704
rect 6840 22701 6868 22732
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 9033 22763 9091 22769
rect 8444 22732 8892 22760
rect 8444 22720 8450 22732
rect 6825 22695 6883 22701
rect 2924 22664 6040 22692
rect 2924 22652 2930 22664
rect 2409 22627 2467 22633
rect 2409 22624 2421 22627
rect 2240 22596 2421 22624
rect 2240 22568 2268 22596
rect 2409 22593 2421 22596
rect 2455 22593 2467 22627
rect 2409 22587 2467 22593
rect 2777 22627 2835 22633
rect 2777 22593 2789 22627
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 2222 22516 2228 22568
rect 2280 22516 2286 22568
rect 2792 22556 2820 22587
rect 3142 22584 3148 22636
rect 3200 22584 3206 22636
rect 3234 22584 3240 22636
rect 3292 22584 3298 22636
rect 3326 22584 3332 22636
rect 3384 22584 3390 22636
rect 3513 22627 3571 22633
rect 3513 22593 3525 22627
rect 3559 22624 3571 22627
rect 3878 22624 3884 22636
rect 3559 22596 3884 22624
rect 3559 22593 3571 22596
rect 3513 22587 3571 22593
rect 2869 22559 2927 22565
rect 2869 22556 2881 22559
rect 2792 22528 2881 22556
rect 2869 22525 2881 22528
rect 2915 22525 2927 22559
rect 2869 22519 2927 22525
rect 3050 22516 3056 22568
rect 3108 22556 3114 22568
rect 3528 22556 3556 22587
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 5350 22584 5356 22636
rect 5408 22584 5414 22636
rect 5736 22633 5764 22664
rect 6012 22636 6040 22664
rect 6825 22661 6837 22695
rect 6871 22661 6883 22695
rect 6825 22655 6883 22661
rect 6917 22695 6975 22701
rect 6917 22661 6929 22695
rect 6963 22692 6975 22695
rect 7653 22695 7711 22701
rect 7653 22692 7665 22695
rect 6963 22664 7665 22692
rect 6963 22661 6975 22664
rect 6917 22655 6975 22661
rect 7653 22661 7665 22664
rect 7699 22661 7711 22695
rect 7653 22655 7711 22661
rect 7742 22652 7748 22704
rect 7800 22692 7806 22704
rect 7800 22664 8708 22692
rect 7800 22652 7806 22664
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22593 5963 22627
rect 5905 22587 5963 22593
rect 3108 22528 3556 22556
rect 4816 22556 4844 22584
rect 5828 22556 5856 22587
rect 4816 22528 5856 22556
rect 3108 22516 3114 22528
rect 2958 22488 2964 22500
rect 1964 22460 2964 22488
rect 2958 22448 2964 22460
rect 3016 22488 3022 22500
rect 4338 22488 4344 22500
rect 3016 22460 4344 22488
rect 3016 22448 3022 22460
rect 4338 22448 4344 22460
rect 4396 22448 4402 22500
rect 1946 22380 1952 22432
rect 2004 22380 2010 22432
rect 2130 22380 2136 22432
rect 2188 22380 2194 22432
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 4890 22420 4896 22432
rect 4304 22392 4896 22420
rect 4304 22380 4310 22392
rect 4890 22380 4896 22392
rect 4948 22420 4954 22432
rect 5920 22420 5948 22587
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6089 22627 6147 22633
rect 6089 22593 6101 22627
rect 6135 22624 6147 22627
rect 6728 22627 6786 22633
rect 6135 22596 6592 22624
rect 6135 22593 6147 22596
rect 6089 22587 6147 22593
rect 6564 22497 6592 22596
rect 6728 22593 6740 22627
rect 6774 22593 6786 22627
rect 6728 22587 6786 22593
rect 6549 22491 6607 22497
rect 6549 22457 6561 22491
rect 6595 22457 6607 22491
rect 6549 22451 6607 22457
rect 4948 22392 5948 22420
rect 4948 22380 4954 22392
rect 6454 22380 6460 22432
rect 6512 22420 6518 22432
rect 6743 22420 6771 22587
rect 7006 22584 7012 22636
rect 7064 22633 7070 22636
rect 7064 22627 7103 22633
rect 7091 22593 7103 22627
rect 7064 22587 7103 22593
rect 7064 22584 7070 22587
rect 7190 22584 7196 22636
rect 7248 22584 7254 22636
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22593 7895 22627
rect 7837 22587 7895 22593
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22624 7987 22627
rect 8018 22624 8024 22636
rect 7975 22596 8024 22624
rect 7975 22593 7987 22596
rect 7929 22587 7987 22593
rect 7852 22488 7880 22587
rect 8018 22584 8024 22596
rect 8076 22584 8082 22636
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8128 22556 8156 22587
rect 8202 22584 8208 22636
rect 8260 22584 8266 22636
rect 8478 22584 8484 22636
rect 8536 22584 8542 22636
rect 8680 22633 8708 22664
rect 8665 22627 8723 22633
rect 8665 22593 8677 22627
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 8386 22556 8392 22568
rect 8128 22528 8392 22556
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 8772 22556 8800 22587
rect 8680 22528 8800 22556
rect 8680 22500 8708 22528
rect 8573 22491 8631 22497
rect 8573 22488 8585 22491
rect 7852 22460 8585 22488
rect 8573 22457 8585 22460
rect 8619 22457 8631 22491
rect 8573 22451 8631 22457
rect 6512 22392 6771 22420
rect 6512 22380 6518 22392
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 8297 22423 8355 22429
rect 8297 22420 8309 22423
rect 7524 22392 8309 22420
rect 7524 22380 7530 22392
rect 8297 22389 8309 22392
rect 8343 22389 8355 22423
rect 8588 22420 8616 22451
rect 8662 22448 8668 22500
rect 8720 22448 8726 22500
rect 8864 22420 8892 22732
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 9306 22760 9312 22772
rect 9079 22732 9312 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 11514 22720 11520 22772
rect 11572 22720 11578 22772
rect 11698 22720 11704 22772
rect 11756 22760 11762 22772
rect 12437 22763 12495 22769
rect 12437 22760 12449 22763
rect 11756 22732 12449 22760
rect 11756 22720 11762 22732
rect 12437 22729 12449 22732
rect 12483 22729 12495 22763
rect 12437 22723 12495 22729
rect 12894 22720 12900 22772
rect 12952 22720 12958 22772
rect 15381 22763 15439 22769
rect 15381 22729 15393 22763
rect 15427 22760 15439 22763
rect 15470 22760 15476 22772
rect 15427 22732 15476 22760
rect 15427 22729 15439 22732
rect 15381 22723 15439 22729
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 16758 22720 16764 22772
rect 16816 22760 16822 22772
rect 17218 22760 17224 22772
rect 16816 22732 17224 22760
rect 16816 22720 16822 22732
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 19610 22760 19616 22772
rect 19428 22732 19616 22760
rect 15013 22695 15071 22701
rect 11900 22664 12271 22692
rect 11900 22636 11928 22664
rect 9125 22627 9183 22633
rect 9125 22593 9137 22627
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9140 22556 9168 22587
rect 11882 22584 11888 22636
rect 11940 22584 11946 22636
rect 11974 22584 11980 22636
rect 12032 22584 12038 22636
rect 12243 22633 12271 22664
rect 15013 22661 15025 22695
rect 15059 22661 15071 22695
rect 15013 22655 15071 22661
rect 15229 22695 15287 22701
rect 15229 22661 15241 22695
rect 15275 22692 15287 22695
rect 15746 22692 15752 22704
rect 15275 22664 15752 22692
rect 15275 22661 15287 22664
rect 15229 22655 15287 22661
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12228 22627 12286 22633
rect 12228 22593 12240 22627
rect 12274 22593 12286 22627
rect 12228 22587 12286 22593
rect 9088 22528 9168 22556
rect 9088 22516 9094 22528
rect 10870 22516 10876 22568
rect 10928 22556 10934 22568
rect 11238 22556 11244 22568
rect 10928 22528 11244 22556
rect 10928 22516 10934 22528
rect 11238 22516 11244 22528
rect 11296 22556 11302 22568
rect 11609 22559 11667 22565
rect 11609 22556 11621 22559
rect 11296 22528 11621 22556
rect 11296 22516 11302 22528
rect 11609 22525 11621 22528
rect 11655 22525 11667 22559
rect 11609 22519 11667 22525
rect 11698 22516 11704 22568
rect 11756 22516 11762 22568
rect 11790 22516 11796 22568
rect 11848 22556 11854 22568
rect 12084 22556 12112 22587
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 12710 22584 12716 22636
rect 12768 22584 12774 22636
rect 13354 22584 13360 22636
rect 13412 22624 13418 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 13412 22596 13461 22624
rect 13412 22584 13418 22596
rect 13449 22593 13461 22596
rect 13495 22593 13507 22627
rect 15028 22624 15056 22655
rect 15746 22652 15752 22664
rect 15804 22652 15810 22704
rect 16132 22664 18368 22692
rect 15470 22624 15476 22636
rect 15028 22596 15476 22624
rect 13449 22587 13507 22593
rect 15470 22584 15476 22596
rect 15528 22584 15534 22636
rect 16132 22624 16160 22664
rect 16040 22596 16160 22624
rect 16945 22627 17003 22633
rect 11848 22528 12112 22556
rect 11848 22516 11854 22528
rect 15378 22516 15384 22568
rect 15436 22556 15442 22568
rect 15654 22556 15660 22568
rect 15436 22528 15660 22556
rect 15436 22516 15442 22528
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 9122 22448 9128 22500
rect 9180 22488 9186 22500
rect 9180 22460 12388 22488
rect 9180 22448 9186 22460
rect 8588 22392 8892 22420
rect 11885 22423 11943 22429
rect 8297 22383 8355 22389
rect 11885 22389 11897 22423
rect 11931 22420 11943 22423
rect 12066 22420 12072 22432
rect 11931 22392 12072 22420
rect 11931 22389 11943 22392
rect 11885 22383 11943 22389
rect 12066 22380 12072 22392
rect 12124 22380 12130 22432
rect 12161 22423 12219 22429
rect 12161 22389 12173 22423
rect 12207 22420 12219 22423
rect 12250 22420 12256 22432
rect 12207 22392 12256 22420
rect 12207 22389 12219 22392
rect 12161 22383 12219 22389
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 12360 22420 12388 22460
rect 13170 22448 13176 22500
rect 13228 22488 13234 22500
rect 16040 22488 16068 22596
rect 16945 22593 16957 22627
rect 16991 22624 17003 22627
rect 17770 22624 17776 22636
rect 16991 22596 17776 22624
rect 16991 22593 17003 22596
rect 16945 22587 17003 22593
rect 17770 22584 17776 22596
rect 17828 22624 17834 22636
rect 17828 22596 18276 22624
rect 17828 22584 17834 22596
rect 16114 22516 16120 22568
rect 16172 22556 16178 22568
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16172 22528 16773 22556
rect 16172 22516 16178 22528
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 13228 22460 16068 22488
rect 16776 22488 16804 22519
rect 18138 22516 18144 22568
rect 18196 22516 18202 22568
rect 18156 22488 18184 22516
rect 16776 22460 18184 22488
rect 18248 22488 18276 22596
rect 18340 22556 18368 22664
rect 18966 22652 18972 22704
rect 19024 22652 19030 22704
rect 19428 22692 19456 22732
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 19705 22763 19763 22769
rect 19705 22729 19717 22763
rect 19751 22760 19763 22763
rect 19751 22732 20085 22760
rect 19751 22729 19763 22732
rect 19705 22723 19763 22729
rect 20057 22701 20085 22732
rect 23934 22720 23940 22772
rect 23992 22720 23998 22772
rect 25774 22720 25780 22772
rect 25832 22720 25838 22772
rect 19352 22664 19456 22692
rect 20042 22695 20100 22701
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18748 22596 18889 22624
rect 18748 22584 18754 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18984 22624 19012 22652
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 18984 22596 19073 22624
rect 18877 22587 18935 22593
rect 19061 22593 19073 22596
rect 19107 22593 19119 22627
rect 19061 22587 19119 22593
rect 19150 22584 19156 22636
rect 19208 22584 19214 22636
rect 19352 22633 19380 22664
rect 20042 22661 20054 22695
rect 20088 22661 20100 22695
rect 20042 22655 20100 22661
rect 20714 22652 20720 22704
rect 20772 22692 20778 22704
rect 22278 22692 22284 22704
rect 20772 22664 22284 22692
rect 20772 22652 20778 22664
rect 22278 22652 22284 22664
rect 22336 22652 22342 22704
rect 24486 22692 24492 22704
rect 23216 22664 24492 22692
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19518 22584 19524 22636
rect 19576 22584 19582 22636
rect 23216 22633 23244 22664
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 25130 22652 25136 22704
rect 25188 22692 25194 22704
rect 25225 22695 25283 22701
rect 25225 22692 25237 22695
rect 25188 22664 25237 22692
rect 25188 22652 25194 22664
rect 25225 22661 25237 22664
rect 25271 22661 25283 22695
rect 25225 22655 25283 22661
rect 23201 22627 23259 22633
rect 23201 22624 23213 22627
rect 19628 22596 23213 22624
rect 18340 22528 18828 22556
rect 18800 22488 18828 22528
rect 18966 22516 18972 22568
rect 19024 22516 19030 22568
rect 19628 22556 19656 22596
rect 23201 22593 23213 22596
rect 23247 22593 23259 22627
rect 23753 22627 23811 22633
rect 23753 22624 23765 22627
rect 23201 22587 23259 22593
rect 23676 22596 23765 22624
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19352 22528 19656 22556
rect 19711 22528 19809 22556
rect 19352 22488 19380 22528
rect 18248 22460 18736 22488
rect 18800 22460 19380 22488
rect 13228 22448 13234 22460
rect 13078 22420 13084 22432
rect 12360 22392 13084 22420
rect 13078 22380 13084 22392
rect 13136 22420 13142 22432
rect 13633 22423 13691 22429
rect 13633 22420 13645 22423
rect 13136 22392 13645 22420
rect 13136 22380 13142 22392
rect 13633 22389 13645 22392
rect 13679 22389 13691 22423
rect 13633 22383 13691 22389
rect 14734 22380 14740 22432
rect 14792 22420 14798 22432
rect 15197 22423 15255 22429
rect 15197 22420 15209 22423
rect 14792 22392 15209 22420
rect 14792 22380 14798 22392
rect 15197 22389 15209 22392
rect 15243 22389 15255 22423
rect 15197 22383 15255 22389
rect 17034 22380 17040 22432
rect 17092 22420 17098 22432
rect 17129 22423 17187 22429
rect 17129 22420 17141 22423
rect 17092 22392 17141 22420
rect 17092 22380 17098 22392
rect 17129 22389 17141 22392
rect 17175 22389 17187 22423
rect 17129 22383 17187 22389
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18601 22423 18659 22429
rect 18601 22420 18613 22423
rect 18104 22392 18613 22420
rect 18104 22380 18110 22392
rect 18601 22389 18613 22392
rect 18647 22389 18659 22423
rect 18708 22420 18736 22460
rect 19426 22448 19432 22500
rect 19484 22488 19490 22500
rect 19711 22488 19739 22528
rect 19797 22525 19809 22528
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 22738 22516 22744 22568
rect 22796 22556 22802 22568
rect 23676 22565 23704 22596
rect 23753 22593 23765 22596
rect 23799 22593 23811 22627
rect 25792 22624 25820 22720
rect 23753 22587 23811 22593
rect 24964 22596 25820 22624
rect 23661 22559 23719 22565
rect 22796 22528 23520 22556
rect 22796 22516 22802 22528
rect 23492 22497 23520 22528
rect 23661 22525 23673 22559
rect 23707 22525 23719 22559
rect 23661 22519 23719 22525
rect 19484 22460 19739 22488
rect 23477 22491 23535 22497
rect 19484 22448 19490 22460
rect 23477 22457 23489 22491
rect 23523 22457 23535 22491
rect 23477 22451 23535 22457
rect 24857 22491 24915 22497
rect 24857 22457 24869 22491
rect 24903 22488 24915 22491
rect 24964 22488 24992 22596
rect 24903 22460 24992 22488
rect 25593 22491 25651 22497
rect 24903 22457 24915 22460
rect 24857 22451 24915 22457
rect 25593 22457 25605 22491
rect 25639 22488 25651 22491
rect 26326 22488 26332 22500
rect 25639 22460 26332 22488
rect 25639 22457 25651 22460
rect 25593 22451 25651 22457
rect 26326 22448 26332 22460
rect 26384 22448 26390 22500
rect 18782 22420 18788 22432
rect 18708 22392 18788 22420
rect 18601 22383 18659 22389
rect 18782 22380 18788 22392
rect 18840 22420 18846 22432
rect 19978 22420 19984 22432
rect 18840 22392 19984 22420
rect 18840 22380 18846 22392
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 20438 22380 20444 22432
rect 20496 22420 20502 22432
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20496 22392 21189 22420
rect 20496 22380 20502 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 21177 22383 21235 22389
rect 24946 22380 24952 22432
rect 25004 22380 25010 22432
rect 25682 22380 25688 22432
rect 25740 22380 25746 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 1670 22176 1676 22228
rect 1728 22216 1734 22228
rect 1946 22216 1952 22228
rect 1728 22188 1952 22216
rect 1728 22176 1734 22188
rect 1946 22176 1952 22188
rect 2004 22176 2010 22228
rect 3970 22176 3976 22228
rect 4028 22176 4034 22228
rect 5718 22216 5724 22228
rect 4080 22188 5724 22216
rect 2314 22148 2320 22160
rect 1596 22120 2320 22148
rect 1596 22021 1624 22120
rect 2314 22108 2320 22120
rect 2372 22148 2378 22160
rect 2685 22151 2743 22157
rect 2685 22148 2697 22151
rect 2372 22120 2697 22148
rect 2372 22108 2378 22120
rect 2685 22117 2697 22120
rect 2731 22117 2743 22151
rect 2685 22111 2743 22117
rect 3786 22108 3792 22160
rect 3844 22108 3850 22160
rect 2774 22080 2780 22092
rect 1780 22052 2780 22080
rect 1780 22021 1808 22052
rect 2774 22040 2780 22052
rect 2832 22040 2838 22092
rect 3510 22040 3516 22092
rect 3568 22080 3574 22092
rect 3804 22080 3832 22108
rect 3988 22080 4016 22176
rect 3568 22052 3832 22080
rect 3896 22052 4016 22080
rect 3568 22040 3574 22052
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 21981 1639 22015
rect 1581 21975 1639 21981
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 1854 21972 1860 22024
rect 1912 21972 1918 22024
rect 2130 21972 2136 22024
rect 2188 22012 2194 22024
rect 3896 22021 3924 22052
rect 2501 22015 2559 22021
rect 2501 22012 2513 22015
rect 2188 21984 2513 22012
rect 2188 21972 2194 21984
rect 2501 21981 2513 21984
rect 2547 21981 2559 22015
rect 2501 21975 2559 21981
rect 3881 22015 3939 22021
rect 3881 21981 3893 22015
rect 3927 21981 3939 22015
rect 3881 21975 3939 21981
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 22012 4031 22015
rect 4080 22012 4108 22188
rect 5718 22176 5724 22188
rect 5776 22176 5782 22228
rect 6638 22216 6644 22228
rect 5828 22188 6644 22216
rect 4157 22151 4215 22157
rect 4157 22117 4169 22151
rect 4203 22117 4215 22151
rect 4157 22111 4215 22117
rect 4172 22080 4200 22111
rect 4525 22083 4583 22089
rect 4172 22052 4476 22080
rect 4019 21984 4108 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 1397 21947 1455 21953
rect 1397 21913 1409 21947
rect 1443 21944 1455 21947
rect 2041 21947 2099 21953
rect 2041 21944 2053 21947
rect 1443 21916 2053 21944
rect 1443 21913 1455 21916
rect 1397 21907 1455 21913
rect 2041 21913 2053 21916
rect 2087 21913 2099 21947
rect 2041 21907 2099 21913
rect 3418 21904 3424 21956
rect 3476 21944 3482 21956
rect 3988 21944 4016 21975
rect 4246 21972 4252 22024
rect 4304 21972 4310 22024
rect 4448 22021 4476 22052
rect 4525 22049 4537 22083
rect 4571 22080 4583 22083
rect 5629 22083 5687 22089
rect 5629 22080 5641 22083
rect 4571 22052 5641 22080
rect 4571 22049 4583 22052
rect 4525 22043 4583 22049
rect 5629 22049 5641 22052
rect 5675 22049 5687 22083
rect 5828 22080 5856 22188
rect 6638 22176 6644 22188
rect 6696 22176 6702 22228
rect 7742 22176 7748 22228
rect 7800 22216 7806 22228
rect 8294 22216 8300 22228
rect 7800 22188 8300 22216
rect 7800 22176 7806 22188
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 10781 22219 10839 22225
rect 10781 22185 10793 22219
rect 10827 22216 10839 22219
rect 10962 22216 10968 22228
rect 10827 22188 10968 22216
rect 10827 22185 10839 22188
rect 10781 22179 10839 22185
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 11517 22219 11575 22225
rect 11517 22185 11529 22219
rect 11563 22216 11575 22219
rect 11698 22216 11704 22228
rect 11563 22188 11704 22216
rect 11563 22185 11575 22188
rect 11517 22179 11575 22185
rect 6362 22108 6368 22160
rect 6420 22148 6426 22160
rect 6420 22120 6776 22148
rect 6420 22108 6426 22120
rect 5629 22043 5687 22049
rect 5736 22052 5856 22080
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 21981 4491 22015
rect 4433 21975 4491 21981
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 22012 4675 22015
rect 4706 22012 4712 22024
rect 4663 21984 4712 22012
rect 4663 21981 4675 21984
rect 4617 21975 4675 21981
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 4798 21972 4804 22024
rect 4856 21972 4862 22024
rect 5261 22015 5319 22021
rect 5261 21981 5273 22015
rect 5307 21981 5319 22015
rect 5261 21975 5319 21981
rect 3476 21916 4016 21944
rect 4157 21947 4215 21953
rect 3476 21904 3482 21916
rect 4157 21913 4169 21947
rect 4203 21944 4215 21947
rect 5077 21947 5135 21953
rect 5077 21944 5089 21947
rect 4203 21916 5089 21944
rect 4203 21913 4215 21916
rect 4157 21907 4215 21913
rect 5077 21913 5089 21916
rect 5123 21913 5135 21947
rect 5276 21944 5304 21975
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 5736 22012 5764 22052
rect 6178 22040 6184 22092
rect 6236 22040 6242 22092
rect 6748 22080 6776 22120
rect 6822 22108 6828 22160
rect 6880 22148 6886 22160
rect 8018 22148 8024 22160
rect 6880 22120 8024 22148
rect 6880 22108 6886 22120
rect 8018 22108 8024 22120
rect 8076 22148 8082 22160
rect 8662 22148 8668 22160
rect 8076 22120 8668 22148
rect 8076 22108 8082 22120
rect 8662 22108 8668 22120
rect 8720 22108 8726 22160
rect 11532 22148 11560 22179
rect 11698 22176 11704 22188
rect 11756 22176 11762 22228
rect 11974 22176 11980 22228
rect 12032 22216 12038 22228
rect 12069 22219 12127 22225
rect 12069 22216 12081 22219
rect 12032 22188 12081 22216
rect 12032 22176 12038 22188
rect 12069 22185 12081 22188
rect 12115 22185 12127 22219
rect 12069 22179 12127 22185
rect 12250 22176 12256 22228
rect 12308 22176 12314 22228
rect 15286 22176 15292 22228
rect 15344 22216 15350 22228
rect 17865 22219 17923 22225
rect 15344 22188 17080 22216
rect 15344 22176 15350 22188
rect 9646 22120 11284 22148
rect 6564 22052 6776 22080
rect 5592 21984 5764 22012
rect 5592 21972 5598 21984
rect 5810 21972 5816 22024
rect 5868 21972 5874 22024
rect 5902 21972 5908 22024
rect 5960 22012 5966 22024
rect 5997 22015 6055 22021
rect 5997 22012 6009 22015
rect 5960 21984 6009 22012
rect 5960 21972 5966 21984
rect 5997 21981 6009 21984
rect 6043 21981 6055 22015
rect 5997 21975 6055 21981
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 6104 21944 6132 21975
rect 6362 21972 6368 22024
rect 6420 21972 6426 22024
rect 6564 22021 6592 22052
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9646 22080 9674 22120
rect 9364 22052 9674 22080
rect 11256 22080 11284 22120
rect 11440 22120 11560 22148
rect 11440 22089 11468 22120
rect 11606 22108 11612 22160
rect 11664 22148 11670 22160
rect 12268 22148 12296 22176
rect 11664 22120 12296 22148
rect 17052 22148 17080 22188
rect 17865 22185 17877 22219
rect 17911 22216 17923 22219
rect 19334 22216 19340 22228
rect 17911 22188 19340 22216
rect 17911 22185 17923 22188
rect 17865 22179 17923 22185
rect 19334 22176 19340 22188
rect 19392 22176 19398 22228
rect 19610 22176 19616 22228
rect 19668 22176 19674 22228
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20806 22216 20812 22228
rect 20036 22188 20812 22216
rect 20036 22176 20042 22188
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 21376 22188 22600 22216
rect 18690 22148 18696 22160
rect 17052 22120 18696 22148
rect 11664 22108 11670 22120
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 19150 22108 19156 22160
rect 19208 22148 19214 22160
rect 20438 22148 20444 22160
rect 19208 22120 20444 22148
rect 19208 22108 19214 22120
rect 11425 22083 11483 22089
rect 11256 22052 11376 22080
rect 9364 22040 9370 22052
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 8202 22012 8208 22024
rect 6696 21984 8208 22012
rect 6696 21972 6702 21984
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 10505 22015 10563 22021
rect 10505 22012 10517 22015
rect 9968 21984 10517 22012
rect 9968 21956 9996 21984
rect 10505 21981 10517 21984
rect 10551 21981 10563 22015
rect 10870 22012 10876 22024
rect 10505 21975 10563 21981
rect 10704 21984 10876 22012
rect 6178 21944 6184 21956
rect 5276 21916 6184 21944
rect 5077 21907 5135 21913
rect 6178 21904 6184 21916
rect 6236 21944 6242 21956
rect 6454 21944 6460 21956
rect 6236 21916 6460 21944
rect 6236 21904 6242 21916
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 7006 21904 7012 21956
rect 7064 21904 7070 21956
rect 9950 21904 9956 21956
rect 10008 21904 10014 21956
rect 10321 21947 10379 21953
rect 10321 21913 10333 21947
rect 10367 21944 10379 21947
rect 10410 21944 10416 21956
rect 10367 21916 10416 21944
rect 10367 21913 10379 21916
rect 10321 21907 10379 21913
rect 2130 21836 2136 21888
rect 2188 21836 2194 21888
rect 4982 21836 4988 21888
rect 5040 21836 5046 21888
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 5408 21848 5457 21876
rect 5408 21836 5414 21848
rect 5445 21845 5457 21848
rect 5491 21845 5503 21879
rect 5445 21839 5503 21845
rect 5994 21836 6000 21888
rect 6052 21876 6058 21888
rect 6822 21876 6828 21888
rect 6052 21848 6828 21876
rect 6052 21836 6058 21848
rect 6822 21836 6828 21848
rect 6880 21836 6886 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 10336 21876 10364 21907
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 10704 21953 10732 21984
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 10962 21972 10968 22024
rect 11020 21972 11026 22024
rect 11054 21972 11060 22024
rect 11112 21972 11118 22024
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 22012 11207 22015
rect 11256 22012 11284 22052
rect 11195 21984 11284 22012
rect 11348 22012 11376 22052
rect 11425 22049 11437 22083
rect 11471 22049 11483 22083
rect 11425 22043 11483 22049
rect 16022 22040 16028 22092
rect 16080 22040 16086 22092
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22049 16175 22083
rect 20254 22080 20260 22092
rect 16117 22043 16175 22049
rect 17880 22052 19380 22080
rect 11348 21984 11468 22012
rect 11195 21981 11207 21984
rect 11149 21975 11207 21981
rect 10689 21947 10747 21953
rect 10689 21913 10701 21947
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 11238 21904 11244 21956
rect 11296 21953 11302 21956
rect 11296 21947 11325 21953
rect 11313 21913 11325 21947
rect 11440 21944 11468 21984
rect 11698 21972 11704 22024
rect 11756 21972 11762 22024
rect 11790 21972 11796 22024
rect 11848 22012 11854 22024
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11848 21984 11989 22012
rect 11848 21972 11854 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12802 21972 12808 22024
rect 12860 22012 12866 22024
rect 13354 22012 13360 22024
rect 12860 21984 13360 22012
rect 12860 21972 12866 21984
rect 13354 21972 13360 21984
rect 13412 22012 13418 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13412 21984 13461 22012
rect 13412 21972 13418 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 14829 22015 14887 22021
rect 14829 22012 14841 22015
rect 14792 21984 14841 22012
rect 14792 21972 14798 21984
rect 14829 21981 14841 21984
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 15746 21972 15752 22024
rect 15804 22012 15810 22024
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15804 21984 15853 22012
rect 15804 21972 15810 21984
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 16132 22012 16160 22043
rect 16942 22012 16948 22024
rect 16132 21984 16948 22012
rect 15841 21975 15899 21981
rect 16942 21972 16948 21984
rect 17000 22012 17006 22024
rect 17880 22012 17908 22052
rect 19352 22024 19380 22052
rect 19720 22052 20260 22080
rect 17000 21984 17908 22012
rect 17000 21972 17006 21984
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18932 21984 19257 22012
rect 18932 21972 18938 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 19334 21972 19340 22024
rect 19392 21972 19398 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19720 22012 19748 22052
rect 20254 22040 20260 22052
rect 20312 22040 20318 22092
rect 19484 21984 19748 22012
rect 19484 21972 19490 21984
rect 19886 21972 19892 22024
rect 19944 22012 19950 22024
rect 20364 22021 20392 22120
rect 20438 22108 20444 22120
rect 20496 22108 20502 22160
rect 21082 22040 21088 22092
rect 21140 22080 21146 22092
rect 21376 22080 21404 22188
rect 21140 22052 21404 22080
rect 22572 22094 22600 22188
rect 22738 22176 22744 22228
rect 22796 22176 22802 22228
rect 22830 22176 22836 22228
rect 22888 22176 22894 22228
rect 23477 22219 23535 22225
rect 23477 22185 23489 22219
rect 23523 22216 23535 22219
rect 26326 22216 26332 22228
rect 23523 22188 26332 22216
rect 23523 22185 23535 22188
rect 23477 22179 23535 22185
rect 26326 22176 26332 22188
rect 26384 22176 26390 22228
rect 23566 22148 23572 22160
rect 23124 22120 23572 22148
rect 23124 22094 23152 22120
rect 23566 22108 23572 22120
rect 23624 22108 23630 22160
rect 22572 22080 23152 22094
rect 23201 22083 23259 22089
rect 23201 22080 23213 22083
rect 22572 22066 23213 22080
rect 23124 22052 23213 22066
rect 21140 22040 21146 22052
rect 23201 22049 23213 22052
rect 23247 22049 23259 22083
rect 23201 22043 23259 22049
rect 24504 22052 25268 22080
rect 20349 22015 20407 22021
rect 19944 21984 20300 22012
rect 19944 21972 19950 21984
rect 12437 21947 12495 21953
rect 12437 21944 12449 21947
rect 11440 21916 12449 21944
rect 11296 21907 11325 21913
rect 12437 21913 12449 21916
rect 12483 21913 12495 21947
rect 12437 21907 12495 21913
rect 11296 21904 11302 21907
rect 12526 21904 12532 21956
rect 12584 21904 12590 21956
rect 13170 21904 13176 21956
rect 13228 21904 13234 21956
rect 16384 21947 16442 21953
rect 13648 21916 15332 21944
rect 7432 21848 10364 21876
rect 7432 21836 7438 21848
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 11606 21876 11612 21888
rect 11112 21848 11612 21876
rect 11112 21836 11118 21848
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 11882 21836 11888 21888
rect 11940 21836 11946 21888
rect 12237 21879 12295 21885
rect 12237 21845 12249 21879
rect 12283 21876 12295 21879
rect 12544 21876 12572 21904
rect 13648 21885 13676 21916
rect 15304 21888 15332 21916
rect 16384 21913 16396 21947
rect 16430 21944 16442 21947
rect 16666 21944 16672 21956
rect 16430 21916 16672 21944
rect 16430 21913 16442 21916
rect 16384 21907 16442 21913
rect 16666 21904 16672 21916
rect 16724 21904 16730 21956
rect 17770 21904 17776 21956
rect 17828 21953 17834 21956
rect 17828 21947 17891 21953
rect 17828 21913 17845 21947
rect 17879 21913 17891 21947
rect 17828 21907 17891 21913
rect 18049 21947 18107 21953
rect 18049 21913 18061 21947
rect 18095 21944 18107 21947
rect 18322 21944 18328 21956
rect 18095 21916 18328 21944
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 17828 21904 17834 21907
rect 18322 21904 18328 21916
rect 18380 21944 18386 21956
rect 19518 21944 19524 21956
rect 18380 21916 19524 21944
rect 18380 21904 18386 21916
rect 19518 21904 19524 21916
rect 19576 21904 19582 21956
rect 19610 21904 19616 21956
rect 19668 21944 19674 21956
rect 19705 21947 19763 21953
rect 19705 21944 19717 21947
rect 19668 21916 19717 21944
rect 19668 21904 19674 21916
rect 19705 21913 19717 21916
rect 19751 21913 19763 21947
rect 19705 21907 19763 21913
rect 20073 21947 20131 21953
rect 20073 21913 20085 21947
rect 20119 21944 20131 21947
rect 20165 21947 20223 21953
rect 20165 21944 20177 21947
rect 20119 21916 20177 21944
rect 20119 21913 20131 21916
rect 20073 21907 20131 21913
rect 20165 21913 20177 21916
rect 20211 21913 20223 21947
rect 20272 21944 20300 21984
rect 20349 21981 20361 22015
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20809 22015 20867 22021
rect 20809 22012 20821 22015
rect 20579 21984 20821 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20809 21981 20821 21984
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 22012 21419 22015
rect 22922 22012 22928 22024
rect 21407 21984 22928 22012
rect 21407 21981 21419 21984
rect 21361 21975 21419 21981
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23014 21972 23020 22024
rect 23072 21972 23078 22024
rect 23290 21972 23296 22024
rect 23348 22012 23354 22024
rect 23348 21984 23704 22012
rect 23348 21972 23354 21984
rect 20272 21916 20760 21944
rect 20165 21907 20223 21913
rect 12283 21848 12572 21876
rect 13633 21879 13691 21885
rect 12283 21845 12295 21848
rect 12237 21839 12295 21845
rect 13633 21845 13645 21879
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 14642 21836 14648 21888
rect 14700 21836 14706 21888
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 15657 21879 15715 21885
rect 15657 21845 15669 21879
rect 15703 21876 15715 21879
rect 16298 21876 16304 21888
rect 15703 21848 16304 21876
rect 15703 21845 15715 21848
rect 15657 21839 15715 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 17494 21836 17500 21888
rect 17552 21836 17558 21888
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 17681 21879 17739 21885
rect 17681 21876 17693 21879
rect 17644 21848 17693 21876
rect 17644 21836 17650 21848
rect 17681 21845 17693 21848
rect 17727 21845 17739 21879
rect 17681 21839 17739 21845
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 19978 21876 19984 21888
rect 18012 21848 19984 21876
rect 18012 21836 18018 21848
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20088 21876 20116 21907
rect 20530 21876 20536 21888
rect 20088 21848 20536 21876
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20622 21836 20628 21888
rect 20680 21836 20686 21888
rect 20732 21876 20760 21916
rect 21450 21904 21456 21956
rect 21508 21944 21514 21956
rect 23676 21953 23704 21984
rect 21606 21947 21664 21953
rect 21606 21944 21618 21947
rect 21508 21916 21618 21944
rect 21508 21904 21514 21916
rect 21606 21913 21618 21916
rect 21652 21913 21664 21947
rect 23661 21947 23719 21953
rect 21606 21907 21664 21913
rect 22066 21916 23612 21944
rect 22066 21876 22094 21916
rect 20732 21848 22094 21876
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 23474 21885 23480 21888
rect 23293 21879 23351 21885
rect 23293 21876 23305 21879
rect 22704 21848 23305 21876
rect 22704 21836 22710 21848
rect 23293 21845 23305 21848
rect 23339 21845 23351 21879
rect 23293 21839 23351 21845
rect 23451 21879 23480 21885
rect 23451 21845 23463 21879
rect 23451 21839 23480 21845
rect 23474 21836 23480 21839
rect 23532 21836 23538 21888
rect 23584 21876 23612 21916
rect 23661 21913 23673 21947
rect 23707 21913 23719 21947
rect 23661 21907 23719 21913
rect 24504 21876 24532 22052
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 22012 24639 22015
rect 24946 22012 24952 22024
rect 24627 21984 24952 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25240 22012 25268 22052
rect 26237 22015 26295 22021
rect 25240 21984 26096 22012
rect 25970 21947 26028 21953
rect 25970 21944 25982 21947
rect 24780 21916 25982 21944
rect 24780 21885 24808 21916
rect 25970 21913 25982 21916
rect 26016 21913 26028 21947
rect 25970 21907 26028 21913
rect 23584 21848 24532 21876
rect 24765 21879 24823 21885
rect 24765 21845 24777 21879
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 24854 21836 24860 21888
rect 24912 21836 24918 21888
rect 26068 21876 26096 21984
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 26326 22012 26332 22024
rect 26283 21984 26332 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 26326 21972 26332 21984
rect 26384 21972 26390 22024
rect 26142 21904 26148 21956
rect 26200 21944 26206 21956
rect 26574 21947 26632 21953
rect 26574 21944 26586 21947
rect 26200 21916 26586 21944
rect 26200 21904 26206 21916
rect 26574 21913 26586 21916
rect 26620 21913 26632 21947
rect 26574 21907 26632 21913
rect 27709 21879 27767 21885
rect 27709 21876 27721 21879
rect 26068 21848 27721 21876
rect 27709 21845 27721 21848
rect 27755 21845 27767 21879
rect 27709 21839 27767 21845
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 2590 21672 2596 21684
rect 1780 21644 2596 21672
rect 1780 21545 1808 21644
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 2685 21675 2743 21681
rect 2685 21641 2697 21675
rect 2731 21672 2743 21675
rect 3050 21672 3056 21684
rect 2731 21644 3056 21672
rect 2731 21641 2743 21644
rect 2685 21635 2743 21641
rect 3050 21632 3056 21644
rect 3108 21632 3114 21684
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 3697 21675 3755 21681
rect 3697 21672 3709 21675
rect 3384 21644 3709 21672
rect 3384 21632 3390 21644
rect 3697 21641 3709 21644
rect 3743 21641 3755 21675
rect 4154 21672 4160 21684
rect 3697 21635 3755 21641
rect 3804 21644 4160 21672
rect 2222 21613 2228 21616
rect 2179 21607 2228 21613
rect 2179 21573 2191 21607
rect 2225 21573 2228 21607
rect 2179 21567 2228 21573
rect 2222 21564 2228 21567
rect 2280 21564 2286 21616
rect 2774 21613 2780 21616
rect 2766 21607 2780 21613
rect 2766 21573 2778 21607
rect 2766 21567 2780 21573
rect 2774 21564 2780 21567
rect 2832 21564 2838 21616
rect 2869 21607 2927 21613
rect 2869 21573 2881 21607
rect 2915 21604 2927 21607
rect 3237 21607 3295 21613
rect 3237 21604 3249 21607
rect 2915 21576 3249 21604
rect 2915 21573 2927 21576
rect 2869 21567 2927 21573
rect 3237 21573 3249 21576
rect 3283 21573 3295 21607
rect 3237 21567 3295 21573
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21536 2467 21539
rect 2501 21539 2559 21545
rect 2501 21536 2513 21539
rect 2455 21508 2513 21536
rect 2455 21505 2467 21508
rect 2409 21499 2467 21505
rect 2501 21505 2513 21508
rect 2547 21505 2559 21539
rect 3145 21539 3203 21545
rect 2501 21499 2559 21505
rect 2608 21508 2774 21536
rect 2130 21428 2136 21480
rect 2188 21468 2194 21480
rect 2608 21468 2636 21508
rect 2188 21440 2636 21468
rect 2746 21468 2774 21508
rect 3145 21505 3157 21539
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 3329 21539 3387 21545
rect 3329 21505 3341 21539
rect 3375 21536 3387 21539
rect 3804 21536 3832 21644
rect 4154 21632 4160 21644
rect 4212 21672 4218 21684
rect 4338 21672 4344 21684
rect 4212 21644 4344 21672
rect 4212 21632 4218 21644
rect 4338 21632 4344 21644
rect 4396 21632 4402 21684
rect 5442 21632 5448 21684
rect 5500 21672 5506 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5500 21644 5641 21672
rect 5500 21632 5506 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5997 21675 6055 21681
rect 5997 21672 6009 21675
rect 5629 21635 5687 21641
rect 5828 21644 6009 21672
rect 4065 21607 4123 21613
rect 4065 21573 4077 21607
rect 4111 21604 4123 21607
rect 5258 21604 5264 21616
rect 4111 21576 5264 21604
rect 4111 21573 4123 21576
rect 4065 21567 4123 21573
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 5828 21604 5856 21644
rect 5997 21641 6009 21644
rect 6043 21641 6055 21675
rect 5997 21635 6055 21641
rect 6454 21632 6460 21684
rect 6512 21632 6518 21684
rect 7466 21632 7472 21684
rect 7524 21672 7530 21684
rect 7524 21644 7604 21672
rect 7524 21632 7530 21644
rect 5644 21576 5856 21604
rect 3375 21508 3832 21536
rect 3876 21539 3934 21545
rect 3375 21505 3387 21508
rect 3329 21499 3387 21505
rect 3876 21505 3888 21539
rect 3922 21505 3934 21539
rect 3876 21499 3934 21505
rect 3160 21468 3188 21499
rect 2746 21440 3188 21468
rect 3896 21468 3924 21499
rect 3970 21496 3976 21548
rect 4028 21496 4034 21548
rect 4248 21539 4306 21545
rect 4248 21505 4260 21539
rect 4294 21505 4306 21539
rect 4248 21499 4306 21505
rect 4154 21468 4160 21480
rect 3896 21440 4160 21468
rect 2188 21428 2194 21440
rect 4154 21428 4160 21440
rect 4212 21428 4218 21480
rect 4264 21468 4292 21499
rect 4338 21496 4344 21548
rect 4396 21496 4402 21548
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4433 21471 4491 21477
rect 4433 21468 4445 21471
rect 4264 21440 4445 21468
rect 4433 21437 4445 21440
rect 4479 21437 4491 21471
rect 4433 21431 4491 21437
rect 1302 21360 1308 21412
rect 1360 21400 1366 21412
rect 3053 21403 3111 21409
rect 3053 21400 3065 21403
rect 1360 21372 3065 21400
rect 1360 21360 1366 21372
rect 3053 21369 3065 21372
rect 3099 21369 3111 21403
rect 3053 21363 3111 21369
rect 4246 21360 4252 21412
rect 4304 21400 4310 21412
rect 4632 21400 4660 21499
rect 4798 21496 4804 21548
rect 4856 21536 4862 21548
rect 5442 21536 5448 21548
rect 4856 21508 5448 21536
rect 4856 21496 4862 21508
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 5534 21496 5540 21548
rect 5592 21496 5598 21548
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 5350 21468 5356 21480
rect 4948 21440 5356 21468
rect 4948 21428 4954 21440
rect 5350 21428 5356 21440
rect 5408 21428 5414 21480
rect 5644 21468 5672 21576
rect 6178 21564 6184 21616
rect 6236 21564 6242 21616
rect 6730 21564 6736 21616
rect 6788 21564 6794 21616
rect 6825 21607 6883 21613
rect 6825 21573 6837 21607
rect 6871 21604 6883 21607
rect 7193 21607 7251 21613
rect 7193 21604 7205 21607
rect 6871 21576 7205 21604
rect 6871 21573 6883 21576
rect 6825 21567 6883 21573
rect 7193 21573 7205 21576
rect 7239 21573 7251 21607
rect 7193 21567 7251 21573
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 5552 21440 5672 21468
rect 5828 21468 5856 21499
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6196 21536 6224 21564
rect 6595 21539 6653 21545
rect 6595 21536 6607 21539
rect 6012 21508 6607 21536
rect 6012 21468 6040 21508
rect 6595 21505 6607 21508
rect 6641 21505 6653 21539
rect 6595 21499 6653 21505
rect 6953 21539 7011 21545
rect 6953 21505 6965 21539
rect 6999 21505 7011 21539
rect 6953 21499 7011 21505
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 5828 21440 6040 21468
rect 6108 21471 6166 21477
rect 5552 21412 5580 21440
rect 6108 21437 6120 21471
rect 6154 21468 6166 21471
rect 6968 21468 6996 21499
rect 6154 21440 6996 21468
rect 7116 21468 7144 21499
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 7340 21508 7389 21536
rect 7340 21496 7346 21508
rect 7377 21505 7389 21508
rect 7423 21505 7435 21539
rect 7466 21530 7472 21582
rect 7524 21530 7530 21582
rect 7576 21536 7604 21644
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 8573 21675 8631 21681
rect 8573 21672 8585 21675
rect 8536 21644 8585 21672
rect 8536 21632 8542 21644
rect 8573 21641 8585 21644
rect 8619 21641 8631 21675
rect 9398 21672 9404 21684
rect 8573 21635 8631 21641
rect 8680 21644 9404 21672
rect 8294 21604 8300 21616
rect 7944 21576 8300 21604
rect 7944 21545 7972 21576
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7377 21499 7435 21505
rect 7469 21505 7481 21530
rect 7515 21505 7527 21530
rect 7576 21508 7665 21536
rect 7469 21499 7527 21505
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7791 21508 7941 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21536 8263 21539
rect 8251 21508 8432 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 7190 21468 7196 21480
rect 7116 21440 7196 21468
rect 6154 21437 6166 21440
rect 6108 21431 6166 21437
rect 4304 21372 4660 21400
rect 4304 21360 4310 21372
rect 5534 21360 5540 21412
rect 5592 21360 5598 21412
rect 5813 21403 5871 21409
rect 5813 21369 5825 21403
rect 5859 21369 5871 21403
rect 5813 21363 5871 21369
rect 2133 21335 2191 21341
rect 2133 21301 2145 21335
rect 2179 21332 2191 21335
rect 2314 21332 2320 21344
rect 2179 21304 2320 21332
rect 2179 21301 2191 21304
rect 2133 21295 2191 21301
rect 2314 21292 2320 21304
rect 2372 21332 2378 21344
rect 3234 21332 3240 21344
rect 2372 21304 3240 21332
rect 2372 21292 2378 21304
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 4798 21292 4804 21344
rect 4856 21292 4862 21344
rect 5828 21332 5856 21363
rect 5902 21360 5908 21412
rect 5960 21400 5966 21412
rect 7116 21400 7144 21440
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 5960 21372 7144 21400
rect 5960 21360 5966 21372
rect 6914 21332 6920 21344
rect 5828 21304 6920 21332
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 7392 21332 7420 21499
rect 7558 21428 7564 21480
rect 7616 21428 7622 21480
rect 7576 21400 7604 21428
rect 7929 21403 7987 21409
rect 7929 21400 7941 21403
rect 7576 21372 7941 21400
rect 7929 21369 7941 21372
rect 7975 21369 7987 21403
rect 8128 21400 8156 21499
rect 8404 21480 8432 21508
rect 8478 21496 8484 21548
rect 8536 21496 8542 21548
rect 8680 21545 8708 21644
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 9766 21672 9772 21684
rect 9539 21644 9772 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 9876 21644 10732 21672
rect 9876 21616 9904 21644
rect 8956 21576 9812 21604
rect 8956 21545 8984 21576
rect 9784 21545 9812 21576
rect 9858 21564 9864 21616
rect 9916 21564 9922 21616
rect 10428 21576 10640 21604
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 8757 21539 8815 21545
rect 8757 21505 8769 21539
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21536 9367 21539
rect 9769 21539 9827 21545
rect 9355 21508 9720 21536
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 8386 21428 8392 21480
rect 8444 21468 8450 21480
rect 8772 21468 8800 21499
rect 8444 21440 8800 21468
rect 9125 21471 9183 21477
rect 8444 21428 8450 21440
rect 9125 21437 9137 21471
rect 9171 21468 9183 21471
rect 9582 21468 9588 21480
rect 9171 21440 9588 21468
rect 9171 21437 9183 21440
rect 9125 21431 9183 21437
rect 9582 21428 9588 21440
rect 9640 21428 9646 21480
rect 9692 21400 9720 21508
rect 9769 21505 9781 21539
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 9784 21468 9812 21499
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 10008 21508 10057 21536
rect 10008 21496 10014 21508
rect 10045 21505 10057 21508
rect 10091 21536 10103 21539
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 10091 21508 10241 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10229 21505 10241 21508
rect 10275 21505 10287 21539
rect 10229 21499 10287 21505
rect 10428 21468 10456 21576
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 9784 21440 10456 21468
rect 9766 21400 9772 21412
rect 8128 21372 9168 21400
rect 9692 21372 9772 21400
rect 7929 21363 7987 21369
rect 9140 21344 9168 21372
rect 9766 21360 9772 21372
rect 9824 21360 9830 21412
rect 9858 21360 9864 21412
rect 9916 21360 9922 21412
rect 9953 21403 10011 21409
rect 9953 21369 9965 21403
rect 9999 21400 10011 21403
rect 10520 21400 10548 21499
rect 10612 21468 10640 21576
rect 10704 21545 10732 21644
rect 10962 21632 10968 21684
rect 11020 21672 11026 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 11020 21644 12081 21672
rect 11020 21632 11026 21644
rect 12069 21641 12081 21644
rect 12115 21672 12127 21675
rect 12526 21672 12532 21684
rect 12115 21644 12532 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 16666 21632 16672 21684
rect 16724 21632 16730 21684
rect 17954 21632 17960 21684
rect 18012 21632 18018 21684
rect 19179 21675 19237 21681
rect 19179 21641 19191 21675
rect 19225 21672 19237 21675
rect 19426 21672 19432 21684
rect 19225 21644 19432 21672
rect 19225 21641 19237 21644
rect 19179 21635 19237 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 19518 21632 19524 21684
rect 19576 21632 19582 21684
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 23474 21672 23480 21684
rect 20312 21644 23480 21672
rect 20312 21632 20318 21644
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 26142 21672 26148 21684
rect 26007 21644 26148 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 10980 21576 12020 21604
rect 10980 21545 11008 21576
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 10980 21468 11008 21499
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 11112 21508 11529 21536
rect 11112 21496 11118 21508
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 10612 21440 11008 21468
rect 11793 21471 11851 21477
rect 11793 21437 11805 21471
rect 11839 21468 11851 21471
rect 11882 21468 11888 21480
rect 11839 21440 11888 21468
rect 11839 21437 11851 21440
rect 11793 21431 11851 21437
rect 9999 21372 10548 21400
rect 10597 21403 10655 21409
rect 9999 21369 10011 21372
rect 9953 21363 10011 21369
rect 10597 21369 10609 21403
rect 10643 21400 10655 21403
rect 11808 21400 11836 21431
rect 11882 21428 11888 21440
rect 11940 21428 11946 21480
rect 11992 21468 12020 21576
rect 12912 21576 14596 21604
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 12802 21536 12808 21548
rect 12391 21508 12808 21536
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 12912 21545 12940 21576
rect 13170 21545 13176 21548
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21505 12955 21539
rect 12897 21499 12955 21505
rect 13164 21499 13176 21545
rect 13170 21496 13176 21499
rect 13228 21496 13234 21548
rect 14568 21480 14596 21576
rect 14642 21564 14648 21616
rect 14700 21604 14706 21616
rect 14798 21607 14856 21613
rect 14798 21604 14810 21607
rect 14700 21576 14810 21604
rect 14700 21564 14706 21576
rect 14798 21573 14810 21576
rect 14844 21573 14856 21607
rect 14798 21567 14856 21573
rect 15654 21564 15660 21616
rect 15712 21604 15718 21616
rect 16025 21607 16083 21613
rect 16025 21604 16037 21607
rect 15712 21576 16037 21604
rect 15712 21564 15718 21576
rect 16025 21573 16037 21576
rect 16071 21604 16083 21607
rect 17972 21604 18000 21632
rect 16071 21576 18000 21604
rect 18969 21607 19027 21613
rect 16071 21573 16083 21576
rect 16025 21567 16083 21573
rect 18969 21573 18981 21607
rect 19015 21604 19027 21607
rect 19536 21604 19564 21632
rect 20340 21607 20398 21613
rect 19015 21576 19196 21604
rect 19536 21576 20300 21604
rect 19015 21573 19027 21576
rect 18969 21567 19027 21573
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21536 16267 21539
rect 16298 21536 16304 21548
rect 16255 21508 16304 21536
rect 16255 21505 16267 21508
rect 16209 21499 16267 21505
rect 12526 21468 12532 21480
rect 11992 21440 12532 21468
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 10643 21372 11836 21400
rect 15933 21403 15991 21409
rect 10643 21369 10655 21372
rect 10597 21363 10655 21369
rect 15933 21369 15945 21403
rect 15979 21400 15991 21403
rect 16224 21400 16252 21499
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 16393 21539 16451 21545
rect 16393 21505 16405 21539
rect 16439 21536 16451 21539
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16439 21508 16865 21536
rect 16439 21505 16451 21508
rect 16393 21499 16451 21505
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17276 21508 17509 21536
rect 17276 21496 17282 21508
rect 17497 21505 17509 21508
rect 17543 21536 17555 21539
rect 17678 21536 17684 21548
rect 17543 21508 17684 21536
rect 17543 21505 17555 21508
rect 17497 21499 17555 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18141 21539 18199 21545
rect 18141 21536 18153 21539
rect 17819 21508 18153 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18141 21505 18153 21508
rect 18187 21536 18199 21539
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 18187 21508 18613 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18601 21505 18613 21508
rect 18647 21536 18659 21539
rect 19168 21536 19196 21576
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 18647 21508 19533 21536
rect 18647 21505 18659 21508
rect 18601 21499 18659 21505
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21468 17647 21471
rect 17788 21468 17816 21499
rect 19168 21480 19196 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20272 21536 20300 21576
rect 20340 21573 20352 21607
rect 20386 21604 20398 21607
rect 20622 21604 20628 21616
rect 20386 21576 20628 21604
rect 20386 21573 20398 21576
rect 20340 21567 20398 21573
rect 20622 21564 20628 21576
rect 20680 21564 20686 21616
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 22129 21607 22187 21613
rect 21959 21576 21993 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 22129 21573 22141 21607
rect 22175 21604 22187 21607
rect 22278 21604 22284 21616
rect 22175 21576 22284 21604
rect 22175 21573 22187 21576
rect 22129 21567 22187 21573
rect 21928 21536 21956 21567
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22756 21576 23152 21604
rect 22756 21548 22784 21576
rect 20272 21508 22692 21536
rect 18322 21468 18328 21480
rect 17635 21440 17816 21468
rect 17972 21440 18328 21468
rect 17635 21437 17647 21440
rect 17589 21431 17647 21437
rect 15979 21372 16252 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 7558 21332 7564 21344
rect 7392 21304 7564 21332
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 8849 21335 8907 21341
rect 8849 21332 8861 21335
rect 7708 21304 8861 21332
rect 7708 21292 7714 21304
rect 8849 21301 8861 21304
rect 8895 21301 8907 21335
rect 8849 21295 8907 21301
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 9968 21332 9996 21363
rect 9180 21304 9996 21332
rect 9180 21292 9186 21304
rect 10778 21292 10784 21344
rect 10836 21332 10842 21344
rect 11609 21335 11667 21341
rect 11609 21332 11621 21335
rect 10836 21304 11621 21332
rect 10836 21292 10842 21304
rect 11609 21301 11621 21304
rect 11655 21332 11667 21335
rect 11790 21332 11796 21344
rect 11655 21304 11796 21332
rect 11655 21301 11667 21304
rect 11609 21295 11667 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12529 21335 12587 21341
rect 12529 21301 12541 21335
rect 12575 21332 12587 21335
rect 12894 21332 12900 21344
rect 12575 21304 12900 21332
rect 12575 21301 12587 21304
rect 12529 21295 12587 21301
rect 12894 21292 12900 21304
rect 12952 21332 12958 21344
rect 13630 21332 13636 21344
rect 12952 21304 13636 21332
rect 12952 21292 12958 21304
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 14277 21335 14335 21341
rect 14277 21301 14289 21335
rect 14323 21332 14335 21335
rect 14826 21332 14832 21344
rect 14323 21304 14832 21332
rect 14323 21301 14335 21304
rect 14277 21295 14335 21301
rect 14826 21292 14832 21304
rect 14884 21292 14890 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17972 21341 18000 21440
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 19150 21428 19156 21480
rect 19208 21428 19214 21480
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21468 19763 21471
rect 19794 21468 19800 21480
rect 19751 21440 19800 21468
rect 19751 21437 19763 21440
rect 19705 21431 19763 21437
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 19904 21400 19932 21496
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21437 20131 21471
rect 22554 21468 22560 21480
rect 20073 21431 20131 21437
rect 22112 21440 22560 21468
rect 19168 21372 19932 21400
rect 17957 21335 18015 21341
rect 17957 21332 17969 21335
rect 16632 21304 17969 21332
rect 16632 21292 16638 21304
rect 17957 21301 17969 21304
rect 18003 21301 18015 21335
rect 17957 21295 18015 21301
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18325 21335 18383 21341
rect 18325 21332 18337 21335
rect 18196 21304 18337 21332
rect 18196 21292 18202 21304
rect 18325 21301 18337 21304
rect 18371 21301 18383 21335
rect 18325 21295 18383 21301
rect 18693 21335 18751 21341
rect 18693 21301 18705 21335
rect 18739 21332 18751 21335
rect 18874 21332 18880 21344
rect 18739 21304 18880 21332
rect 18739 21301 18751 21304
rect 18693 21295 18751 21301
rect 18874 21292 18880 21304
rect 18932 21292 18938 21344
rect 19168 21341 19196 21372
rect 19153 21335 19211 21341
rect 19153 21301 19165 21335
rect 19199 21301 19211 21335
rect 19153 21295 19211 21301
rect 19334 21292 19340 21344
rect 19392 21292 19398 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19886 21332 19892 21344
rect 19484 21304 19892 21332
rect 19484 21292 19490 21304
rect 19886 21292 19892 21304
rect 19944 21332 19950 21344
rect 20088 21332 20116 21431
rect 19944 21304 20116 21332
rect 19944 21292 19950 21304
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 22112 21341 22140 21440
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 22664 21468 22692 21508
rect 22738 21496 22744 21548
rect 22796 21496 22802 21548
rect 23124 21545 23152 21576
rect 23198 21564 23204 21616
rect 23256 21564 23262 21616
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23109 21539 23167 21545
rect 23109 21505 23121 21539
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 22940 21468 22968 21499
rect 25774 21496 25780 21548
rect 25832 21496 25838 21548
rect 24854 21468 24860 21480
rect 22664 21440 22876 21468
rect 22940 21440 24860 21468
rect 22281 21403 22339 21409
rect 22281 21369 22293 21403
rect 22327 21400 22339 21403
rect 22741 21403 22799 21409
rect 22741 21400 22753 21403
rect 22327 21372 22753 21400
rect 22327 21369 22339 21372
rect 22281 21363 22339 21369
rect 22741 21369 22753 21372
rect 22787 21369 22799 21403
rect 22848 21400 22876 21440
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 22848 21372 22968 21400
rect 22741 21363 22799 21369
rect 21453 21335 21511 21341
rect 21453 21332 21465 21335
rect 21324 21304 21465 21332
rect 21324 21292 21330 21304
rect 21453 21301 21465 21304
rect 21499 21301 21511 21335
rect 21453 21295 21511 21301
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21301 22155 21335
rect 22097 21295 22155 21301
rect 22370 21292 22376 21344
rect 22428 21292 22434 21344
rect 22646 21292 22652 21344
rect 22704 21292 22710 21344
rect 22830 21292 22836 21344
rect 22888 21292 22894 21344
rect 22940 21332 22968 21372
rect 23106 21360 23112 21412
rect 23164 21400 23170 21412
rect 23477 21403 23535 21409
rect 23477 21400 23489 21403
rect 23164 21372 23489 21400
rect 23164 21360 23170 21372
rect 23477 21369 23489 21372
rect 23523 21369 23535 21403
rect 23477 21363 23535 21369
rect 23198 21332 23204 21344
rect 22940 21304 23204 21332
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 23658 21292 23664 21344
rect 23716 21292 23722 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 2225 21131 2283 21137
rect 2225 21097 2237 21131
rect 2271 21128 2283 21131
rect 2406 21128 2412 21140
rect 2271 21100 2412 21128
rect 2271 21097 2283 21100
rect 2225 21091 2283 21097
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 2774 21088 2780 21140
rect 2832 21128 2838 21140
rect 4709 21131 4767 21137
rect 4709 21128 4721 21131
rect 2832 21100 4721 21128
rect 2832 21088 2838 21100
rect 4709 21097 4721 21100
rect 4755 21097 4767 21131
rect 4709 21091 4767 21097
rect 4890 21088 4896 21140
rect 4948 21128 4954 21140
rect 4948 21100 5396 21128
rect 4948 21088 4954 21100
rect 3050 21060 3056 21072
rect 2240 21032 3056 21060
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2240 20924 2268 21032
rect 3050 21020 3056 21032
rect 3108 21020 3114 21072
rect 3145 21063 3203 21069
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 3510 21060 3516 21072
rect 3191 21032 3516 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 3510 21020 3516 21032
rect 3568 21020 3574 21072
rect 2682 20952 2688 21004
rect 2740 20952 2746 21004
rect 2792 20964 3188 20992
rect 2087 20896 2268 20924
rect 2317 20927 2375 20933
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 2317 20893 2329 20927
rect 2363 20924 2375 20927
rect 2792 20924 2820 20964
rect 3160 20936 3188 20964
rect 3234 20952 3240 21004
rect 3292 20952 3298 21004
rect 2363 20896 2820 20924
rect 2869 20927 2927 20933
rect 2363 20893 2375 20896
rect 2317 20887 2375 20893
rect 2869 20893 2881 20927
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 2884 20856 2912 20887
rect 3142 20884 3148 20936
rect 3200 20884 3206 20936
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 4847 20927 4905 20933
rect 4847 20924 4859 20927
rect 4212 20896 4859 20924
rect 4212 20884 4218 20896
rect 4847 20893 4859 20896
rect 4893 20893 4905 20927
rect 4847 20887 4905 20893
rect 5166 20884 5172 20936
rect 5224 20933 5230 20936
rect 5368 20933 5396 21100
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 6270 21128 6276 21140
rect 5592 21100 6276 21128
rect 5592 21088 5598 21100
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 7009 21131 7067 21137
rect 7009 21097 7021 21131
rect 7055 21128 7067 21131
rect 7098 21128 7104 21140
rect 7055 21100 7104 21128
rect 7055 21097 7067 21100
rect 7009 21091 7067 21097
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 7190 21088 7196 21140
rect 7248 21128 7254 21140
rect 8573 21131 8631 21137
rect 7248 21100 7880 21128
rect 7248 21088 7254 21100
rect 6196 20964 6771 20992
rect 6196 20936 6224 20964
rect 5224 20927 5273 20933
rect 5224 20893 5227 20927
rect 5261 20893 5273 20927
rect 5224 20887 5273 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 5224 20884 5230 20887
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 6638 20924 6644 20936
rect 6599 20896 6644 20924
rect 6638 20884 6644 20896
rect 6696 20884 6702 20936
rect 6743 20924 6771 20964
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7101 20995 7159 21001
rect 7101 20992 7113 20995
rect 6972 20964 7113 20992
rect 6972 20952 6978 20964
rect 7101 20961 7113 20964
rect 7147 20961 7159 20995
rect 7101 20955 7159 20961
rect 7331 20927 7389 20933
rect 7331 20924 7343 20927
rect 6743 20896 7343 20924
rect 7331 20893 7343 20896
rect 7377 20893 7389 20927
rect 7331 20887 7389 20893
rect 7466 20884 7472 20936
rect 7524 20884 7530 20936
rect 7650 20884 7656 20936
rect 7708 20933 7714 20936
rect 7852 20933 7880 21100
rect 8573 21097 8585 21131
rect 8619 21097 8631 21131
rect 8573 21091 8631 21097
rect 8588 21060 8616 21091
rect 8754 21088 8760 21140
rect 8812 21088 8818 21140
rect 9122 21088 9128 21140
rect 9180 21088 9186 21140
rect 10428 21100 11008 21128
rect 8846 21060 8852 21072
rect 8588 21032 8852 21060
rect 8846 21020 8852 21032
rect 8904 21020 8910 21072
rect 9490 21020 9496 21072
rect 9548 21060 9554 21072
rect 9858 21060 9864 21072
rect 9548 21032 9864 21060
rect 9548 21020 9554 21032
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 8205 20995 8263 21001
rect 8205 20961 8217 20995
rect 8251 20992 8263 20995
rect 9398 20992 9404 21004
rect 8251 20964 9404 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 9398 20952 9404 20964
rect 9456 20992 9462 21004
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9456 20964 9689 20992
rect 9456 20952 9462 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 7708 20927 7747 20933
rect 7735 20893 7747 20927
rect 7708 20887 7747 20893
rect 7837 20927 7895 20933
rect 7837 20893 7849 20927
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 7708 20884 7714 20887
rect 9214 20884 9220 20936
rect 9272 20924 9278 20936
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 9272 20896 9505 20924
rect 9272 20884 9278 20896
rect 9493 20893 9505 20896
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 9640 20896 10333 20924
rect 9640 20884 9646 20896
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 4706 20856 4712 20868
rect 2884 20828 4712 20856
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 4985 20859 5043 20865
rect 4985 20825 4997 20859
rect 5031 20825 5043 20859
rect 4985 20819 5043 20825
rect 5077 20859 5135 20865
rect 5077 20825 5089 20859
rect 5123 20825 5135 20859
rect 7561 20859 7619 20865
rect 5077 20819 5135 20825
rect 5460 20828 7236 20856
rect 1857 20791 1915 20797
rect 1857 20757 1869 20791
rect 1903 20788 1915 20791
rect 2314 20788 2320 20800
rect 1903 20760 2320 20788
rect 1903 20757 1915 20760
rect 1857 20751 1915 20757
rect 2314 20748 2320 20760
rect 2372 20748 2378 20800
rect 4614 20748 4620 20800
rect 4672 20788 4678 20800
rect 5000 20788 5028 20819
rect 4672 20760 5028 20788
rect 5092 20788 5120 20819
rect 5460 20788 5488 20828
rect 5092 20760 5488 20788
rect 4672 20748 4678 20760
rect 5810 20748 5816 20800
rect 5868 20788 5874 20800
rect 6457 20791 6515 20797
rect 6457 20788 6469 20791
rect 5868 20760 6469 20788
rect 5868 20748 5874 20760
rect 6457 20757 6469 20760
rect 6503 20757 6515 20791
rect 6457 20751 6515 20757
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 7208 20797 7236 20828
rect 7561 20825 7573 20859
rect 7607 20856 7619 20859
rect 8754 20856 8760 20868
rect 7607 20828 8760 20856
rect 7607 20825 7619 20828
rect 7561 20819 7619 20825
rect 8754 20816 8760 20828
rect 8812 20816 8818 20868
rect 8846 20816 8852 20868
rect 8904 20856 8910 20868
rect 10428 20856 10456 21100
rect 10873 21063 10931 21069
rect 10873 21029 10885 21063
rect 10919 21029 10931 21063
rect 10980 21060 11008 21100
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13357 21131 13415 21137
rect 13357 21128 13369 21131
rect 13228 21100 13369 21128
rect 13228 21088 13234 21100
rect 13357 21097 13369 21100
rect 13403 21097 13415 21131
rect 13357 21091 13415 21097
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 14921 21131 14979 21137
rect 14921 21128 14933 21131
rect 14792 21100 14933 21128
rect 14792 21088 14798 21100
rect 14921 21097 14933 21100
rect 14967 21097 14979 21131
rect 14921 21091 14979 21097
rect 15194 21088 15200 21140
rect 15252 21088 15258 21140
rect 15841 21131 15899 21137
rect 15841 21097 15853 21131
rect 15887 21097 15899 21131
rect 15841 21091 15899 21097
rect 17129 21131 17187 21137
rect 17129 21097 17141 21131
rect 17175 21128 17187 21131
rect 17494 21128 17500 21140
rect 17175 21100 17500 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 12802 21060 12808 21072
rect 10980 21032 12808 21060
rect 10873 21023 10931 21029
rect 10888 20992 10916 21023
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 14826 21020 14832 21072
rect 14884 21060 14890 21072
rect 15856 21060 15884 21091
rect 17494 21088 17500 21100
rect 17552 21088 17558 21140
rect 18690 21088 18696 21140
rect 18748 21088 18754 21140
rect 19150 21128 19156 21140
rect 19076 21100 19156 21128
rect 14884 21032 15884 21060
rect 14884 21020 14890 21032
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 10888 20964 11161 20992
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 12066 20952 12072 21004
rect 12124 20952 12130 21004
rect 19076 21001 19104 21100
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19521 21131 19579 21137
rect 19521 21128 19533 21131
rect 19392 21100 19533 21128
rect 19392 21088 19398 21100
rect 19521 21097 19533 21100
rect 19567 21097 19579 21131
rect 19521 21091 19579 21097
rect 20533 21131 20591 21137
rect 20533 21097 20545 21131
rect 20579 21128 20591 21131
rect 21174 21128 21180 21140
rect 20579 21100 21180 21128
rect 20579 21097 20591 21100
rect 20533 21091 20591 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 21450 21088 21456 21140
rect 21508 21088 21514 21140
rect 22830 21088 22836 21140
rect 22888 21088 22894 21140
rect 23017 21131 23075 21137
rect 23017 21097 23029 21131
rect 23063 21128 23075 21131
rect 23106 21128 23112 21140
rect 23063 21100 23112 21128
rect 23063 21097 23075 21100
rect 23017 21091 23075 21097
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 23658 21088 23664 21140
rect 23716 21088 23722 21140
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 24912 21100 24992 21128
rect 24912 21088 24918 21100
rect 19242 21020 19248 21072
rect 19300 21060 19306 21072
rect 19613 21063 19671 21069
rect 19613 21060 19625 21063
rect 19300 21032 19625 21060
rect 19300 21020 19306 21032
rect 19613 21029 19625 21032
rect 19659 21029 19671 21063
rect 19613 21023 19671 21029
rect 20438 21020 20444 21072
rect 20496 21060 20502 21072
rect 20496 21032 23520 21060
rect 20496 21020 20502 21032
rect 19061 20995 19119 21001
rect 14292 20964 17954 20992
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10778 20924 10784 20936
rect 10735 20896 10784 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 13538 20884 13544 20936
rect 13596 20884 13602 20936
rect 14292 20933 14320 20964
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 14016 20896 14289 20924
rect 8904 20828 10456 20856
rect 10505 20859 10563 20865
rect 8904 20816 8910 20828
rect 10505 20825 10517 20859
rect 10551 20825 10563 20859
rect 10505 20819 10563 20825
rect 10597 20859 10655 20865
rect 10597 20825 10609 20859
rect 10643 20856 10655 20859
rect 11698 20856 11704 20868
rect 10643 20828 11704 20856
rect 10643 20825 10655 20828
rect 10597 20819 10655 20825
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 6604 20760 6653 20788
rect 6604 20748 6610 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 7193 20791 7251 20797
rect 7193 20757 7205 20791
rect 7239 20757 7251 20791
rect 7193 20751 7251 20757
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 8573 20791 8631 20797
rect 8573 20788 8585 20791
rect 7432 20760 8585 20788
rect 7432 20748 7438 20760
rect 8573 20757 8585 20760
rect 8619 20757 8631 20791
rect 8573 20751 8631 20757
rect 9582 20748 9588 20800
rect 9640 20748 9646 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 10520 20788 10548 20819
rect 11698 20816 11704 20828
rect 11756 20816 11762 20868
rect 12897 20859 12955 20865
rect 12897 20825 12909 20859
rect 12943 20856 12955 20859
rect 13354 20856 13360 20868
rect 12943 20828 13360 20856
rect 12943 20825 12955 20828
rect 12897 20819 12955 20825
rect 13354 20816 13360 20828
rect 13412 20816 13418 20868
rect 14016 20800 14044 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 14826 20924 14832 20936
rect 14783 20896 14832 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 15013 20927 15071 20933
rect 15013 20893 15025 20927
rect 15059 20893 15071 20927
rect 15013 20887 15071 20893
rect 14366 20816 14372 20868
rect 14424 20856 14430 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 14424 20828 14565 20856
rect 14424 20816 14430 20828
rect 14553 20825 14565 20828
rect 14599 20856 14611 20859
rect 14642 20856 14648 20868
rect 14599 20828 14648 20856
rect 14599 20825 14611 20828
rect 14553 20819 14611 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 15028 20856 15056 20887
rect 15470 20884 15476 20936
rect 15528 20924 15534 20936
rect 16574 20924 16580 20936
rect 15528 20896 16580 20924
rect 15528 20884 15534 20896
rect 16574 20884 16580 20896
rect 16632 20924 16638 20936
rect 17926 20924 17954 20964
rect 19061 20961 19073 20995
rect 19107 20961 19119 20995
rect 19061 20955 19119 20961
rect 19978 20952 19984 21004
rect 20036 20992 20042 21004
rect 20346 20992 20352 21004
rect 20036 20964 20352 20992
rect 20036 20952 20042 20964
rect 20346 20952 20352 20964
rect 20404 20992 20410 21004
rect 20404 20964 20852 20992
rect 20404 20952 20410 20964
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 16632 20896 16988 20924
rect 17926 20896 18889 20924
rect 16632 20884 16638 20896
rect 14752 20828 15056 20856
rect 15657 20859 15715 20865
rect 14752 20800 14780 20828
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16114 20856 16120 20868
rect 15703 20828 16120 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16482 20816 16488 20868
rect 16540 20856 16546 20868
rect 16960 20865 16988 20896
rect 18877 20893 18889 20896
rect 18923 20924 18935 20927
rect 18966 20924 18972 20936
rect 18923 20896 18972 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19242 20927 19300 20933
rect 19242 20924 19254 20927
rect 19076 20896 19254 20924
rect 16945 20859 17003 20865
rect 16540 20828 16896 20856
rect 16540 20816 16546 20828
rect 11054 20788 11060 20800
rect 9824 20760 11060 20788
rect 9824 20748 9830 20760
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 12986 20748 12992 20800
rect 13044 20748 13050 20800
rect 13998 20748 14004 20800
rect 14056 20748 14062 20800
rect 14090 20748 14096 20800
rect 14148 20748 14154 20800
rect 14734 20748 14740 20800
rect 14792 20748 14798 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15857 20791 15915 20797
rect 15857 20788 15869 20791
rect 15252 20760 15869 20788
rect 15252 20748 15258 20760
rect 15857 20757 15869 20760
rect 15903 20757 15915 20791
rect 15857 20751 15915 20757
rect 16025 20791 16083 20797
rect 16025 20757 16037 20791
rect 16071 20788 16083 20791
rect 16758 20788 16764 20800
rect 16071 20760 16764 20788
rect 16071 20757 16083 20760
rect 16025 20751 16083 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 16868 20788 16896 20828
rect 16945 20825 16957 20859
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 18690 20816 18696 20868
rect 18748 20856 18754 20868
rect 19076 20856 19104 20896
rect 19242 20893 19254 20896
rect 19288 20893 19300 20927
rect 19242 20887 19300 20893
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 20824 20933 20852 20964
rect 20916 20964 22232 20992
rect 19705 20927 19763 20933
rect 19705 20924 19717 20927
rect 19392 20896 19717 20924
rect 19392 20884 19398 20896
rect 19705 20893 19717 20896
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 20809 20927 20867 20933
rect 20809 20893 20821 20927
rect 20855 20893 20867 20927
rect 20809 20887 20867 20893
rect 20916 20868 20944 20964
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20924 21235 20927
rect 21269 20927 21327 20933
rect 21269 20924 21281 20927
rect 21223 20896 21281 20924
rect 21223 20893 21235 20896
rect 21177 20887 21235 20893
rect 21269 20893 21281 20896
rect 21315 20893 21327 20927
rect 21269 20887 21327 20893
rect 18748 20828 19104 20856
rect 18748 20816 18754 20828
rect 19518 20816 19524 20868
rect 19576 20856 19582 20868
rect 20349 20859 20407 20865
rect 20349 20856 20361 20859
rect 19576 20828 20361 20856
rect 19576 20816 19582 20828
rect 20349 20825 20361 20828
rect 20395 20825 20407 20859
rect 20349 20819 20407 20825
rect 20898 20816 20904 20868
rect 20956 20816 20962 20868
rect 20993 20859 21051 20865
rect 20993 20825 21005 20859
rect 21039 20856 21051 20859
rect 21082 20856 21088 20868
rect 21039 20828 21088 20856
rect 21039 20825 21051 20828
rect 20993 20819 21051 20825
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 17145 20791 17203 20797
rect 17145 20788 17157 20791
rect 16868 20760 17157 20788
rect 17145 20757 17157 20760
rect 17191 20757 17203 20791
rect 17145 20751 17203 20757
rect 17313 20791 17371 20797
rect 17313 20757 17325 20791
rect 17359 20788 17371 20791
rect 17678 20788 17684 20800
rect 17359 20760 17684 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 19058 20748 19064 20800
rect 19116 20788 19122 20800
rect 19337 20791 19395 20797
rect 19337 20788 19349 20791
rect 19116 20760 19349 20788
rect 19116 20748 19122 20760
rect 19337 20757 19349 20760
rect 19383 20757 19395 20791
rect 19337 20751 19395 20757
rect 19978 20748 19984 20800
rect 20036 20748 20042 20800
rect 20070 20748 20076 20800
rect 20128 20788 20134 20800
rect 20549 20791 20607 20797
rect 20549 20788 20561 20791
rect 20128 20760 20561 20788
rect 20128 20748 20134 20760
rect 20549 20757 20561 20760
rect 20595 20757 20607 20791
rect 20549 20751 20607 20757
rect 20717 20791 20775 20797
rect 20717 20757 20729 20791
rect 20763 20788 20775 20791
rect 21174 20788 21180 20800
rect 20763 20760 21180 20788
rect 20763 20757 20775 20760
rect 20717 20751 20775 20757
rect 21174 20748 21180 20760
rect 21232 20748 21238 20800
rect 22204 20788 22232 20964
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 22830 20992 22836 21004
rect 22336 20964 22836 20992
rect 22336 20952 22342 20964
rect 22830 20952 22836 20964
rect 22888 20952 22894 21004
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 22922 20924 22928 20936
rect 22612 20896 22928 20924
rect 22612 20884 22618 20896
rect 22922 20884 22928 20896
rect 22980 20884 22986 20936
rect 23106 20816 23112 20868
rect 23164 20856 23170 20868
rect 23201 20859 23259 20865
rect 23201 20856 23213 20859
rect 23164 20828 23213 20856
rect 23164 20816 23170 20828
rect 23201 20825 23213 20828
rect 23247 20825 23259 20859
rect 23492 20856 23520 21032
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 23676 20924 23704 21088
rect 24964 21069 24992 21100
rect 24949 21063 25007 21069
rect 24949 21029 24961 21063
rect 24995 21029 25007 21063
rect 24949 21023 25007 21029
rect 24486 20952 24492 21004
rect 24544 20992 24550 21004
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 24544 20964 24593 20992
rect 24544 20952 24550 20964
rect 24581 20961 24593 20964
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 23615 20896 23704 20924
rect 25056 20924 25084 20955
rect 25225 20927 25283 20933
rect 25225 20924 25237 20927
rect 25056 20896 25237 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 25225 20893 25237 20896
rect 25271 20893 25283 20927
rect 25225 20887 25283 20893
rect 23492 20828 23888 20856
rect 23201 20819 23259 20825
rect 23014 20797 23020 20800
rect 22991 20791 23020 20797
rect 22991 20788 23003 20791
rect 22204 20760 23003 20788
rect 22991 20757 23003 20760
rect 22991 20751 23020 20757
rect 23014 20748 23020 20751
rect 23072 20748 23078 20800
rect 23750 20748 23756 20800
rect 23808 20748 23814 20800
rect 23860 20788 23888 20828
rect 25130 20788 25136 20800
rect 23860 20760 25136 20788
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 25409 20791 25467 20797
rect 25409 20757 25421 20791
rect 25455 20788 25467 20791
rect 26234 20788 26240 20800
rect 25455 20760 26240 20788
rect 25455 20757 25467 20760
rect 25409 20751 25467 20757
rect 26234 20748 26240 20760
rect 26292 20748 26298 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 3142 20544 3148 20596
rect 3200 20584 3206 20596
rect 3237 20587 3295 20593
rect 3237 20584 3249 20587
rect 3200 20556 3249 20584
rect 3200 20544 3206 20556
rect 3237 20553 3249 20556
rect 3283 20553 3295 20587
rect 3237 20547 3295 20553
rect 3602 20544 3608 20596
rect 3660 20584 3666 20596
rect 3881 20587 3939 20593
rect 3881 20584 3893 20587
rect 3660 20556 3893 20584
rect 3660 20544 3666 20556
rect 3881 20553 3893 20556
rect 3927 20553 3939 20587
rect 3881 20547 3939 20553
rect 4338 20544 4344 20596
rect 4396 20544 4402 20596
rect 4982 20584 4988 20596
rect 4908 20556 4988 20584
rect 2976 20488 3648 20516
rect 2976 20389 3004 20488
rect 3421 20451 3479 20457
rect 3421 20448 3433 20451
rect 3160 20420 3433 20448
rect 3160 20392 3188 20420
rect 3421 20417 3433 20420
rect 3467 20448 3479 20451
rect 3513 20451 3571 20457
rect 3513 20448 3525 20451
rect 3467 20420 3525 20448
rect 3467 20417 3479 20420
rect 3421 20411 3479 20417
rect 3513 20417 3525 20420
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20349 3019 20383
rect 2961 20343 3019 20349
rect 2884 20244 2912 20343
rect 3142 20340 3148 20392
rect 3200 20340 3206 20392
rect 3234 20340 3240 20392
rect 3292 20340 3298 20392
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3620 20389 3648 20488
rect 4154 20476 4160 20528
rect 4212 20476 4218 20528
rect 4356 20516 4384 20544
rect 4908 20516 4936 20556
rect 4982 20544 4988 20556
rect 5040 20544 5046 20596
rect 5166 20544 5172 20596
rect 5224 20544 5230 20596
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 7098 20584 7104 20596
rect 6144 20556 7104 20584
rect 6144 20544 6150 20556
rect 7098 20544 7104 20556
rect 7156 20584 7162 20596
rect 7653 20587 7711 20593
rect 7653 20584 7665 20587
rect 7156 20556 7665 20584
rect 7156 20544 7162 20556
rect 7653 20553 7665 20556
rect 7699 20553 7711 20587
rect 7653 20547 7711 20553
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11238 20584 11244 20596
rect 11011 20556 11244 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 13262 20584 13268 20596
rect 12452 20556 13268 20584
rect 6178 20516 6184 20528
rect 4356 20488 4476 20516
rect 4172 20448 4200 20476
rect 4249 20451 4307 20457
rect 4249 20448 4261 20451
rect 4172 20420 4261 20448
rect 4249 20417 4261 20420
rect 4295 20417 4307 20451
rect 4249 20411 4307 20417
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3384 20352 3617 20380
rect 3384 20340 3390 20352
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 4356 20380 4384 20411
rect 3605 20343 3663 20349
rect 4172 20352 4384 20380
rect 4448 20380 4476 20488
rect 4540 20488 4936 20516
rect 5276 20488 6184 20516
rect 4540 20457 4568 20488
rect 5276 20460 5304 20488
rect 6178 20476 6184 20488
rect 6236 20476 6242 20528
rect 6822 20516 6828 20528
rect 6288 20488 6828 20516
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 4617 20451 4675 20457
rect 4617 20417 4629 20451
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 4632 20380 4660 20411
rect 4706 20408 4712 20460
rect 4764 20408 4770 20460
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 4985 20451 5043 20457
rect 4985 20417 4997 20451
rect 5031 20448 5043 20451
rect 5031 20420 5120 20448
rect 5031 20417 5043 20420
rect 4985 20411 5043 20417
rect 4890 20380 4896 20392
rect 4448 20352 4896 20380
rect 3252 20312 3280 20340
rect 3252 20284 3648 20312
rect 3620 20256 3648 20284
rect 3234 20244 3240 20256
rect 2884 20216 3240 20244
rect 3234 20204 3240 20216
rect 3292 20244 3298 20256
rect 3513 20247 3571 20253
rect 3513 20244 3525 20247
rect 3292 20216 3525 20244
rect 3292 20204 3298 20216
rect 3513 20213 3525 20216
rect 3559 20213 3571 20247
rect 3513 20207 3571 20213
rect 3602 20204 3608 20256
rect 3660 20204 3666 20256
rect 4062 20204 4068 20256
rect 4120 20204 4126 20256
rect 4172 20244 4200 20352
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 4246 20272 4252 20324
rect 4304 20312 4310 20324
rect 5092 20312 5120 20420
rect 5258 20408 5264 20460
rect 5316 20408 5322 20460
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20448 6055 20451
rect 6288 20448 6316 20488
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 7834 20476 7840 20528
rect 7892 20516 7898 20528
rect 12452 20525 12480 20556
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 16317 20587 16375 20593
rect 16317 20584 16329 20587
rect 15212 20556 16329 20584
rect 15212 20528 15240 20556
rect 16317 20553 16329 20556
rect 16363 20584 16375 20587
rect 16482 20584 16488 20596
rect 16363 20556 16488 20584
rect 16363 20553 16375 20556
rect 16317 20547 16375 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18969 20587 19027 20593
rect 18012 20556 18920 20584
rect 18012 20544 18018 20556
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 7892 20488 12449 20516
rect 7892 20476 7898 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12437 20479 12495 20485
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 13081 20519 13139 20525
rect 13081 20516 13093 20519
rect 13044 20488 13093 20516
rect 13044 20476 13050 20488
rect 13081 20485 13093 20488
rect 13127 20485 13139 20519
rect 13081 20479 13139 20485
rect 13188 20488 13860 20516
rect 13188 20460 13216 20488
rect 6043 20420 6316 20448
rect 6043 20417 6055 20420
rect 5997 20411 6055 20417
rect 5920 20380 5948 20411
rect 6362 20408 6368 20460
rect 6420 20408 6426 20460
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 7374 20448 7380 20460
rect 6788 20420 7380 20448
rect 6788 20408 6794 20420
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7466 20408 7472 20460
rect 7524 20448 7530 20460
rect 8205 20451 8263 20457
rect 8205 20448 8217 20451
rect 7524 20420 8217 20448
rect 7524 20408 7530 20420
rect 8205 20417 8217 20420
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20448 8447 20451
rect 9398 20448 9404 20460
rect 8435 20420 9404 20448
rect 8435 20417 8447 20420
rect 8389 20411 8447 20417
rect 6178 20380 6184 20392
rect 5920 20352 6184 20380
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 4304 20284 5120 20312
rect 6564 20312 6592 20408
rect 8220 20380 8248 20411
rect 8478 20380 8484 20392
rect 8220 20352 8484 20380
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 8205 20315 8263 20321
rect 8205 20312 8217 20315
rect 6564 20284 8217 20312
rect 4304 20272 4310 20284
rect 8205 20281 8217 20284
rect 8251 20281 8263 20315
rect 8205 20275 8263 20281
rect 9232 20256 9260 20420
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 10870 20408 10876 20460
rect 10928 20408 10934 20460
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 12406 20420 12541 20448
rect 9766 20272 9772 20324
rect 9824 20312 9830 20324
rect 12406 20312 12434 20420
rect 12529 20417 12541 20420
rect 12575 20417 12587 20451
rect 12529 20411 12587 20417
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 13170 20448 13176 20460
rect 12667 20420 13176 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 13262 20408 13268 20460
rect 13320 20408 13326 20460
rect 13832 20457 13860 20488
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 14700 20488 14964 20516
rect 14700 20476 14706 20488
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13446 20380 13452 20392
rect 13035 20352 13452 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13556 20312 13584 20411
rect 13998 20408 14004 20460
rect 14056 20408 14062 20460
rect 14090 20408 14096 20460
rect 14148 20448 14154 20460
rect 14734 20448 14740 20460
rect 14148 20420 14740 20448
rect 14148 20408 14154 20420
rect 14734 20408 14740 20420
rect 14792 20448 14798 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14792 20420 14841 20448
rect 14792 20408 14798 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 14936 20448 14964 20488
rect 15194 20476 15200 20528
rect 15252 20476 15258 20528
rect 15565 20519 15623 20525
rect 15565 20485 15577 20519
rect 15611 20516 15623 20519
rect 16117 20519 16175 20525
rect 15611 20488 16068 20516
rect 15611 20485 15623 20488
rect 15565 20479 15623 20485
rect 15654 20448 15660 20460
rect 14936 20420 15660 20448
rect 14829 20411 14887 20417
rect 15654 20408 15660 20420
rect 15712 20448 15718 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15712 20420 15761 20448
rect 15712 20408 15718 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 16040 20448 16068 20488
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 16206 20516 16212 20528
rect 16163 20488 16212 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 18138 20476 18144 20528
rect 18196 20516 18202 20528
rect 18601 20519 18659 20525
rect 18601 20516 18613 20519
rect 18196 20488 18613 20516
rect 18196 20476 18202 20488
rect 18601 20485 18613 20488
rect 18647 20485 18659 20519
rect 18801 20519 18859 20525
rect 18801 20516 18813 20519
rect 18601 20479 18659 20485
rect 18708 20488 18813 20516
rect 18708 20460 18736 20488
rect 18801 20485 18813 20488
rect 18847 20485 18859 20519
rect 18892 20516 18920 20556
rect 18969 20553 18981 20587
rect 19015 20584 19027 20587
rect 19334 20584 19340 20596
rect 19015 20556 19340 20584
rect 19015 20553 19027 20556
rect 18969 20547 19027 20553
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 23385 20587 23443 20593
rect 23385 20584 23397 20587
rect 22204 20556 23397 20584
rect 22094 20516 22100 20528
rect 18892 20488 22100 20516
rect 18801 20479 18859 20485
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 16040 20420 17172 20448
rect 15749 20411 15807 20417
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 15562 20380 15568 20392
rect 13688 20352 15568 20380
rect 13688 20340 13694 20352
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 13814 20312 13820 20324
rect 9824 20284 13820 20312
rect 9824 20272 9830 20284
rect 13814 20272 13820 20284
rect 13872 20272 13878 20324
rect 14274 20272 14280 20324
rect 14332 20272 14338 20324
rect 17144 20256 17172 20420
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 17862 20448 17868 20460
rect 17543 20420 17868 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20349 20451 20407 20457
rect 20349 20448 20361 20451
rect 20036 20420 20361 20448
rect 20036 20408 20042 20420
rect 20349 20417 20361 20420
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 20772 20420 21833 20448
rect 20772 20408 20778 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21994 20451 22052 20457
rect 21994 20448 22006 20451
rect 21821 20411 21879 20417
rect 21928 20420 22006 20448
rect 17310 20340 17316 20392
rect 17368 20340 17374 20392
rect 21928 20380 21956 20420
rect 21994 20417 22006 20420
rect 22040 20448 22052 20451
rect 22204 20448 22232 20556
rect 23385 20553 23397 20556
rect 23431 20553 23443 20587
rect 23385 20547 23443 20553
rect 26326 20544 26332 20596
rect 26384 20584 26390 20596
rect 26384 20556 26740 20584
rect 26384 20544 26390 20556
rect 23750 20476 23756 20528
rect 23808 20516 23814 20528
rect 24498 20519 24556 20525
rect 24498 20516 24510 20519
rect 23808 20488 24510 20516
rect 23808 20476 23814 20488
rect 24498 20485 24510 20488
rect 24544 20485 24556 20519
rect 24498 20479 24556 20485
rect 26234 20476 26240 20528
rect 26292 20516 26298 20528
rect 26430 20519 26488 20525
rect 26430 20516 26442 20519
rect 26292 20488 26442 20516
rect 26292 20476 26298 20488
rect 26430 20485 26442 20488
rect 26476 20485 26488 20519
rect 26430 20479 26488 20485
rect 22040 20420 22232 20448
rect 22040 20417 22052 20420
rect 21994 20411 22052 20417
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 22336 20420 22385 20448
rect 22336 20408 22342 20420
rect 22373 20417 22385 20420
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 22554 20408 22560 20460
rect 22612 20408 22618 20460
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 18800 20352 21956 20380
rect 22189 20383 22247 20389
rect 6086 20244 6092 20256
rect 4172 20216 6092 20244
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 6181 20247 6239 20253
rect 6181 20213 6193 20247
rect 6227 20244 6239 20247
rect 7650 20244 7656 20256
rect 6227 20216 7656 20244
rect 6227 20213 6239 20216
rect 6181 20207 6239 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 9214 20204 9220 20256
rect 9272 20244 9278 20256
rect 10962 20244 10968 20256
rect 9272 20216 10968 20244
rect 9272 20204 9278 20216
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 14918 20204 14924 20256
rect 14976 20204 14982 20256
rect 15378 20204 15384 20256
rect 15436 20204 15442 20256
rect 16298 20204 16304 20256
rect 16356 20204 16362 20256
rect 16482 20204 16488 20256
rect 16540 20204 16546 20256
rect 17034 20204 17040 20256
rect 17092 20204 17098 20256
rect 17126 20204 17132 20256
rect 17184 20204 17190 20256
rect 17402 20204 17408 20256
rect 17460 20204 17466 20256
rect 18800 20253 18828 20352
rect 22189 20349 22201 20383
rect 22235 20380 22247 20383
rect 22664 20380 22692 20411
rect 22922 20408 22928 20460
rect 22980 20448 22986 20460
rect 24765 20451 24823 20457
rect 24765 20448 24777 20451
rect 22980 20420 24777 20448
rect 22980 20408 22986 20420
rect 24765 20417 24777 20420
rect 24811 20448 24823 20451
rect 24946 20448 24952 20460
rect 24811 20420 24952 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 26712 20457 26740 20556
rect 26697 20451 26755 20457
rect 26697 20417 26709 20451
rect 26743 20417 26755 20451
rect 26697 20411 26755 20417
rect 22235 20352 22692 20380
rect 22235 20349 22247 20352
rect 22189 20343 22247 20349
rect 19150 20272 19156 20324
rect 19208 20312 19214 20324
rect 25317 20315 25375 20321
rect 19208 20284 23704 20312
rect 19208 20272 19214 20284
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20213 18843 20247
rect 18785 20207 18843 20213
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 20070 20244 20076 20256
rect 19024 20216 20076 20244
rect 19024 20204 19030 20216
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20533 20247 20591 20253
rect 20533 20213 20545 20247
rect 20579 20244 20591 20247
rect 20622 20244 20628 20256
rect 20579 20216 20628 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22738 20244 22744 20256
rect 22152 20216 22744 20244
rect 22152 20204 22158 20216
rect 22738 20204 22744 20216
rect 22796 20204 22802 20256
rect 22833 20247 22891 20253
rect 22833 20213 22845 20247
rect 22879 20244 22891 20247
rect 22922 20244 22928 20256
rect 22879 20216 22928 20244
rect 22879 20213 22891 20216
rect 22833 20207 22891 20213
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 23676 20244 23704 20284
rect 25317 20281 25329 20315
rect 25363 20281 25375 20315
rect 25317 20275 25375 20281
rect 25332 20244 25360 20275
rect 23676 20216 25360 20244
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 2590 20000 2596 20052
rect 2648 20000 2654 20052
rect 2682 20000 2688 20052
rect 2740 20040 2746 20052
rect 3053 20043 3111 20049
rect 3053 20040 3065 20043
rect 2740 20012 3065 20040
rect 2740 20000 2746 20012
rect 3053 20009 3065 20012
rect 3099 20040 3111 20043
rect 3142 20040 3148 20052
rect 3099 20012 3148 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3476 20012 3985 20040
rect 3476 20000 3482 20012
rect 3973 20009 3985 20012
rect 4019 20009 4031 20043
rect 3973 20003 4031 20009
rect 4709 20043 4767 20049
rect 4709 20009 4721 20043
rect 4755 20040 4767 20043
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 4755 20012 5365 20040
rect 4755 20009 4767 20012
rect 4709 20003 4767 20009
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7650 20040 7656 20052
rect 6972 20012 7656 20040
rect 6972 20000 6978 20012
rect 7650 20000 7656 20012
rect 7708 20040 7714 20052
rect 8386 20040 8392 20052
rect 7708 20012 8392 20040
rect 7708 20000 7714 20012
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 8754 20000 8760 20052
rect 8812 20000 8818 20052
rect 8941 20043 8999 20049
rect 8941 20009 8953 20043
rect 8987 20040 8999 20043
rect 9030 20040 9036 20052
rect 8987 20012 9036 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 9858 20000 9864 20052
rect 9916 20040 9922 20052
rect 9953 20043 10011 20049
rect 9953 20040 9965 20043
rect 9916 20012 9965 20040
rect 9916 20000 9922 20012
rect 9953 20009 9965 20012
rect 9999 20009 10011 20043
rect 9953 20003 10011 20009
rect 10318 20000 10324 20052
rect 10376 20040 10382 20052
rect 10870 20040 10876 20052
rect 10376 20012 10876 20040
rect 10376 20000 10382 20012
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 11517 20043 11575 20049
rect 11517 20009 11529 20043
rect 11563 20040 11575 20043
rect 11698 20040 11704 20052
rect 11563 20012 11704 20040
rect 11563 20009 11575 20012
rect 11517 20003 11575 20009
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 14090 20000 14096 20052
rect 14148 20000 14154 20052
rect 15378 20040 15384 20052
rect 14752 20012 15384 20040
rect 2608 19972 2636 20000
rect 2958 19972 2964 19984
rect 2240 19944 2964 19972
rect 2240 19845 2268 19944
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 3234 19932 3240 19984
rect 3292 19972 3298 19984
rect 3878 19972 3884 19984
rect 3292 19944 3884 19972
rect 3292 19932 3298 19944
rect 3878 19932 3884 19944
rect 3936 19932 3942 19984
rect 4985 19975 5043 19981
rect 4985 19972 4997 19975
rect 4908 19944 4997 19972
rect 2314 19864 2320 19916
rect 2372 19904 2378 19916
rect 2869 19907 2927 19913
rect 2869 19904 2881 19907
rect 2372 19876 2881 19904
rect 2372 19864 2378 19876
rect 2869 19873 2881 19876
rect 2915 19873 2927 19907
rect 4062 19904 4068 19916
rect 2869 19867 2927 19873
rect 3160 19893 3740 19904
rect 3804 19893 4068 19904
rect 3160 19876 4068 19893
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19805 2007 19839
rect 1949 19799 2007 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19836 2467 19839
rect 2498 19836 2504 19848
rect 2455 19808 2504 19836
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 750 19728 756 19780
rect 808 19768 814 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 808 19740 1501 19768
rect 808 19728 814 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 1489 19731 1547 19737
rect 1964 19700 1992 19799
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 3160 19836 3188 19876
rect 3712 19865 3832 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4908 19913 4936 19944
rect 4985 19941 4997 19944
rect 5031 19941 5043 19975
rect 4985 19935 5043 19941
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 5684 19944 5948 19972
rect 5684 19932 5690 19944
rect 4893 19907 4951 19913
rect 4893 19873 4905 19907
rect 4939 19873 4951 19907
rect 4893 19867 4951 19873
rect 5000 19876 5304 19904
rect 2823 19808 3188 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 3234 19796 3240 19848
rect 3292 19796 3298 19848
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 3605 19839 3663 19845
rect 3605 19836 3617 19839
rect 3476 19808 3617 19836
rect 3476 19796 3482 19808
rect 3605 19805 3617 19808
rect 3651 19805 3663 19839
rect 3605 19799 3663 19805
rect 3620 19768 3648 19799
rect 3878 19796 3884 19848
rect 3936 19796 3942 19848
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 3988 19768 4016 19799
rect 4338 19796 4344 19848
rect 4396 19796 4402 19848
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 5000 19836 5028 19876
rect 5276 19848 5304 19876
rect 5810 19864 5816 19916
rect 5868 19864 5874 19916
rect 5920 19913 5948 19944
rect 5994 19932 6000 19984
rect 6052 19972 6058 19984
rect 6178 19972 6184 19984
rect 6052 19944 6184 19972
rect 6052 19932 6058 19944
rect 6178 19932 6184 19944
rect 6236 19972 6242 19984
rect 8294 19972 8300 19984
rect 6236 19944 8300 19972
rect 6236 19932 6242 19944
rect 8294 19932 8300 19944
rect 8352 19972 8358 19984
rect 11072 19972 11100 20000
rect 8352 19944 8616 19972
rect 8352 19932 8358 19944
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 8478 19864 8484 19916
rect 8536 19864 8542 19916
rect 4663 19808 5028 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 5132 19808 5181 19836
rect 5132 19796 5138 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 5258 19796 5264 19848
rect 5316 19796 5322 19848
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 7800 19808 8217 19836
rect 7800 19796 7806 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8496 19836 8524 19864
rect 8588 19845 8616 19944
rect 10244 19944 11100 19972
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 10244 19913 10272 19944
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 9272 19876 9505 19904
rect 9272 19864 9278 19876
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 10229 19907 10287 19913
rect 10229 19873 10241 19907
rect 10275 19873 10287 19907
rect 10229 19867 10287 19873
rect 10318 19864 10324 19916
rect 10376 19904 10382 19916
rect 10781 19907 10839 19913
rect 10781 19904 10793 19907
rect 10376 19876 10793 19904
rect 10376 19864 10382 19876
rect 10781 19873 10793 19876
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 11072 19904 11100 19944
rect 11149 19907 11207 19913
rect 11149 19904 11161 19907
rect 11072 19876 11161 19904
rect 11149 19873 11161 19876
rect 11195 19873 11207 19907
rect 14090 19904 14096 19916
rect 11149 19867 11207 19873
rect 13004 19876 14096 19904
rect 13004 19848 13032 19876
rect 14090 19864 14096 19876
rect 14148 19904 14154 19916
rect 14461 19907 14519 19913
rect 14461 19904 14473 19907
rect 14148 19876 14473 19904
rect 14148 19864 14154 19876
rect 14461 19873 14473 19876
rect 14507 19873 14519 19907
rect 14461 19867 14519 19873
rect 8343 19808 8524 19836
rect 8573 19839 8631 19845
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 9858 19796 9864 19848
rect 9916 19796 9922 19848
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19836 10011 19839
rect 9999 19808 10364 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 3620 19740 4016 19768
rect 4706 19728 4712 19780
rect 4764 19768 4770 19780
rect 4985 19771 5043 19777
rect 4985 19768 4997 19771
rect 4764 19740 4997 19768
rect 4764 19728 4770 19740
rect 4985 19737 4997 19740
rect 5031 19768 5043 19771
rect 5902 19768 5908 19780
rect 5031 19740 5908 19768
rect 5031 19737 5043 19740
rect 4985 19731 5043 19737
rect 5902 19728 5908 19740
rect 5960 19728 5966 19780
rect 9309 19771 9367 19777
rect 9309 19768 9321 19771
rect 6104 19740 9321 19768
rect 6104 19712 6132 19740
rect 9309 19737 9321 19740
rect 9355 19768 9367 19771
rect 9766 19768 9772 19780
rect 9355 19740 9772 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9766 19728 9772 19740
rect 9824 19728 9830 19780
rect 10336 19768 10364 19808
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11330 19846 11336 19848
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10652 19808 10701 19836
rect 10652 19796 10658 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 11256 19818 11336 19846
rect 11256 19768 11284 19818
rect 11330 19796 11336 19818
rect 11388 19796 11394 19848
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14182 19836 14188 19848
rect 13872 19808 14188 19836
rect 13872 19796 13878 19808
rect 14182 19796 14188 19808
rect 14240 19836 14246 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14240 19808 14289 19836
rect 14240 19796 14246 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19836 14611 19839
rect 14642 19836 14648 19848
rect 14599 19808 14648 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 10336 19740 11284 19768
rect 13280 19768 13308 19796
rect 13722 19768 13728 19780
rect 13280 19740 13728 19768
rect 13722 19728 13728 19740
rect 13780 19768 13786 19780
rect 14384 19768 14412 19799
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 14752 19845 14780 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 16758 20000 16764 20052
rect 16816 20000 16822 20052
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17310 20040 17316 20052
rect 17175 20012 17316 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17310 20000 17316 20012
rect 17368 20000 17374 20052
rect 17954 20000 17960 20052
rect 18012 20000 18018 20052
rect 18601 20043 18659 20049
rect 18601 20009 18613 20043
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 16776 19972 16804 20000
rect 17405 19975 17463 19981
rect 17405 19972 17417 19975
rect 16776 19944 17417 19972
rect 17405 19941 17417 19944
rect 17451 19941 17463 19975
rect 17405 19935 17463 19941
rect 17589 19975 17647 19981
rect 17589 19941 17601 19975
rect 17635 19972 17647 19975
rect 18417 19975 18475 19981
rect 18417 19972 18429 19975
rect 17635 19944 18429 19972
rect 17635 19941 17647 19944
rect 17589 19935 17647 19941
rect 18417 19941 18429 19944
rect 18463 19941 18475 19975
rect 18616 19972 18644 20003
rect 18782 20000 18788 20052
rect 18840 20040 18846 20052
rect 19242 20040 19248 20052
rect 18840 20012 19248 20040
rect 18840 20000 18846 20012
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20257 20043 20315 20049
rect 20257 20040 20269 20043
rect 20036 20012 20269 20040
rect 20036 20000 20042 20012
rect 20257 20009 20269 20012
rect 20303 20009 20315 20043
rect 20990 20040 20996 20052
rect 20257 20003 20315 20009
rect 20364 20012 20996 20040
rect 18966 19972 18972 19984
rect 18616 19944 18972 19972
rect 18417 19935 18475 19941
rect 18966 19932 18972 19944
rect 19024 19972 19030 19984
rect 20364 19972 20392 20012
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 21358 20000 21364 20052
rect 21416 20040 21422 20052
rect 21729 20043 21787 20049
rect 21729 20040 21741 20043
rect 21416 20012 21741 20040
rect 21416 20000 21422 20012
rect 21729 20009 21741 20012
rect 21775 20009 21787 20043
rect 21729 20003 21787 20009
rect 22278 20000 22284 20052
rect 22336 20000 22342 20052
rect 22554 20000 22560 20052
rect 22612 20040 22618 20052
rect 22612 20012 23244 20040
rect 22612 20000 22618 20012
rect 22296 19972 22324 20000
rect 19024 19944 20392 19972
rect 21376 19944 22324 19972
rect 19024 19932 19030 19944
rect 17126 19864 17132 19916
rect 17184 19904 17190 19916
rect 19150 19904 19156 19916
rect 17184 19876 19156 19904
rect 17184 19864 17190 19876
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19805 14795 19839
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 14737 19799 14795 19805
rect 14844 19808 15025 19836
rect 14844 19768 14872 19808
rect 15013 19805 15025 19808
rect 15059 19805 15071 19839
rect 15013 19799 15071 19805
rect 17494 19796 17500 19848
rect 17552 19796 17558 19848
rect 17696 19845 17724 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 19944 19876 20392 19904
rect 19944 19864 19950 19876
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 17681 19799 17739 19805
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19836 17923 19839
rect 17954 19836 17960 19848
rect 17911 19808 17960 19836
rect 17911 19805 17923 19808
rect 17865 19799 17923 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 15258 19771 15316 19777
rect 15258 19768 15270 19771
rect 13780 19740 14412 19768
rect 14568 19740 14872 19768
rect 14936 19740 15270 19768
rect 13780 19728 13786 19740
rect 14568 19712 14596 19740
rect 2222 19700 2228 19712
rect 1964 19672 2228 19700
rect 2222 19660 2228 19672
rect 2280 19700 2286 19712
rect 2406 19700 2412 19712
rect 2280 19672 2412 19700
rect 2280 19660 2286 19672
rect 2406 19660 2412 19672
rect 2464 19660 2470 19712
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 3142 19700 3148 19712
rect 2924 19672 3148 19700
rect 2924 19660 2930 19672
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 4798 19700 4804 19712
rect 3467 19672 4804 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 4890 19660 4896 19712
rect 4948 19660 4954 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 5721 19703 5779 19709
rect 5721 19700 5733 19703
rect 5592 19672 5733 19700
rect 5592 19660 5598 19672
rect 5721 19669 5733 19672
rect 5767 19700 5779 19703
rect 5810 19700 5816 19712
rect 5767 19672 5816 19700
rect 5767 19669 5779 19672
rect 5721 19663 5779 19669
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 6086 19660 6092 19712
rect 6144 19660 6150 19712
rect 6914 19660 6920 19712
rect 6972 19660 6978 19712
rect 8386 19660 8392 19712
rect 8444 19660 8450 19712
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 9858 19700 9864 19712
rect 9447 19672 9864 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 10045 19703 10103 19709
rect 10045 19669 10057 19703
rect 10091 19700 10103 19703
rect 10134 19700 10140 19712
rect 10091 19672 10140 19700
rect 10091 19669 10103 19672
rect 10045 19663 10103 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 14550 19660 14556 19712
rect 14608 19660 14614 19712
rect 14936 19709 14964 19740
rect 15258 19737 15270 19740
rect 15304 19737 15316 19771
rect 15258 19731 15316 19737
rect 15562 19728 15568 19780
rect 15620 19768 15626 19780
rect 16022 19768 16028 19780
rect 15620 19740 16028 19768
rect 15620 19728 15626 19740
rect 16022 19728 16028 19740
rect 16080 19768 16086 19780
rect 18156 19768 18184 19799
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 18690 19836 18696 19848
rect 18564 19808 18696 19836
rect 18564 19796 18570 19808
rect 18690 19796 18696 19808
rect 18748 19836 18754 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18748 19808 19257 19836
rect 18748 19796 18754 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20364 19845 20392 19876
rect 20349 19839 20407 19845
rect 19392 19808 20116 19836
rect 19392 19796 19398 19808
rect 16080 19740 18184 19768
rect 18248 19768 18276 19796
rect 18785 19771 18843 19777
rect 18785 19768 18797 19771
rect 18248 19740 18797 19768
rect 16080 19728 16086 19740
rect 18785 19737 18797 19740
rect 18831 19768 18843 19771
rect 19058 19768 19064 19780
rect 18831 19740 19064 19768
rect 18831 19737 18843 19740
rect 18785 19731 18843 19737
rect 19058 19728 19064 19740
rect 19116 19728 19122 19780
rect 19889 19771 19947 19777
rect 19889 19737 19901 19771
rect 19935 19768 19947 19771
rect 19978 19768 19984 19780
rect 19935 19740 19984 19768
rect 19935 19737 19947 19740
rect 19889 19731 19947 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 20088 19777 20116 19808
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 21376 19836 21404 19944
rect 23216 19913 23244 20012
rect 23201 19907 23259 19913
rect 23201 19873 23213 19907
rect 23247 19873 23259 19907
rect 23201 19867 23259 19873
rect 20395 19808 21404 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 22922 19796 22928 19848
rect 22980 19845 22986 19848
rect 22980 19836 22992 19845
rect 22980 19808 23025 19836
rect 22980 19799 22992 19808
rect 22980 19796 22986 19799
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 24946 19796 24952 19848
rect 25004 19836 25010 19848
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25004 19808 25789 19836
rect 25004 19796 25010 19808
rect 25777 19805 25789 19808
rect 25823 19836 25835 19839
rect 25958 19836 25964 19848
rect 25823 19808 25964 19836
rect 25823 19805 25835 19808
rect 25777 19799 25835 19805
rect 25958 19796 25964 19808
rect 26016 19836 26022 19848
rect 26326 19836 26332 19848
rect 26016 19808 26332 19836
rect 26016 19796 26022 19808
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 20622 19777 20628 19780
rect 20073 19771 20131 19777
rect 20073 19737 20085 19771
rect 20119 19768 20131 19771
rect 20119 19740 20576 19768
rect 20119 19737 20131 19740
rect 20073 19731 20131 19737
rect 14921 19703 14979 19709
rect 14921 19669 14933 19703
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 16114 19660 16120 19712
rect 16172 19700 16178 19712
rect 16393 19703 16451 19709
rect 16393 19700 16405 19703
rect 16172 19672 16405 19700
rect 16172 19660 16178 19672
rect 16393 19669 16405 19672
rect 16439 19669 16451 19703
rect 16393 19663 16451 19669
rect 17310 19660 17316 19712
rect 17368 19700 17374 19712
rect 17770 19700 17776 19712
rect 17368 19672 17776 19700
rect 17368 19660 17374 19672
rect 17770 19660 17776 19672
rect 17828 19660 17834 19712
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 18575 19703 18633 19709
rect 18575 19700 18587 19703
rect 18380 19672 18587 19700
rect 18380 19660 18386 19672
rect 18575 19669 18587 19672
rect 18621 19669 18633 19703
rect 18575 19663 18633 19669
rect 19242 19660 19248 19712
rect 19300 19700 19306 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 19300 19672 19441 19700
rect 19300 19660 19306 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 20548 19700 20576 19740
rect 20616 19731 20628 19777
rect 20680 19768 20686 19780
rect 20680 19740 20716 19768
rect 20622 19728 20628 19731
rect 20680 19728 20686 19740
rect 20990 19728 20996 19780
rect 21048 19768 21054 19780
rect 21048 19740 24440 19768
rect 21048 19728 21054 19740
rect 21821 19703 21879 19709
rect 21821 19700 21833 19703
rect 20548 19672 21833 19700
rect 19429 19663 19487 19669
rect 21821 19669 21833 19672
rect 21867 19669 21879 19703
rect 21821 19663 21879 19669
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 24412 19709 24440 19740
rect 25406 19728 25412 19780
rect 25464 19768 25470 19780
rect 25510 19771 25568 19777
rect 25510 19768 25522 19771
rect 25464 19740 25522 19768
rect 25464 19728 25470 19740
rect 25510 19737 25522 19740
rect 25556 19737 25568 19771
rect 25510 19731 25568 19737
rect 24397 19703 24455 19709
rect 24397 19669 24409 19703
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 2498 19496 2504 19508
rect 2096 19468 2504 19496
rect 2096 19456 2102 19468
rect 2498 19456 2504 19468
rect 2556 19496 2562 19508
rect 4341 19499 4399 19505
rect 4341 19496 4353 19499
rect 2556 19468 4353 19496
rect 2556 19456 2562 19468
rect 4341 19465 4353 19468
rect 4387 19465 4399 19499
rect 4341 19459 4399 19465
rect 4617 19499 4675 19505
rect 4617 19465 4629 19499
rect 4663 19465 4675 19499
rect 4617 19459 4675 19465
rect 1397 19431 1455 19437
rect 1397 19397 1409 19431
rect 1443 19397 1455 19431
rect 1397 19391 1455 19397
rect 2409 19431 2467 19437
rect 2409 19397 2421 19431
rect 2455 19428 2467 19431
rect 3237 19431 3295 19437
rect 3237 19428 3249 19431
rect 2455 19400 3249 19428
rect 2455 19397 2467 19400
rect 2409 19391 2467 19397
rect 3237 19397 3249 19400
rect 3283 19397 3295 19431
rect 4632 19428 4660 19459
rect 5258 19456 5264 19508
rect 5316 19496 5322 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 5316 19468 6561 19496
rect 5316 19456 5322 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 6549 19459 6607 19465
rect 6822 19456 6828 19508
rect 6880 19496 6886 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 6880 19468 7481 19496
rect 6880 19456 6886 19468
rect 7469 19465 7481 19468
rect 7515 19465 7527 19499
rect 7469 19459 7527 19465
rect 8205 19499 8263 19505
rect 8205 19465 8217 19499
rect 8251 19496 8263 19499
rect 8386 19496 8392 19508
rect 8251 19468 8392 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 9306 19456 9312 19508
rect 9364 19456 9370 19508
rect 9674 19505 9680 19508
rect 9670 19496 9680 19505
rect 9635 19468 9680 19496
rect 9670 19459 9680 19468
rect 9674 19456 9680 19459
rect 9732 19456 9738 19508
rect 9950 19456 9956 19508
rect 10008 19456 10014 19508
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19496 10563 19499
rect 11054 19496 11060 19508
rect 10551 19468 11060 19496
rect 10551 19465 10563 19468
rect 10505 19459 10563 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11330 19456 11336 19508
rect 11388 19456 11394 19508
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 14792 19468 15700 19496
rect 14792 19456 14798 19468
rect 6730 19428 6736 19440
rect 3237 19391 3295 19397
rect 3712 19400 4660 19428
rect 4908 19400 6736 19428
rect 1412 19360 1440 19391
rect 1412 19332 2728 19360
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19261 1639 19295
rect 1581 19255 1639 19261
rect 1596 19156 1624 19255
rect 1670 19252 1676 19304
rect 1728 19252 1734 19304
rect 1762 19252 1768 19304
rect 1820 19252 1826 19304
rect 2700 19301 2728 19332
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 2869 19363 2927 19369
rect 2869 19329 2881 19363
rect 2915 19360 2927 19363
rect 3142 19360 3148 19372
rect 2915 19332 3148 19360
rect 2915 19329 2927 19332
rect 2869 19323 2927 19329
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3510 19320 3516 19372
rect 3568 19320 3574 19372
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 3712 19369 3740 19400
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 3878 19320 3884 19372
rect 3936 19320 3942 19372
rect 4154 19320 4160 19372
rect 4212 19320 4218 19372
rect 4430 19320 4436 19372
rect 4488 19320 4494 19372
rect 4908 19369 4936 19400
rect 5552 19372 5580 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 4755 19363 4813 19369
rect 4755 19360 4767 19363
rect 4540 19332 4767 19360
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2643 19264 2697 19292
rect 2685 19261 2697 19264
rect 2731 19292 2743 19295
rect 4172 19292 4200 19320
rect 4540 19292 4568 19332
rect 4755 19329 4767 19332
rect 4801 19329 4813 19363
rect 4755 19323 4813 19329
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 2731 19264 2912 19292
rect 4172 19264 4568 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 2225 19227 2283 19233
rect 2225 19193 2237 19227
rect 2271 19224 2283 19227
rect 2774 19224 2780 19236
rect 2271 19196 2780 19224
rect 2271 19193 2283 19196
rect 2225 19187 2283 19193
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 2884 19168 2912 19264
rect 4157 19227 4215 19233
rect 4157 19193 4169 19227
rect 4203 19224 4215 19227
rect 5000 19224 5028 19323
rect 5074 19320 5080 19372
rect 5132 19369 5138 19372
rect 5132 19363 5171 19369
rect 5159 19329 5171 19363
rect 5132 19323 5171 19329
rect 5261 19363 5319 19369
rect 5261 19329 5273 19363
rect 5307 19360 5319 19363
rect 5307 19332 5341 19360
rect 5307 19329 5319 19332
rect 5261 19323 5319 19329
rect 5132 19320 5138 19323
rect 5276 19292 5304 19323
rect 5534 19320 5540 19372
rect 5592 19320 5598 19372
rect 6365 19363 6423 19369
rect 5644 19332 6316 19360
rect 5184 19264 5304 19292
rect 5184 19236 5212 19264
rect 4203 19196 5028 19224
rect 4203 19193 4215 19196
rect 4157 19187 4215 19193
rect 5166 19184 5172 19236
rect 5224 19184 5230 19236
rect 5644 19224 5672 19332
rect 6288 19292 6316 19332
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 6546 19360 6552 19372
rect 6411 19332 6552 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 6840 19360 6868 19456
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 8938 19428 8944 19440
rect 7607 19400 8944 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 8938 19388 8944 19400
rect 8996 19388 9002 19440
rect 6656 19332 6868 19360
rect 7285 19363 7343 19369
rect 6656 19292 6684 19332
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 7742 19360 7748 19372
rect 7331 19332 7748 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7742 19320 7748 19332
rect 7800 19360 7806 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7800 19332 7849 19360
rect 7800 19320 7806 19332
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19360 8079 19363
rect 8205 19363 8263 19369
rect 8067 19332 8101 19360
rect 8067 19329 8079 19332
rect 8021 19323 8079 19329
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 9030 19360 9036 19372
rect 8251 19332 9036 19360
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 6288 19264 6684 19292
rect 7650 19252 7656 19304
rect 7708 19292 7714 19304
rect 8036 19292 8064 19323
rect 9030 19320 9036 19332
rect 9088 19360 9094 19372
rect 9324 19360 9352 19456
rect 10413 19431 10471 19437
rect 10413 19397 10425 19431
rect 10459 19428 10471 19431
rect 10962 19428 10968 19440
rect 10459 19400 10968 19428
rect 10459 19397 10471 19400
rect 10413 19391 10471 19397
rect 10962 19388 10968 19400
rect 11020 19388 11026 19440
rect 11072 19391 11192 19394
rect 11058 19385 11192 19391
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 14369 19431 14427 19437
rect 14369 19428 14381 19431
rect 11480 19400 14381 19428
rect 11480 19388 11486 19400
rect 14369 19397 14381 19400
rect 14415 19428 14427 19431
rect 15194 19428 15200 19440
rect 14415 19400 15200 19428
rect 14415 19397 14427 19400
rect 14369 19391 14427 19397
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 9088 19332 9352 19360
rect 9088 19320 9094 19332
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9769 19363 9827 19369
rect 9640 19332 9720 19360
rect 9640 19320 9646 19332
rect 7708 19264 8064 19292
rect 9508 19292 9536 19320
rect 9692 19292 9720 19332
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 10137 19363 10195 19369
rect 10137 19360 10149 19363
rect 9815 19332 10149 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 10137 19329 10149 19332
rect 10183 19360 10195 19363
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10183 19332 10701 19360
rect 10183 19329 10195 19332
rect 10137 19323 10195 19329
rect 10689 19329 10701 19332
rect 10735 19360 10747 19363
rect 10735 19332 11008 19360
rect 11058 19351 11070 19385
rect 11104 19366 11192 19385
rect 11104 19351 11116 19366
rect 11058 19345 11116 19351
rect 11164 19360 11192 19366
rect 11238 19360 11244 19372
rect 11164 19332 11244 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 10321 19295 10379 19301
rect 9508 19264 9628 19292
rect 9692 19264 10272 19292
rect 7708 19252 7714 19264
rect 9600 19236 9628 19264
rect 6454 19224 6460 19236
rect 5644 19196 6460 19224
rect 6454 19184 6460 19196
rect 6512 19184 6518 19236
rect 9582 19184 9588 19236
rect 9640 19184 9646 19236
rect 2682 19156 2688 19168
rect 1596 19128 2688 19156
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 2866 19116 2872 19168
rect 2924 19116 2930 19168
rect 3970 19116 3976 19168
rect 4028 19156 4034 19168
rect 4890 19156 4896 19168
rect 4028 19128 4896 19156
rect 4028 19116 4034 19128
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 7006 19116 7012 19168
rect 7064 19116 7070 19168
rect 10134 19116 10140 19168
rect 10192 19116 10198 19168
rect 10244 19156 10272 19264
rect 10321 19261 10333 19295
rect 10367 19292 10379 19295
rect 10410 19292 10416 19304
rect 10367 19264 10416 19292
rect 10367 19261 10379 19264
rect 10321 19255 10379 19261
rect 10410 19252 10416 19264
rect 10468 19292 10474 19304
rect 10873 19295 10931 19301
rect 10873 19292 10885 19295
rect 10468 19264 10885 19292
rect 10468 19252 10474 19264
rect 10873 19261 10885 19264
rect 10919 19261 10931 19295
rect 10980 19292 11008 19332
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13044 19332 13461 19360
rect 13044 19320 13050 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13449 19323 13507 19329
rect 13722 19320 13728 19372
rect 13780 19320 13786 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 13872 19332 13921 19360
rect 13872 19320 13878 19332
rect 13909 19329 13921 19332
rect 13955 19329 13967 19363
rect 13909 19323 13967 19329
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14047 19332 15240 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 10980 19264 11345 19292
rect 10873 19255 10931 19261
rect 11333 19261 11345 19264
rect 11379 19292 11391 19295
rect 12345 19295 12403 19301
rect 11379 19264 11836 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 10888 19224 10916 19255
rect 11808 19236 11836 19264
rect 12345 19261 12357 19295
rect 12391 19261 12403 19295
rect 13740 19292 13768 19320
rect 14016 19292 14044 19323
rect 13740 19264 14044 19292
rect 14461 19295 14519 19301
rect 12345 19255 12403 19261
rect 14461 19261 14473 19295
rect 14507 19292 14519 19295
rect 14642 19292 14648 19304
rect 14507 19264 14648 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 10888 19196 11284 19224
rect 11256 19168 11284 19196
rect 11790 19184 11796 19236
rect 11848 19184 11854 19236
rect 12360 19168 12388 19255
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 15028 19264 15117 19292
rect 10870 19156 10876 19168
rect 10244 19128 10876 19156
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 11020 19128 11161 19156
rect 11020 19116 11026 19128
rect 11149 19125 11161 19128
rect 11195 19125 11207 19159
rect 11149 19119 11207 19125
rect 11238 19116 11244 19168
rect 11296 19116 11302 19168
rect 12342 19116 12348 19168
rect 12400 19116 12406 19168
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 12529 19159 12587 19165
rect 12529 19125 12541 19159
rect 12575 19156 12587 19159
rect 12710 19156 12716 19168
rect 12575 19128 12716 19156
rect 12575 19125 12587 19128
rect 12529 19119 12587 19125
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14274 19156 14280 19168
rect 13412 19128 14280 19156
rect 13412 19116 13418 19128
rect 14274 19116 14280 19128
rect 14332 19156 14338 19168
rect 15028 19156 15056 19264
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15212 19292 15240 19332
rect 15470 19320 15476 19372
rect 15528 19360 15534 19372
rect 15672 19369 15700 19468
rect 17494 19456 17500 19508
rect 17552 19456 17558 19508
rect 18598 19456 18604 19508
rect 18656 19456 18662 19508
rect 18690 19456 18696 19508
rect 18748 19496 18754 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18748 19468 18981 19496
rect 18748 19456 18754 19468
rect 18969 19465 18981 19468
rect 19015 19496 19027 19499
rect 19518 19496 19524 19508
rect 19015 19468 19524 19496
rect 19015 19465 19027 19468
rect 18969 19459 19027 19465
rect 19518 19456 19524 19468
rect 19576 19496 19582 19508
rect 19889 19499 19947 19505
rect 19576 19468 19840 19496
rect 19576 19456 19582 19468
rect 16022 19388 16028 19440
rect 16080 19388 16086 19440
rect 17660 19431 17718 19437
rect 17660 19397 17672 19431
rect 17706 19428 17718 19431
rect 17770 19428 17776 19440
rect 17706 19400 17776 19428
rect 17706 19397 17718 19400
rect 17660 19391 17718 19397
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 17865 19431 17923 19437
rect 17865 19397 17877 19431
rect 17911 19428 17923 19431
rect 17954 19428 17960 19440
rect 17911 19400 17960 19428
rect 17911 19397 17923 19400
rect 17865 19391 17923 19397
rect 17954 19388 17960 19400
rect 18012 19428 18018 19440
rect 18138 19428 18144 19440
rect 18012 19400 18144 19428
rect 18012 19388 18018 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18230 19388 18236 19440
rect 18288 19388 18294 19440
rect 18449 19431 18507 19437
rect 18449 19397 18461 19431
rect 18495 19428 18507 19431
rect 19242 19428 19248 19440
rect 18495 19400 19248 19428
rect 18495 19397 18507 19400
rect 18449 19391 18507 19397
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19429 19431 19487 19437
rect 19429 19397 19441 19431
rect 19475 19428 19487 19431
rect 19610 19428 19616 19440
rect 19475 19400 19616 19428
rect 19475 19397 19487 19400
rect 19429 19391 19487 19397
rect 19610 19388 19616 19400
rect 19668 19388 19674 19440
rect 19812 19437 19840 19468
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 19978 19496 19984 19508
rect 19935 19468 19984 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 19797 19431 19855 19437
rect 19797 19397 19809 19431
rect 19843 19397 19855 19431
rect 19904 19428 19932 19459
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 23566 19456 23572 19508
rect 23624 19456 23630 19508
rect 25133 19499 25191 19505
rect 25133 19465 25145 19499
rect 25179 19465 25191 19499
rect 25133 19459 25191 19465
rect 20438 19428 20444 19440
rect 19904 19400 20444 19428
rect 19797 19391 19855 19397
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 23468 19431 23526 19437
rect 23468 19397 23480 19431
rect 23514 19428 23526 19431
rect 23584 19428 23612 19456
rect 23514 19400 23612 19428
rect 23514 19397 23526 19400
rect 23468 19391 23526 19397
rect 24486 19388 24492 19440
rect 24544 19428 24550 19440
rect 24673 19431 24731 19437
rect 24673 19428 24685 19431
rect 24544 19400 24685 19428
rect 24544 19388 24550 19400
rect 24673 19397 24685 19400
rect 24719 19397 24731 19431
rect 24673 19391 24731 19397
rect 15565 19363 15623 19369
rect 15565 19360 15577 19363
rect 15528 19332 15577 19360
rect 15528 19320 15534 19332
rect 15565 19329 15577 19332
rect 15611 19329 15623 19363
rect 15565 19323 15623 19329
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 19628 19360 19656 19388
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 15703 19332 19472 19360
rect 19628 19332 19993 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15378 19292 15384 19304
rect 15212 19264 15384 19292
rect 15105 19255 15163 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 16132 19224 16160 19255
rect 16666 19252 16672 19304
rect 16724 19292 16730 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16724 19264 16957 19292
rect 16724 19252 16730 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 16945 19255 17003 19261
rect 17236 19264 18889 19292
rect 16298 19224 16304 19236
rect 15344 19196 16304 19224
rect 15344 19184 15350 19196
rect 16298 19184 16304 19196
rect 16356 19184 16362 19236
rect 15102 19156 15108 19168
rect 14332 19128 15108 19156
rect 14332 19116 14338 19128
rect 15102 19116 15108 19128
rect 15160 19156 15166 19168
rect 17236 19156 17264 19264
rect 18877 19261 18889 19264
rect 18923 19292 18935 19295
rect 19334 19292 19340 19304
rect 18923 19264 19340 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 17313 19227 17371 19233
rect 17313 19193 17325 19227
rect 17359 19224 17371 19227
rect 18693 19227 18751 19233
rect 17359 19196 18644 19224
rect 17359 19193 17371 19196
rect 17313 19187 17371 19193
rect 15160 19128 17264 19156
rect 15160 19116 15166 19128
rect 17402 19116 17408 19168
rect 17460 19116 17466 19168
rect 17696 19165 17724 19196
rect 17681 19159 17739 19165
rect 17681 19125 17693 19159
rect 17727 19125 17739 19159
rect 17681 19119 17739 19125
rect 18417 19159 18475 19165
rect 18417 19125 18429 19159
rect 18463 19156 18475 19159
rect 18506 19156 18512 19168
rect 18463 19128 18512 19156
rect 18463 19125 18475 19128
rect 18417 19119 18475 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18616 19156 18644 19196
rect 18693 19193 18705 19227
rect 18739 19224 18751 19227
rect 18782 19224 18788 19236
rect 18739 19196 18788 19224
rect 18739 19193 18751 19196
rect 18693 19187 18751 19193
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 19444 19233 19472 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 19429 19227 19487 19233
rect 19429 19193 19441 19227
rect 19475 19224 19487 19227
rect 19886 19224 19892 19236
rect 19475 19196 19892 19224
rect 19475 19193 19487 19196
rect 19429 19187 19487 19193
rect 19886 19184 19892 19196
rect 19944 19184 19950 19236
rect 19996 19224 20024 19323
rect 20530 19320 20536 19372
rect 20588 19320 20594 19372
rect 25148 19360 25176 19459
rect 25406 19456 25412 19508
rect 25464 19456 25470 19508
rect 25225 19363 25283 19369
rect 25225 19360 25237 19363
rect 23216 19332 24256 19360
rect 25148 19332 25237 19360
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20312 19264 20361 19292
rect 20312 19252 20318 19264
rect 20349 19261 20361 19264
rect 20395 19292 20407 19295
rect 21634 19292 21640 19304
rect 20395 19264 21640 19292
rect 20395 19261 20407 19264
rect 20349 19255 20407 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 23216 19301 23244 19332
rect 23201 19295 23259 19301
rect 23201 19261 23213 19295
rect 23247 19261 23259 19295
rect 24228 19292 24256 19332
rect 25225 19329 25237 19332
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25866 19320 25872 19372
rect 25924 19360 25930 19372
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 25924 19332 26065 19360
rect 25924 19320 25930 19332
rect 26053 19329 26065 19332
rect 26099 19329 26111 19363
rect 26053 19323 26111 19329
rect 24486 19292 24492 19304
rect 24228 19264 24492 19292
rect 23201 19255 23259 19261
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 20622 19224 20628 19236
rect 19996 19196 20628 19224
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 20990 19184 20996 19236
rect 21048 19224 21054 19236
rect 21726 19224 21732 19236
rect 21048 19196 21732 19224
rect 21048 19184 21054 19196
rect 21726 19184 21732 19196
rect 21784 19184 21790 19236
rect 24949 19227 25007 19233
rect 24949 19224 24961 19227
rect 24596 19196 24961 19224
rect 24596 19168 24624 19196
rect 24949 19193 24961 19196
rect 24995 19193 25007 19227
rect 24949 19187 25007 19193
rect 23934 19156 23940 19168
rect 18616 19128 23940 19156
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 24578 19116 24584 19168
rect 24636 19116 24642 19168
rect 26234 19116 26240 19168
rect 26292 19116 26298 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 2501 18955 2559 18961
rect 1728 18924 2176 18952
rect 1728 18912 1734 18924
rect 2041 18887 2099 18893
rect 2041 18853 2053 18887
rect 2087 18853 2099 18887
rect 2041 18847 2099 18853
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18748 2007 18751
rect 2056 18748 2084 18847
rect 2148 18816 2176 18924
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2682 18952 2688 18964
rect 2547 18924 2688 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2682 18912 2688 18924
rect 2740 18912 2746 18964
rect 4246 18912 4252 18964
rect 4304 18912 4310 18964
rect 7282 18952 7288 18964
rect 6748 18924 7288 18952
rect 4154 18844 4160 18896
rect 4212 18884 4218 18896
rect 4709 18887 4767 18893
rect 4709 18884 4721 18887
rect 4212 18856 4721 18884
rect 4212 18844 4218 18856
rect 4709 18853 4721 18856
rect 4755 18853 4767 18887
rect 4709 18847 4767 18853
rect 2314 18816 2320 18828
rect 2148 18788 2320 18816
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 2685 18819 2743 18825
rect 2685 18816 2697 18819
rect 2464 18788 2697 18816
rect 2464 18776 2470 18788
rect 2685 18785 2697 18788
rect 2731 18785 2743 18819
rect 2685 18779 2743 18785
rect 3988 18788 4660 18816
rect 1995 18720 2084 18748
rect 1995 18717 2007 18720
rect 1949 18711 2007 18717
rect 2590 18708 2596 18760
rect 2648 18708 2654 18760
rect 2866 18708 2872 18760
rect 2924 18708 2930 18760
rect 3050 18708 3056 18760
rect 3108 18748 3114 18760
rect 3878 18748 3884 18760
rect 3108 18720 3884 18748
rect 3108 18708 3114 18720
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 1765 18615 1823 18621
rect 1765 18581 1777 18615
rect 1811 18612 1823 18615
rect 3068 18612 3096 18708
rect 3988 18689 4016 18788
rect 4632 18757 4660 18788
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 4172 18720 4445 18748
rect 4172 18689 4200 18720
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6236 18720 6653 18748
rect 6236 18708 6242 18720
rect 6641 18717 6653 18720
rect 6687 18748 6699 18751
rect 6748 18748 6776 18924
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 9582 18912 9588 18964
rect 9640 18952 9646 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 9640 18924 10609 18952
rect 9640 18912 9646 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 11790 18912 11796 18964
rect 11848 18912 11854 18964
rect 13354 18952 13360 18964
rect 11900 18924 13360 18952
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 11900 18884 11928 18924
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 18601 18955 18659 18961
rect 16356 18924 18552 18952
rect 16356 18912 16362 18924
rect 9364 18856 11928 18884
rect 9364 18844 9370 18856
rect 12526 18844 12532 18896
rect 12584 18844 12590 18896
rect 18524 18884 18552 18924
rect 18601 18921 18613 18955
rect 18647 18952 18659 18955
rect 19150 18952 19156 18964
rect 18647 18924 19156 18952
rect 18647 18921 18659 18924
rect 18601 18915 18659 18921
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 19242 18912 19248 18964
rect 19300 18912 19306 18964
rect 19610 18952 19616 18964
rect 19444 18924 19616 18952
rect 19444 18884 19472 18924
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 20162 18912 20168 18964
rect 20220 18912 20226 18964
rect 22370 18912 22376 18964
rect 22428 18912 22434 18964
rect 23750 18912 23756 18964
rect 23808 18912 23814 18964
rect 23934 18912 23940 18964
rect 23992 18912 23998 18964
rect 24029 18955 24087 18961
rect 24029 18921 24041 18955
rect 24075 18952 24087 18955
rect 24578 18952 24584 18964
rect 24075 18924 24584 18952
rect 24075 18921 24087 18924
rect 24029 18915 24087 18921
rect 24578 18912 24584 18924
rect 24636 18912 24642 18964
rect 25866 18912 25872 18964
rect 25924 18912 25930 18964
rect 27341 18955 27399 18961
rect 27341 18952 27353 18955
rect 25976 18924 27353 18952
rect 18524 18856 19472 18884
rect 20438 18844 20444 18896
rect 20496 18884 20502 18896
rect 20496 18856 21680 18884
rect 20496 18844 20502 18856
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 6963 18788 7389 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 9401 18819 9459 18825
rect 9401 18785 9413 18819
rect 9447 18816 9459 18819
rect 10042 18816 10048 18828
rect 9447 18788 10048 18816
rect 9447 18785 9459 18788
rect 9401 18779 9459 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10962 18816 10968 18828
rect 10275 18788 10968 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 6687 18720 6776 18748
rect 6825 18751 6883 18757
rect 6687 18717 6699 18720
rect 6641 18711 6699 18717
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 7006 18748 7012 18760
rect 6871 18720 7012 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 3973 18683 4031 18689
rect 3973 18680 3985 18683
rect 3528 18652 3985 18680
rect 3528 18624 3556 18652
rect 3973 18649 3985 18652
rect 4019 18649 4031 18683
rect 3973 18643 4031 18649
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18649 4215 18683
rect 4157 18643 4215 18649
rect 1811 18584 3096 18612
rect 1811 18581 1823 18584
rect 1765 18575 1823 18581
rect 3510 18572 3516 18624
rect 3568 18572 3574 18624
rect 3602 18572 3608 18624
rect 3660 18612 3666 18624
rect 4172 18612 4200 18643
rect 6730 18640 6736 18692
rect 6788 18680 6794 18692
rect 7116 18680 7144 18711
rect 7742 18708 7748 18760
rect 7800 18748 7806 18760
rect 9033 18751 9091 18757
rect 9033 18748 9045 18751
rect 7800 18720 9045 18748
rect 7800 18708 7806 18720
rect 9033 18717 9045 18720
rect 9079 18717 9091 18751
rect 9033 18711 9091 18717
rect 9214 18708 9220 18760
rect 9272 18708 9278 18760
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 10008 18720 10149 18748
rect 10008 18708 10014 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 6788 18652 7144 18680
rect 8757 18683 8815 18689
rect 6788 18640 6794 18652
rect 8757 18649 8769 18683
rect 8803 18680 8815 18683
rect 10042 18680 10048 18692
rect 8803 18652 10048 18680
rect 8803 18649 8815 18652
rect 8757 18643 8815 18649
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10336 18680 10364 18711
rect 10410 18708 10416 18760
rect 10468 18708 10474 18760
rect 10612 18757 10640 18788
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 12434 18816 12440 18828
rect 11992 18788 12440 18816
rect 11992 18757 12020 18788
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12728 18788 13001 18816
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12728 18748 12756 18788
rect 12989 18785 13001 18788
rect 13035 18816 13047 18819
rect 13814 18816 13820 18828
rect 13035 18788 13820 18816
rect 13035 18785 13047 18788
rect 12989 18779 13047 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15197 18819 15255 18825
rect 15197 18816 15209 18819
rect 14108 18788 15209 18816
rect 14108 18760 14136 18788
rect 15197 18785 15209 18788
rect 15243 18785 15255 18819
rect 17954 18816 17960 18828
rect 15197 18779 15255 18785
rect 16316 18788 17960 18816
rect 12299 18720 12756 18748
rect 12805 18751 12863 18757
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12805 18717 12817 18751
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 11146 18680 11152 18692
rect 10336 18652 11152 18680
rect 10428 18624 10456 18652
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 12161 18683 12219 18689
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 12820 18680 12848 18711
rect 13262 18708 13268 18760
rect 13320 18708 13326 18760
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13722 18708 13728 18760
rect 13780 18708 13786 18760
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18748 13967 18751
rect 13998 18748 14004 18760
rect 13955 18720 14004 18748
rect 13955 18717 13967 18720
rect 13909 18711 13967 18717
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14090 18708 14096 18760
rect 14148 18708 14154 18760
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 14369 18751 14427 18757
rect 14369 18748 14381 18751
rect 14240 18720 14381 18748
rect 14240 18708 14246 18720
rect 14369 18717 14381 18720
rect 14415 18717 14427 18751
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14369 18711 14427 18717
rect 14476 18720 14657 18748
rect 12207 18652 13032 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 13004 18624 13032 18652
rect 13170 18640 13176 18692
rect 13228 18680 13234 18692
rect 13740 18680 13768 18708
rect 14476 18680 14504 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15105 18751 15163 18757
rect 15105 18748 15117 18751
rect 14792 18720 15117 18748
rect 14792 18708 14798 18720
rect 15105 18717 15117 18720
rect 15151 18717 15163 18751
rect 15470 18748 15476 18760
rect 15105 18711 15163 18717
rect 15304 18720 15476 18748
rect 15304 18680 15332 18720
rect 15470 18708 15476 18720
rect 15528 18748 15534 18760
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 15528 18720 15577 18748
rect 15528 18708 15534 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16316 18757 16344 18788
rect 17954 18776 17960 18788
rect 18012 18776 18018 18828
rect 19426 18825 19432 18828
rect 19404 18819 19432 18825
rect 19404 18785 19416 18819
rect 19404 18779 19432 18785
rect 19426 18776 19432 18779
rect 19484 18776 19490 18828
rect 19886 18776 19892 18828
rect 19944 18816 19950 18828
rect 19944 18788 20576 18816
rect 19944 18776 19950 18788
rect 20548 18760 20576 18788
rect 20622 18776 20628 18828
rect 20680 18776 20686 18828
rect 20717 18819 20775 18825
rect 20717 18785 20729 18819
rect 20763 18816 20775 18819
rect 20806 18816 20812 18828
rect 20763 18788 20812 18816
rect 20763 18785 20775 18788
rect 20717 18779 20775 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 20990 18776 20996 18828
rect 21048 18776 21054 18828
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15712 18720 16037 18748
rect 15712 18708 15718 18720
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 16301 18751 16359 18757
rect 16301 18717 16313 18751
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17402 18748 17408 18760
rect 17359 18720 17408 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 19536 18720 20500 18748
rect 13228 18652 14504 18680
rect 14660 18652 15332 18680
rect 13228 18640 13234 18652
rect 14660 18624 14688 18652
rect 15378 18640 15384 18692
rect 15436 18640 15442 18692
rect 18785 18683 18843 18689
rect 18785 18649 18797 18683
rect 18831 18680 18843 18683
rect 18874 18680 18880 18692
rect 18831 18652 18880 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 18874 18640 18880 18652
rect 18932 18680 18938 18692
rect 19150 18680 19156 18692
rect 18932 18652 19156 18680
rect 18932 18640 18938 18652
rect 19150 18640 19156 18652
rect 19208 18640 19214 18692
rect 19536 18624 19564 18720
rect 19794 18640 19800 18692
rect 19852 18680 19858 18692
rect 20162 18689 20168 18692
rect 20149 18683 20168 18689
rect 19852 18652 20116 18680
rect 19852 18640 19858 18652
rect 3660 18584 4200 18612
rect 3660 18572 3666 18584
rect 10410 18572 10416 18624
rect 10468 18572 10474 18624
rect 12986 18572 12992 18624
rect 13044 18572 13050 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13596 18584 13737 18612
rect 13596 18572 13602 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 13725 18575 13783 18581
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 13964 18584 14197 18612
rect 13964 18572 13970 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 14642 18572 14648 18624
rect 14700 18572 14706 18624
rect 15470 18572 15476 18624
rect 15528 18572 15534 18624
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16022 18612 16028 18624
rect 15804 18584 16028 18612
rect 15804 18572 15810 18584
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16206 18572 16212 18624
rect 16264 18572 16270 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 17034 18612 17040 18624
rect 16816 18584 17040 18612
rect 16816 18572 16822 18584
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18572 17190 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 18417 18615 18475 18621
rect 18417 18612 18429 18615
rect 18196 18584 18429 18612
rect 18196 18572 18202 18584
rect 18417 18581 18429 18584
rect 18463 18581 18475 18615
rect 18417 18575 18475 18581
rect 18585 18615 18643 18621
rect 18585 18581 18597 18615
rect 18631 18612 18643 18615
rect 19058 18612 19064 18624
rect 18631 18584 19064 18612
rect 18631 18581 18643 18584
rect 18585 18575 18643 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 19518 18572 19524 18624
rect 19576 18572 19582 18624
rect 19610 18572 19616 18624
rect 19668 18572 19674 18624
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 19981 18615 20039 18621
rect 19981 18612 19993 18615
rect 19944 18584 19993 18612
rect 19944 18572 19950 18584
rect 19981 18581 19993 18584
rect 20027 18581 20039 18615
rect 20088 18612 20116 18652
rect 20149 18649 20161 18683
rect 20149 18643 20168 18649
rect 20162 18640 20168 18643
rect 20220 18640 20226 18692
rect 20349 18683 20407 18689
rect 20349 18649 20361 18683
rect 20395 18649 20407 18683
rect 20472 18680 20500 18720
rect 20530 18708 20536 18760
rect 20588 18748 20594 18760
rect 21008 18748 21036 18776
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20588 18720 21097 18748
rect 20588 18708 20594 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21181 18751 21239 18757
rect 21181 18717 21193 18751
rect 21227 18748 21239 18751
rect 21284 18748 21312 18856
rect 21227 18720 21312 18748
rect 21227 18717 21239 18720
rect 21181 18711 21239 18717
rect 21269 18683 21327 18689
rect 20472 18652 21129 18680
rect 20349 18643 20407 18649
rect 20364 18612 20392 18643
rect 20990 18612 20996 18624
rect 20088 18584 20996 18612
rect 19981 18575 20039 18581
rect 20990 18572 20996 18584
rect 21048 18572 21054 18624
rect 21101 18612 21129 18652
rect 21269 18649 21281 18683
rect 21315 18649 21327 18683
rect 21269 18643 21327 18649
rect 21545 18683 21603 18689
rect 21545 18649 21557 18683
rect 21591 18649 21603 18683
rect 21652 18680 21680 18856
rect 21726 18844 21732 18896
rect 21784 18884 21790 18896
rect 21784 18856 22968 18884
rect 21784 18844 21790 18856
rect 21928 18825 21956 18856
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18785 21971 18819
rect 21913 18779 21971 18785
rect 22278 18776 22284 18828
rect 22336 18816 22342 18828
rect 22830 18816 22836 18828
rect 22336 18788 22836 18816
rect 22336 18776 22342 18788
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 22940 18816 22968 18856
rect 23566 18844 23572 18896
rect 23624 18844 23630 18896
rect 23952 18884 23980 18912
rect 25976 18884 26004 18924
rect 27341 18921 27353 18924
rect 27387 18921 27399 18955
rect 27341 18915 27399 18921
rect 23952 18856 26004 18884
rect 25682 18816 25688 18828
rect 22940 18788 25688 18816
rect 25682 18776 25688 18788
rect 25740 18776 25746 18828
rect 25958 18776 25964 18828
rect 26016 18776 26022 18828
rect 22554 18708 22560 18760
rect 22612 18708 22618 18760
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 26234 18757 26240 18760
rect 25501 18751 25559 18757
rect 23716 18720 24256 18748
rect 23716 18708 23722 18720
rect 24228 18692 24256 18720
rect 25501 18717 25513 18751
rect 25547 18748 25559 18751
rect 26228 18748 26240 18757
rect 25547 18720 26096 18748
rect 26195 18720 26240 18748
rect 25547 18717 25559 18720
rect 25501 18711 25559 18717
rect 22005 18683 22063 18689
rect 22005 18680 22017 18683
rect 21652 18652 22017 18680
rect 21545 18643 21603 18649
rect 22005 18649 22017 18652
rect 22051 18649 22063 18683
rect 22373 18683 22431 18689
rect 22373 18680 22385 18683
rect 22005 18643 22063 18649
rect 22112 18652 22385 18680
rect 21284 18612 21312 18643
rect 21560 18612 21588 18643
rect 21101 18584 21588 18612
rect 21818 18572 21824 18624
rect 21876 18572 21882 18624
rect 21910 18572 21916 18624
rect 21968 18612 21974 18624
rect 22112 18612 22140 18652
rect 22373 18649 22385 18652
rect 22419 18649 22431 18683
rect 22373 18643 22431 18649
rect 23293 18683 23351 18689
rect 23293 18649 23305 18683
rect 23339 18680 23351 18683
rect 23474 18680 23480 18692
rect 23339 18652 23480 18680
rect 23339 18649 23351 18652
rect 23293 18643 23351 18649
rect 23474 18640 23480 18652
rect 23532 18680 23538 18692
rect 24118 18680 24124 18692
rect 23532 18652 24124 18680
rect 23532 18640 23538 18652
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 24210 18640 24216 18692
rect 24268 18640 24274 18692
rect 25685 18683 25743 18689
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 26068 18680 26096 18720
rect 26228 18711 26240 18720
rect 26234 18708 26240 18711
rect 26292 18708 26298 18760
rect 26694 18680 26700 18692
rect 25731 18652 26004 18680
rect 26068 18652 26700 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 25976 18624 26004 18652
rect 26694 18640 26700 18652
rect 26752 18640 26758 18692
rect 21968 18584 22140 18612
rect 22189 18615 22247 18621
rect 21968 18572 21974 18584
rect 22189 18581 22201 18615
rect 22235 18612 22247 18615
rect 22278 18612 22284 18624
rect 22235 18584 22284 18612
rect 22235 18581 22247 18584
rect 22189 18575 22247 18581
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 22833 18615 22891 18621
rect 22833 18612 22845 18615
rect 22796 18584 22845 18612
rect 22796 18572 22802 18584
rect 22833 18581 22845 18584
rect 22879 18581 22891 18615
rect 22833 18575 22891 18581
rect 23842 18572 23848 18624
rect 23900 18572 23906 18624
rect 24026 18621 24032 18624
rect 24013 18615 24032 18621
rect 24013 18581 24025 18615
rect 24013 18575 24032 18581
rect 24026 18572 24032 18575
rect 24084 18572 24090 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 1762 18368 1768 18420
rect 1820 18368 1826 18420
rect 2314 18368 2320 18420
rect 2372 18368 2378 18420
rect 3234 18368 3240 18420
rect 3292 18368 3298 18420
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4856 18380 4905 18408
rect 4856 18368 4862 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5166 18368 5172 18420
rect 5224 18368 5230 18420
rect 6914 18408 6920 18420
rect 5552 18380 6920 18408
rect 1780 18340 1808 18368
rect 2590 18340 2596 18352
rect 1780 18312 2596 18340
rect 2590 18300 2596 18312
rect 2648 18340 2654 18352
rect 3252 18340 3280 18368
rect 2648 18312 3004 18340
rect 2648 18300 2654 18312
rect 1762 18232 1768 18284
rect 1820 18272 1826 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1820 18244 2053 18272
rect 1820 18232 1826 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2314 18232 2320 18284
rect 2372 18232 2378 18284
rect 2498 18232 2504 18284
rect 2556 18232 2562 18284
rect 2976 18281 3004 18312
rect 3252 18312 3832 18340
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2608 18244 2881 18272
rect 2332 18204 2360 18232
rect 2608 18204 2636 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3252 18272 3280 18312
rect 3007 18244 3280 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 2332 18176 2636 18204
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18173 2835 18207
rect 2884 18204 2912 18235
rect 3326 18232 3332 18284
rect 3384 18232 3390 18284
rect 3528 18281 3556 18312
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 3602 18232 3608 18284
rect 3660 18232 3666 18284
rect 3804 18281 3832 18312
rect 4430 18300 4436 18352
rect 4488 18340 4494 18352
rect 5442 18340 5448 18352
rect 4488 18312 5448 18340
rect 4488 18300 4494 18312
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 4338 18272 4344 18284
rect 3789 18235 3847 18241
rect 3896 18244 4344 18272
rect 3620 18204 3648 18232
rect 2884 18176 3648 18204
rect 2777 18167 2835 18173
rect 2682 18096 2688 18148
rect 2740 18136 2746 18148
rect 2792 18136 2820 18167
rect 3326 18136 3332 18148
rect 2740 18108 3332 18136
rect 2740 18096 2746 18108
rect 3326 18096 3332 18108
rect 3384 18136 3390 18148
rect 3896 18136 3924 18244
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5077 18235 5135 18241
rect 5092 18204 5120 18235
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5353 18275 5411 18281
rect 5353 18272 5365 18275
rect 5316 18244 5365 18272
rect 5316 18232 5322 18244
rect 5353 18241 5365 18244
rect 5399 18272 5411 18275
rect 5552 18272 5580 18380
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 7929 18411 7987 18417
rect 7929 18377 7941 18411
rect 7975 18408 7987 18411
rect 9306 18408 9312 18420
rect 7975 18380 9312 18408
rect 7975 18377 7987 18380
rect 7929 18371 7987 18377
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 9490 18408 9496 18420
rect 9447 18380 9496 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9416 18340 9444 18371
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 9585 18411 9643 18417
rect 9585 18377 9597 18411
rect 9631 18408 9643 18411
rect 9674 18408 9680 18420
rect 9631 18380 9680 18408
rect 9631 18377 9643 18380
rect 9585 18371 9643 18377
rect 8772 18312 9444 18340
rect 5399 18244 5580 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 5902 18232 5908 18284
rect 5960 18232 5966 18284
rect 6089 18275 6147 18281
rect 6089 18241 6101 18275
rect 6135 18272 6147 18275
rect 6641 18275 6699 18281
rect 6641 18272 6653 18275
rect 6135 18244 6653 18272
rect 6135 18241 6147 18244
rect 6089 18235 6147 18241
rect 6641 18241 6653 18244
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 6730 18232 6736 18284
rect 6788 18232 6794 18284
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 8772 18281 8800 18312
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 7800 18244 8493 18272
rect 7800 18232 7806 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18241 8815 18275
rect 8757 18235 8815 18241
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 3384 18108 3924 18136
rect 4264 18176 5120 18204
rect 3384 18096 3390 18108
rect 4264 18080 4292 18176
rect 5994 18164 6000 18216
rect 6052 18164 6058 18216
rect 6178 18164 6184 18216
rect 6236 18164 6242 18216
rect 6362 18164 6368 18216
rect 6420 18204 6426 18216
rect 6748 18204 6776 18232
rect 6420 18176 6776 18204
rect 6420 18164 6426 18176
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 6012 18136 6040 18164
rect 4856 18108 6040 18136
rect 8864 18136 8892 18235
rect 9030 18232 9036 18284
rect 9088 18232 9094 18284
rect 9122 18232 9128 18284
rect 9180 18232 9186 18284
rect 9490 18232 9496 18284
rect 9548 18232 9554 18284
rect 9398 18164 9404 18216
rect 9456 18164 9462 18216
rect 9600 18136 9628 18371
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 11296 18380 11713 18408
rect 11296 18368 11302 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 11701 18371 11759 18377
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 12216 18380 12449 18408
rect 12216 18368 12222 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13909 18411 13967 18417
rect 13909 18408 13921 18411
rect 13044 18380 13921 18408
rect 13044 18368 13050 18380
rect 13909 18377 13921 18380
rect 13955 18377 13967 18411
rect 16758 18408 16764 18420
rect 13909 18371 13967 18377
rect 14568 18380 16764 18408
rect 9950 18300 9956 18352
rect 10008 18340 10014 18352
rect 14369 18343 14427 18349
rect 14369 18340 14381 18343
rect 10008 18312 12296 18340
rect 10008 18300 10014 18312
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 10042 18272 10048 18284
rect 9723 18244 10048 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 11882 18232 11888 18284
rect 11940 18232 11946 18284
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 12032 18244 12173 18272
rect 12032 18232 12038 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12268 18272 12296 18312
rect 13924 18312 14381 18340
rect 13924 18284 13952 18312
rect 14369 18309 14381 18312
rect 14415 18309 14427 18343
rect 14369 18303 14427 18309
rect 12342 18272 12348 18284
rect 12268 18244 12348 18272
rect 12161 18235 12219 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 13906 18232 13912 18284
rect 13964 18232 13970 18284
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 14182 18272 14188 18284
rect 14139 18244 14188 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18204 12127 18207
rect 14568 18204 14596 18380
rect 16758 18368 16764 18380
rect 16816 18368 16822 18420
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 17460 18380 21925 18408
rect 17460 18368 17466 18380
rect 21913 18377 21925 18380
rect 21959 18377 21971 18411
rect 21913 18371 21971 18377
rect 22554 18368 22560 18420
rect 22612 18368 22618 18420
rect 24489 18411 24547 18417
rect 24489 18377 24501 18411
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 14642 18300 14648 18352
rect 14700 18300 14706 18352
rect 15473 18343 15531 18349
rect 15473 18309 15485 18343
rect 15519 18309 15531 18343
rect 15473 18303 15531 18309
rect 15657 18343 15715 18349
rect 15657 18309 15669 18343
rect 15703 18340 15715 18343
rect 15930 18340 15936 18352
rect 15703 18312 15936 18340
rect 15703 18309 15715 18312
rect 15657 18303 15715 18309
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15102 18272 15108 18284
rect 14967 18244 15108 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15194 18232 15200 18284
rect 15252 18272 15258 18284
rect 15488 18272 15516 18303
rect 15930 18300 15936 18312
rect 15988 18300 15994 18352
rect 17126 18349 17132 18352
rect 16025 18343 16083 18349
rect 16025 18309 16037 18343
rect 16071 18340 16083 18343
rect 16225 18343 16283 18349
rect 16071 18312 16176 18340
rect 16071 18309 16083 18312
rect 16025 18303 16083 18309
rect 15252 18244 15516 18272
rect 15252 18232 15258 18244
rect 15746 18232 15752 18284
rect 15804 18272 15810 18284
rect 15841 18275 15899 18281
rect 15841 18272 15853 18275
rect 15804 18244 15853 18272
rect 15804 18232 15810 18244
rect 15841 18241 15853 18244
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 12115 18176 14596 18204
rect 12115 18173 12127 18176
rect 12069 18167 12127 18173
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15470 18204 15476 18216
rect 14884 18176 15476 18204
rect 14884 18164 14890 18176
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 16022 18164 16028 18216
rect 16080 18164 16086 18216
rect 16148 18204 16176 18312
rect 16225 18309 16237 18343
rect 16271 18340 16283 18343
rect 17109 18343 17132 18349
rect 16271 18312 16436 18340
rect 16271 18309 16283 18312
rect 16225 18303 16283 18309
rect 16298 18204 16304 18216
rect 16148 18176 16304 18204
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 8864 18108 9628 18136
rect 11977 18139 12035 18145
rect 4856 18096 4862 18108
rect 11977 18105 11989 18139
rect 12023 18105 12035 18139
rect 11977 18099 12035 18105
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 4246 18068 4252 18080
rect 3191 18040 4252 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 8570 18028 8576 18080
rect 8628 18028 8634 18080
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18068 9275 18071
rect 9674 18068 9680 18080
rect 9263 18040 9680 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 11992 18068 12020 18099
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 14553 18139 14611 18145
rect 13228 18108 13584 18136
rect 13228 18096 13234 18108
rect 13446 18068 13452 18080
rect 11992 18040 13452 18068
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 13556 18068 13584 18108
rect 14553 18105 14565 18139
rect 14599 18136 14611 18139
rect 15378 18136 15384 18148
rect 14599 18108 15384 18136
rect 14599 18105 14611 18108
rect 14553 18099 14611 18105
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 16040 18136 16068 18164
rect 16408 18136 16436 18312
rect 17109 18309 17121 18343
rect 17109 18303 17132 18309
rect 17126 18300 17132 18303
rect 17184 18300 17190 18352
rect 17310 18300 17316 18352
rect 17368 18340 17374 18352
rect 17368 18312 18552 18340
rect 17368 18300 17374 18312
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18272 16911 18275
rect 16942 18272 16948 18284
rect 16899 18244 16948 18272
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 16040 18108 16436 18136
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 13556 18040 14657 18068
rect 14645 18037 14657 18040
rect 14691 18068 14703 18071
rect 14734 18068 14740 18080
rect 14691 18040 14740 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15286 18068 15292 18080
rect 15151 18040 15292 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15286 18028 15292 18040
rect 15344 18068 15350 18080
rect 15654 18068 15660 18080
rect 15344 18040 15660 18068
rect 15344 18028 15350 18040
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 16209 18071 16267 18077
rect 16209 18068 16221 18071
rect 15988 18040 16221 18068
rect 15988 18028 15994 18040
rect 16209 18037 16221 18040
rect 16255 18037 16267 18071
rect 16209 18031 16267 18037
rect 16393 18071 16451 18077
rect 16393 18037 16405 18071
rect 16439 18068 16451 18071
rect 16758 18068 16764 18080
rect 16439 18040 16764 18068
rect 16439 18037 16451 18040
rect 16393 18031 16451 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 16868 18068 16896 18235
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18524 18281 18552 18312
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 20898 18349 20904 18352
rect 20885 18343 20904 18349
rect 18748 18312 20852 18340
rect 18748 18300 18754 18312
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 18012 18244 18337 18272
rect 18012 18232 18018 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19300 18244 19533 18272
rect 19300 18232 19306 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 20824 18272 20852 18312
rect 20885 18309 20897 18343
rect 20885 18303 20904 18309
rect 20898 18300 20904 18303
rect 20956 18300 20962 18352
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 21085 18343 21143 18349
rect 21085 18340 21097 18343
rect 21048 18312 21097 18340
rect 21048 18300 21054 18312
rect 21085 18309 21097 18312
rect 21131 18309 21143 18343
rect 21085 18303 21143 18309
rect 22370 18300 22376 18352
rect 22428 18300 22434 18352
rect 24504 18340 24532 18371
rect 25958 18368 25964 18420
rect 26016 18368 26022 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18377 26295 18411
rect 26237 18371 26295 18377
rect 24826 18343 24884 18349
rect 24826 18340 24838 18343
rect 22848 18312 23427 18340
rect 24504 18312 24838 18340
rect 22848 18281 22876 18312
rect 22104 18275 22162 18281
rect 20824 18244 22064 18272
rect 19521 18235 19579 18241
rect 18230 18164 18236 18216
rect 18288 18164 18294 18216
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18204 18751 18207
rect 19058 18204 19064 18216
rect 18739 18176 19064 18204
rect 18739 18173 18751 18176
rect 18693 18167 18751 18173
rect 19058 18164 19064 18176
rect 19116 18204 19122 18216
rect 21910 18204 21916 18216
rect 19116 18176 21916 18204
rect 19116 18164 19122 18176
rect 21910 18164 21916 18176
rect 21968 18164 21974 18216
rect 18248 18136 18276 18164
rect 20530 18136 20536 18148
rect 18248 18108 20536 18136
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20717 18139 20775 18145
rect 20717 18105 20729 18139
rect 20763 18136 20775 18139
rect 21450 18136 21456 18148
rect 20763 18108 21456 18136
rect 20763 18105 20775 18108
rect 20717 18099 20775 18105
rect 21450 18096 21456 18108
rect 21508 18096 21514 18148
rect 22036 18136 22064 18244
rect 22104 18241 22116 18275
rect 22150 18272 22162 18275
rect 22833 18275 22891 18281
rect 22150 18244 22416 18272
rect 22150 18241 22162 18244
rect 22104 18235 22162 18241
rect 22388 18216 22416 18244
rect 22833 18241 22845 18275
rect 22879 18241 22891 18275
rect 22833 18235 22891 18241
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 22278 18164 22284 18216
rect 22336 18164 22342 18216
rect 22370 18164 22376 18216
rect 22428 18164 22434 18216
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23017 18207 23075 18213
rect 23017 18204 23029 18207
rect 22980 18176 23029 18204
rect 22980 18164 22986 18176
rect 23017 18173 23029 18176
rect 23063 18173 23075 18207
rect 23124 18204 23152 18235
rect 23198 18232 23204 18284
rect 23256 18272 23262 18284
rect 23293 18275 23351 18281
rect 23293 18272 23305 18275
rect 23256 18244 23305 18272
rect 23256 18232 23262 18244
rect 23293 18241 23305 18244
rect 23339 18241 23351 18275
rect 23399 18272 23427 18312
rect 24826 18309 24838 18312
rect 24872 18309 24884 18343
rect 24826 18303 24884 18309
rect 23842 18272 23848 18284
rect 23399 18244 23848 18272
rect 23293 18235 23351 18241
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 24302 18232 24308 18284
rect 24360 18232 24366 18284
rect 25976 18272 26004 18368
rect 26252 18340 26280 18371
rect 27218 18343 27276 18349
rect 27218 18340 27230 18343
rect 26252 18312 27230 18340
rect 27218 18309 27230 18312
rect 27264 18309 27276 18343
rect 27218 18303 27276 18309
rect 24504 18244 26004 18272
rect 26053 18275 26111 18281
rect 24504 18204 24532 18244
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 26329 18275 26387 18281
rect 26329 18272 26341 18275
rect 26099 18244 26341 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 26329 18241 26341 18244
rect 26375 18241 26387 18275
rect 26329 18235 26387 18241
rect 26513 18275 26571 18281
rect 26513 18241 26525 18275
rect 26559 18241 26571 18275
rect 26513 18235 26571 18241
rect 23124 18176 24532 18204
rect 23017 18167 23075 18173
rect 24578 18164 24584 18216
rect 24636 18164 24642 18216
rect 22036 18108 24633 18136
rect 17770 18068 17776 18080
rect 16868 18040 17776 18068
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 18230 18028 18236 18080
rect 18288 18028 18294 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19518 18068 19524 18080
rect 19383 18040 19524 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21358 18068 21364 18080
rect 20947 18040 21364 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 22373 18071 22431 18077
rect 22373 18037 22385 18071
rect 22419 18068 22431 18071
rect 22462 18068 22468 18080
rect 22419 18040 22468 18068
rect 22419 18037 22431 18040
rect 22373 18031 22431 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 22922 18028 22928 18080
rect 22980 18028 22986 18080
rect 24605 18068 24633 18108
rect 26528 18080 26556 18235
rect 26694 18232 26700 18284
rect 26752 18232 26758 18284
rect 26970 18164 26976 18216
rect 27028 18164 27034 18216
rect 26510 18068 26516 18080
rect 24605 18040 26516 18068
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 26878 18028 26884 18080
rect 26936 18068 26942 18080
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 26936 18040 28365 18068
rect 26936 18028 26942 18040
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 28353 18031 28411 18037
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1820 17836 1869 17864
rect 1820 17824 1826 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 1857 17827 1915 17833
rect 3510 17824 3516 17876
rect 3568 17824 3574 17876
rect 3786 17824 3792 17876
rect 3844 17864 3850 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 3844 17836 4261 17864
rect 3844 17824 3850 17836
rect 4249 17833 4261 17836
rect 4295 17833 4307 17867
rect 4249 17827 4307 17833
rect 4798 17824 4804 17876
rect 4856 17824 4862 17876
rect 10229 17867 10287 17873
rect 10229 17833 10241 17867
rect 10275 17864 10287 17867
rect 10318 17864 10324 17876
rect 10275 17836 10324 17864
rect 10275 17833 10287 17836
rect 10229 17827 10287 17833
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10778 17824 10784 17876
rect 10836 17864 10842 17876
rect 10873 17867 10931 17873
rect 10873 17864 10885 17867
rect 10836 17836 10885 17864
rect 10836 17824 10842 17836
rect 10873 17833 10885 17836
rect 10919 17833 10931 17867
rect 10873 17827 10931 17833
rect 11149 17867 11207 17873
rect 11149 17833 11161 17867
rect 11195 17833 11207 17867
rect 11149 17827 11207 17833
rect 4065 17799 4123 17805
rect 4065 17765 4077 17799
rect 4111 17796 4123 17799
rect 4816 17796 4844 17824
rect 4111 17768 4844 17796
rect 5077 17799 5135 17805
rect 4111 17765 4123 17768
rect 4065 17759 4123 17765
rect 5077 17765 5089 17799
rect 5123 17796 5135 17799
rect 5902 17796 5908 17808
rect 5123 17768 5908 17796
rect 5123 17765 5135 17768
rect 5077 17759 5135 17765
rect 5902 17756 5908 17768
rect 5960 17756 5966 17808
rect 7377 17799 7435 17805
rect 7377 17765 7389 17799
rect 7423 17796 7435 17799
rect 7650 17796 7656 17808
rect 7423 17768 7656 17796
rect 7423 17765 7435 17768
rect 7377 17759 7435 17765
rect 7650 17756 7656 17768
rect 7708 17756 7714 17808
rect 8570 17756 8576 17808
rect 8628 17796 8634 17808
rect 9398 17796 9404 17808
rect 8628 17768 9404 17796
rect 8628 17756 8634 17768
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 9456 17768 9536 17796
rect 9456 17756 9462 17768
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4212 17700 4798 17728
rect 4212 17688 4218 17700
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17629 2651 17663
rect 2593 17623 2651 17629
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 2498 17592 2504 17604
rect 1728 17564 2504 17592
rect 1728 17552 1734 17564
rect 2498 17552 2504 17564
rect 2556 17592 2562 17604
rect 2608 17592 2636 17623
rect 3234 17620 3240 17672
rect 3292 17620 3298 17672
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3878 17620 3884 17672
rect 3936 17620 3942 17672
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4770 17669 4798 17700
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 8846 17728 8852 17740
rect 5224 17700 8852 17728
rect 5224 17688 5230 17700
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 9508 17728 9536 17768
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 9769 17799 9827 17805
rect 9769 17796 9781 17799
rect 9732 17768 9781 17796
rect 9732 17756 9738 17768
rect 9769 17765 9781 17768
rect 9815 17765 9827 17799
rect 9769 17759 9827 17765
rect 9861 17799 9919 17805
rect 9861 17765 9873 17799
rect 9907 17796 9919 17799
rect 10137 17799 10195 17805
rect 10137 17796 10149 17799
rect 9907 17768 10149 17796
rect 9907 17765 9919 17768
rect 9861 17759 9919 17765
rect 10137 17765 10149 17768
rect 10183 17796 10195 17799
rect 10505 17799 10563 17805
rect 10505 17796 10517 17799
rect 10183 17768 10517 17796
rect 10183 17765 10195 17768
rect 10137 17759 10195 17765
rect 10505 17765 10517 17768
rect 10551 17765 10563 17799
rect 10505 17759 10563 17765
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9508 17700 9965 17728
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 9953 17691 10011 17697
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17728 10379 17731
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10367 17700 10977 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 4433 17663 4491 17669
rect 4433 17660 4445 17663
rect 4304 17632 4445 17660
rect 4304 17620 4310 17632
rect 4433 17629 4445 17632
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 4719 17663 4798 17669
rect 4719 17629 4731 17663
rect 4765 17632 4798 17663
rect 4765 17629 4777 17632
rect 4719 17623 4777 17629
rect 4890 17620 4896 17672
rect 4948 17620 4954 17672
rect 5031 17663 5089 17669
rect 5031 17629 5043 17663
rect 5077 17654 5089 17663
rect 5258 17660 5264 17672
rect 5184 17654 5264 17660
rect 5077 17632 5264 17654
rect 5077 17629 5212 17632
rect 5031 17626 5212 17629
rect 5031 17623 5089 17626
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 7009 17663 7067 17669
rect 6196 17632 6500 17660
rect 6196 17592 6224 17632
rect 2556 17564 2636 17592
rect 3988 17564 6224 17592
rect 2556 17552 2562 17564
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 1873 17527 1931 17533
rect 1873 17524 1885 17527
rect 1636 17496 1885 17524
rect 1636 17484 1642 17496
rect 1873 17493 1885 17496
rect 1919 17493 1931 17527
rect 1873 17487 1931 17493
rect 2041 17527 2099 17533
rect 2041 17493 2053 17527
rect 2087 17524 2099 17527
rect 3988 17524 4016 17564
rect 6362 17552 6368 17604
rect 6420 17552 6426 17604
rect 6472 17592 6500 17632
rect 7009 17629 7021 17663
rect 7055 17660 7067 17663
rect 7098 17660 7104 17672
rect 7055 17632 7104 17660
rect 7055 17629 7067 17632
rect 7009 17623 7067 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8757 17663 8815 17669
rect 8757 17660 8769 17663
rect 8628 17632 8769 17660
rect 8628 17620 8634 17632
rect 8757 17629 8769 17632
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 7193 17595 7251 17601
rect 7193 17592 7205 17595
rect 6472 17564 7205 17592
rect 7193 17561 7205 17564
rect 7239 17561 7251 17595
rect 7193 17555 7251 17561
rect 2087 17496 4016 17524
rect 4617 17527 4675 17533
rect 2087 17493 2099 17496
rect 2041 17487 2099 17493
rect 4617 17493 4629 17527
rect 4663 17524 4675 17527
rect 5074 17524 5080 17536
rect 4663 17496 5080 17524
rect 4663 17493 4675 17496
rect 4617 17487 4675 17493
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 5626 17484 5632 17536
rect 5684 17524 5690 17536
rect 5721 17527 5779 17533
rect 5721 17524 5733 17527
rect 5684 17496 5733 17524
rect 5684 17484 5690 17496
rect 5721 17493 5733 17496
rect 5767 17524 5779 17527
rect 6380 17524 6408 17552
rect 5767 17496 6408 17524
rect 8772 17524 8800 17623
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9456 17632 9689 17660
rect 9456 17620 9462 17632
rect 9677 17629 9689 17632
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 9968 17592 9996 17691
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10091 17632 10425 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10413 17629 10425 17632
rect 10459 17660 10471 17663
rect 10502 17660 10508 17672
rect 10459 17632 10508 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 10704 17669 10732 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 11164 17592 11192 17827
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 12676 17836 13277 17864
rect 12676 17824 12682 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 13872 17836 14657 17864
rect 13872 17824 13878 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16574 17864 16580 17876
rect 15896 17836 16580 17864
rect 15896 17824 15902 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16758 17824 16764 17876
rect 16816 17824 16822 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 19343 17864 19349 17876
rect 16908 17836 19349 17864
rect 16908 17824 16914 17836
rect 19343 17824 19349 17836
rect 19401 17824 19407 17876
rect 19469 17867 19527 17873
rect 19469 17833 19481 17867
rect 19515 17864 19527 17867
rect 19515 17833 19544 17864
rect 19469 17827 19544 17833
rect 11698 17756 11704 17808
rect 11756 17756 11762 17808
rect 13170 17756 13176 17808
rect 13228 17756 13234 17808
rect 14274 17756 14280 17808
rect 14332 17796 14338 17808
rect 14369 17799 14427 17805
rect 14369 17796 14381 17799
rect 14332 17768 14381 17796
rect 14332 17756 14338 17768
rect 14369 17765 14381 17768
rect 14415 17765 14427 17799
rect 14369 17759 14427 17765
rect 16669 17799 16727 17805
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 19245 17799 19303 17805
rect 19245 17796 19257 17799
rect 16715 17768 19257 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 19245 17765 19257 17768
rect 19291 17765 19303 17799
rect 19516 17796 19544 17827
rect 22278 17824 22284 17876
rect 22336 17864 22342 17876
rect 23017 17867 23075 17873
rect 23017 17864 23029 17867
rect 22336 17836 23029 17864
rect 22336 17824 22342 17836
rect 23017 17833 23029 17836
rect 23063 17833 23075 17867
rect 23017 17827 23075 17833
rect 23492 17836 24256 17864
rect 23492 17796 23520 17836
rect 19516 17768 23520 17796
rect 19245 17759 19303 17765
rect 23566 17756 23572 17808
rect 23624 17756 23630 17808
rect 23934 17756 23940 17808
rect 23992 17756 23998 17808
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 11716 17660 11744 17756
rect 11471 17632 11744 17660
rect 11885 17663 11943 17669
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 11885 17629 11897 17663
rect 11931 17660 11943 17663
rect 13188 17660 13216 17756
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13320 17700 13829 17728
rect 13320 17688 13326 17700
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 14550 17728 14556 17740
rect 13817 17691 13875 17697
rect 13924 17700 14556 17728
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 11931 17632 12434 17660
rect 13188 17632 13553 17660
rect 11931 17629 11943 17632
rect 11885 17623 11943 17629
rect 12158 17601 12164 17604
rect 9968 17564 11192 17592
rect 12152 17555 12164 17601
rect 12158 17552 12164 17555
rect 12216 17552 12222 17604
rect 12406 17592 12434 17632
rect 13541 17629 13553 17632
rect 13587 17629 13599 17663
rect 13924 17660 13952 17700
rect 14550 17688 14556 17700
rect 14608 17728 14614 17740
rect 14921 17731 14979 17737
rect 14921 17728 14933 17731
rect 14608 17700 14933 17728
rect 14608 17688 14614 17700
rect 14921 17697 14933 17700
rect 14967 17697 14979 17731
rect 14921 17691 14979 17697
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 16853 17731 16911 17737
rect 16356 17700 16528 17728
rect 16356 17688 16362 17700
rect 13541 17623 13599 17629
rect 13832 17632 13952 17660
rect 13170 17592 13176 17604
rect 12406 17564 13176 17592
rect 13170 17552 13176 17564
rect 13228 17592 13234 17604
rect 13832 17592 13860 17632
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14792 17632 14841 17660
rect 14792 17620 14798 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16264 17632 16405 17660
rect 16264 17620 16270 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 13228 17564 13860 17592
rect 13228 17552 13234 17564
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 14056 17564 14197 17592
rect 14056 17552 14062 17564
rect 14185 17561 14197 17564
rect 14231 17561 14243 17595
rect 14185 17555 14243 17561
rect 15188 17595 15246 17601
rect 15188 17561 15200 17595
rect 15234 17592 15246 17595
rect 15378 17592 15384 17604
rect 15234 17564 15384 17592
rect 15234 17561 15246 17564
rect 15188 17555 15246 17561
rect 9950 17524 9956 17536
rect 8772 17496 9956 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 13078 17524 13084 17536
rect 11848 17496 13084 17524
rect 11848 17484 11854 17496
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 14200 17524 14228 17555
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 16500 17592 16528 17700
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 19886 17728 19892 17740
rect 16899 17700 19892 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 23106 17688 23112 17740
rect 23164 17688 23170 17740
rect 23584 17728 23612 17756
rect 23308 17700 23612 17728
rect 24228 17728 24256 17836
rect 24302 17824 24308 17876
rect 24360 17864 24366 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 24360 17836 24409 17864
rect 24360 17824 24366 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 24397 17827 24455 17833
rect 25130 17824 25136 17876
rect 25188 17864 25194 17876
rect 28537 17867 28595 17873
rect 28537 17864 28549 17867
rect 25188 17836 28549 17864
rect 25188 17824 25194 17836
rect 28537 17833 28549 17836
rect 28583 17833 28595 17867
rect 28537 17827 28595 17833
rect 26510 17756 26516 17808
rect 26568 17796 26574 17808
rect 26605 17799 26663 17805
rect 26605 17796 26617 17799
rect 26568 17768 26617 17796
rect 26568 17756 26574 17768
rect 26605 17765 26617 17768
rect 26651 17765 26663 17799
rect 26605 17759 26663 17765
rect 24228 17700 25360 17728
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 19518 17660 19524 17672
rect 19398 17635 19524 17660
rect 19383 17632 19524 17635
rect 19383 17629 19441 17632
rect 16942 17592 16948 17604
rect 16500 17564 16948 17592
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 19383 17595 19395 17629
rect 19429 17595 19441 17629
rect 19518 17620 19524 17632
rect 19576 17660 19582 17672
rect 19576 17632 19932 17660
rect 19576 17620 19582 17632
rect 19383 17589 19441 17595
rect 19610 17552 19616 17604
rect 19668 17552 19674 17604
rect 19904 17592 19932 17632
rect 19978 17620 19984 17672
rect 20036 17620 20042 17672
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21048 17632 21373 17660
rect 21048 17620 21054 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 20622 17592 20628 17604
rect 19904 17564 20628 17592
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 23124 17592 23152 17688
rect 23198 17669 23204 17672
rect 23196 17623 23204 17669
rect 23198 17620 23204 17623
rect 23256 17620 23262 17672
rect 23308 17669 23336 17700
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23568 17663 23626 17669
rect 23568 17629 23580 17663
rect 23614 17629 23626 17663
rect 23568 17623 23626 17629
rect 23382 17592 23388 17604
rect 23124 17564 23388 17592
rect 23382 17552 23388 17564
rect 23440 17552 23446 17604
rect 23583 17592 23611 17623
rect 23658 17620 23664 17672
rect 23716 17620 23722 17672
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 25130 17660 25136 17672
rect 24627 17632 25136 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24596 17592 24624 17623
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17629 25283 17663
rect 25332 17660 25360 17700
rect 26878 17660 26884 17672
rect 25332 17632 26884 17660
rect 25225 17623 25283 17629
rect 23583 17564 24624 17592
rect 24762 17552 24768 17604
rect 24820 17552 24826 17604
rect 14826 17524 14832 17536
rect 14200 17496 14832 17524
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 16298 17484 16304 17536
rect 16356 17484 16362 17536
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16632 17496 17141 17524
rect 16632 17484 16638 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 20165 17527 20223 17533
rect 20165 17493 20177 17527
rect 20211 17524 20223 17527
rect 20254 17524 20260 17536
rect 20211 17496 20260 17524
rect 20211 17493 20223 17496
rect 20165 17487 20223 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 21358 17484 21364 17536
rect 21416 17524 21422 17536
rect 21545 17527 21603 17533
rect 21545 17524 21557 17527
rect 21416 17496 21557 17524
rect 21416 17484 21422 17496
rect 21545 17493 21557 17496
rect 21591 17524 21603 17527
rect 24578 17524 24584 17536
rect 21591 17496 24584 17524
rect 21591 17493 21603 17496
rect 21545 17487 21603 17493
rect 24578 17484 24584 17496
rect 24636 17524 24642 17536
rect 25240 17524 25268 17623
rect 26878 17620 26884 17632
rect 26936 17620 26942 17672
rect 26970 17620 26976 17672
rect 27028 17660 27034 17672
rect 27157 17663 27215 17669
rect 27157 17660 27169 17663
rect 27028 17632 27169 17660
rect 27028 17620 27034 17632
rect 27157 17629 27169 17632
rect 27203 17629 27215 17663
rect 27157 17623 27215 17629
rect 25498 17601 25504 17604
rect 25492 17555 25504 17601
rect 25498 17552 25504 17555
rect 25556 17552 25562 17604
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 26694 17592 26700 17604
rect 26292 17564 26700 17592
rect 26292 17552 26298 17564
rect 26694 17552 26700 17564
rect 26752 17552 26758 17604
rect 26988 17524 27016 17620
rect 27430 17601 27436 17604
rect 27424 17555 27436 17601
rect 27430 17552 27436 17555
rect 27488 17552 27494 17604
rect 24636 17496 27016 17524
rect 24636 17484 24642 17496
rect 27062 17484 27068 17536
rect 27120 17484 27126 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 2130 17280 2136 17332
rect 2188 17280 2194 17332
rect 2777 17323 2835 17329
rect 2777 17289 2789 17323
rect 2823 17289 2835 17323
rect 2777 17283 2835 17289
rect 1670 17212 1676 17264
rect 1728 17252 1734 17264
rect 1949 17255 2007 17261
rect 1949 17252 1961 17255
rect 1728 17224 1961 17252
rect 1728 17212 1734 17224
rect 1949 17221 1961 17224
rect 1995 17252 2007 17255
rect 2593 17255 2651 17261
rect 2593 17252 2605 17255
rect 1995 17224 2605 17252
rect 1995 17221 2007 17224
rect 1949 17215 2007 17221
rect 2593 17221 2605 17224
rect 2639 17221 2651 17255
rect 2792 17252 2820 17283
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 3326 17280 3332 17332
rect 3384 17280 3390 17332
rect 3878 17280 3884 17332
rect 3936 17280 3942 17332
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 5350 17320 5356 17332
rect 5307 17292 5356 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 7653 17323 7711 17329
rect 7653 17320 7665 17323
rect 5592 17292 7665 17320
rect 5592 17280 5598 17292
rect 7653 17289 7665 17292
rect 7699 17320 7711 17323
rect 12066 17320 12072 17332
rect 7699 17292 12072 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13004 17292 13829 17320
rect 3896 17252 3924 17280
rect 2792 17224 3924 17252
rect 5552 17252 5580 17280
rect 5552 17224 5672 17252
rect 2593 17215 2651 17221
rect 2866 17144 2872 17196
rect 2924 17144 2930 17196
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 3252 17116 3280 17147
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 5644 17193 5672 17224
rect 6086 17212 6092 17264
rect 6144 17252 6150 17264
rect 6144 17224 6675 17252
rect 6144 17212 6150 17224
rect 6647 17193 6675 17224
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 7929 17255 7987 17261
rect 7929 17252 7941 17255
rect 7800 17224 7941 17252
rect 7800 17212 7806 17224
rect 7929 17221 7941 17224
rect 7975 17252 7987 17255
rect 7975 17224 9352 17252
rect 7975 17221 7987 17224
rect 7929 17215 7987 17221
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5905 17187 5963 17193
rect 5905 17184 5917 17187
rect 5828 17168 5917 17184
rect 5629 17147 5687 17153
rect 5736 17156 5917 17168
rect 5736 17140 5856 17156
rect 5905 17153 5917 17156
rect 5951 17184 5963 17187
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 5951 17156 6561 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 1596 17088 3280 17116
rect 1596 17060 1624 17088
rect 1578 17008 1584 17060
rect 1636 17008 1642 17060
rect 2225 17051 2283 17057
rect 2225 17048 2237 17051
rect 1964 17020 2237 17048
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 1964 16989 1992 17020
rect 2225 17017 2237 17020
rect 2271 17017 2283 17051
rect 2225 17011 2283 17017
rect 2608 16989 2636 17088
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 5736 17116 5764 17140
rect 4948 17088 5764 17116
rect 6564 17116 6592 17147
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7006 17144 7012 17196
rect 7064 17144 7070 17196
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8662 17184 8668 17196
rect 8159 17156 8668 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 9324 17184 9352 17224
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 11756 17224 12664 17252
rect 11756 17212 11762 17224
rect 12250 17184 12256 17196
rect 9324 17156 12256 17184
rect 8849 17147 8907 17153
rect 6932 17116 6960 17144
rect 6564 17088 6960 17116
rect 8573 17119 8631 17125
rect 4948 17076 4954 17088
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8864 17116 8892 17147
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 12345 17187 12403 17193
rect 12345 17153 12357 17187
rect 12391 17184 12403 17187
rect 12526 17184 12532 17196
rect 12391 17156 12532 17184
rect 12391 17153 12403 17156
rect 12345 17147 12403 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 8619 17088 8892 17116
rect 12636 17116 12664 17224
rect 13004 17193 13032 17292
rect 13817 17289 13829 17292
rect 13863 17320 13875 17323
rect 14274 17320 14280 17332
rect 13863 17292 14280 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 14642 17320 14648 17332
rect 14599 17292 14648 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15194 17280 15200 17332
rect 15252 17280 15258 17332
rect 15378 17280 15384 17332
rect 15436 17280 15442 17332
rect 21082 17280 21088 17332
rect 21140 17320 21146 17332
rect 21361 17323 21419 17329
rect 21361 17320 21373 17323
rect 21140 17292 21373 17320
rect 21140 17280 21146 17292
rect 21361 17289 21373 17292
rect 21407 17289 21419 17323
rect 21361 17283 21419 17289
rect 21542 17280 21548 17332
rect 21600 17320 21606 17332
rect 21600 17292 22324 17320
rect 21600 17280 21606 17292
rect 13096 17224 13860 17252
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13096 17125 13124 17224
rect 13262 17144 13268 17196
rect 13320 17144 13326 17196
rect 13354 17144 13360 17196
rect 13412 17188 13418 17196
rect 13412 17184 13492 17188
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13412 17160 13645 17184
rect 13412 17144 13418 17160
rect 13464 17156 13645 17160
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13722 17144 13728 17196
rect 13780 17144 13786 17196
rect 13832 17184 13860 17224
rect 14090 17212 14096 17264
rect 14148 17252 14154 17264
rect 14148 17224 14688 17252
rect 14148 17212 14154 17224
rect 14660 17193 14688 17224
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 13832 17156 14381 17184
rect 14369 17153 14381 17156
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 15212 17184 15240 17280
rect 22296 17261 22324 17292
rect 23198 17280 23204 17332
rect 23256 17280 23262 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 23566 17320 23572 17332
rect 23523 17292 23572 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 23934 17280 23940 17332
rect 23992 17280 23998 17332
rect 24670 17280 24676 17332
rect 24728 17280 24734 17332
rect 25498 17280 25504 17332
rect 25556 17280 25562 17332
rect 27430 17280 27436 17332
rect 27488 17280 27494 17332
rect 22281 17255 22339 17261
rect 15672 17224 20392 17252
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15212 17156 15577 17184
rect 14645 17147 14703 17153
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 12636 17088 13093 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13081 17079 13139 17085
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13372 17116 13400 17144
rect 13219 17088 13400 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 14182 17076 14188 17128
rect 14240 17076 14246 17128
rect 5902 17008 5908 17060
rect 5960 17008 5966 17060
rect 5994 17008 6000 17060
rect 6052 17048 6058 17060
rect 6457 17051 6515 17057
rect 6457 17048 6469 17051
rect 6052 17020 6469 17048
rect 6052 17008 6058 17020
rect 6457 17017 6469 17020
rect 6503 17017 6515 17051
rect 6457 17011 6515 17017
rect 8481 17051 8539 17057
rect 8481 17017 8493 17051
rect 8527 17048 8539 17051
rect 9122 17048 9128 17060
rect 8527 17020 9128 17048
rect 8527 17017 8539 17020
rect 8481 17011 8539 17017
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 15672 17048 15700 17224
rect 17770 17144 17776 17196
rect 17828 17144 17834 17196
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 18012 17156 18061 17184
rect 18012 17144 18018 17156
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17184 18291 17187
rect 18598 17184 18604 17196
rect 18279 17156 18604 17184
rect 18279 17153 18291 17156
rect 18233 17147 18291 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 18782 17193 18788 17196
rect 18776 17147 18788 17193
rect 18782 17144 18788 17147
rect 18840 17144 18846 17196
rect 20254 17193 20260 17196
rect 20237 17187 20260 17193
rect 20237 17153 20249 17187
rect 20237 17147 20260 17153
rect 20254 17144 20260 17147
rect 20312 17144 20318 17196
rect 20364 17184 20392 17224
rect 22281 17221 22293 17255
rect 22327 17221 22339 17255
rect 23952 17252 23980 17280
rect 24590 17255 24648 17261
rect 24590 17252 24602 17255
rect 23952 17224 24602 17252
rect 22281 17215 22339 17221
rect 24590 17221 24602 17224
rect 24636 17221 24648 17255
rect 24590 17215 24648 17221
rect 20364 17156 21036 17184
rect 17788 17116 17816 17144
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 17788 17088 18521 17116
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 21008 17116 21036 17156
rect 21542 17144 21548 17196
rect 21600 17184 21606 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21600 17156 22017 17184
rect 21600 17144 21606 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22152 17156 23029 17184
rect 22152 17144 22158 17156
rect 23017 17153 23029 17156
rect 23063 17184 23075 17187
rect 24026 17184 24032 17196
rect 23063 17156 24032 17184
rect 23063 17153 23075 17156
rect 23017 17147 23075 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 24688 17184 24716 17280
rect 26234 17212 26240 17264
rect 26292 17252 26298 17264
rect 26973 17255 27031 17261
rect 26973 17252 26985 17255
rect 26292 17224 26985 17252
rect 26292 17212 26298 17224
rect 26973 17221 26985 17224
rect 27019 17221 27031 17255
rect 26973 17215 27031 17221
rect 24857 17187 24915 17193
rect 24857 17184 24869 17187
rect 24688 17156 24869 17184
rect 24857 17153 24869 17156
rect 24903 17153 24915 17187
rect 24857 17147 24915 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17184 25375 17187
rect 25590 17184 25596 17196
rect 25363 17156 25596 17184
rect 25363 17153 25375 17156
rect 25317 17147 25375 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 27154 17144 27160 17196
rect 27212 17144 27218 17196
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17184 27399 17187
rect 27617 17187 27675 17193
rect 27617 17184 27629 17187
rect 27387 17156 27629 17184
rect 27387 17153 27399 17156
rect 27341 17147 27399 17153
rect 27617 17153 27629 17156
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 22189 17119 22247 17125
rect 20027 17085 20040 17116
rect 21008 17088 21864 17116
rect 19981 17079 20040 17085
rect 20012 17048 20040 17079
rect 9968 17020 15700 17048
rect 19444 17020 20040 17048
rect 9968 16992 9996 17020
rect 19444 16992 19472 17020
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1820 16952 1961 16980
rect 1820 16940 1826 16952
rect 1949 16949 1961 16952
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 2593 16983 2651 16989
rect 2593 16949 2605 16983
rect 2639 16949 2651 16983
rect 2593 16943 2651 16949
rect 7098 16940 7104 16992
rect 7156 16940 7162 16992
rect 8662 16940 8668 16992
rect 8720 16940 8726 16992
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 12250 16980 12256 16992
rect 10928 16952 12256 16980
rect 10928 16940 10934 16952
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 13449 16983 13507 16989
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 15746 16980 15752 16992
rect 13495 16952 15752 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 18417 16983 18475 16989
rect 18417 16949 18429 16983
rect 18463 16980 18475 16983
rect 18690 16980 18696 16992
rect 18463 16952 18696 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 19426 16940 19432 16992
rect 19484 16940 19490 16992
rect 19886 16940 19892 16992
rect 19944 16940 19950 16992
rect 20012 16980 20040 17020
rect 20990 17008 20996 17060
rect 21048 17008 21054 17060
rect 21836 17057 21864 17088
rect 22189 17085 22201 17119
rect 22235 17116 22247 17119
rect 22462 17116 22468 17128
rect 22235 17088 22468 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 22833 17119 22891 17125
rect 22833 17085 22845 17119
rect 22879 17116 22891 17119
rect 23106 17116 23112 17128
rect 22879 17088 23112 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 21821 17051 21879 17057
rect 21821 17017 21833 17051
rect 21867 17017 21879 17051
rect 21821 17011 21879 17017
rect 21008 16980 21036 17008
rect 20012 16952 21036 16980
rect 22186 16940 22192 16992
rect 22244 16940 22250 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 5994 16776 6000 16788
rect 5368 16748 6000 16776
rect 5368 16649 5396 16748
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9122 16776 9128 16788
rect 8803 16748 9128 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 9916 16748 10149 16776
rect 9916 16736 9922 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 11149 16779 11207 16785
rect 11149 16745 11161 16779
rect 11195 16776 11207 16779
rect 11974 16776 11980 16788
rect 11195 16748 11980 16776
rect 11195 16745 11207 16748
rect 11149 16739 11207 16745
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12176 16748 12388 16776
rect 9398 16668 9404 16720
rect 9456 16668 9462 16720
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 11241 16711 11299 16717
rect 11241 16708 11253 16711
rect 10284 16680 11253 16708
rect 10284 16668 10290 16680
rect 11241 16677 11253 16680
rect 11287 16677 11299 16711
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 11241 16671 11299 16677
rect 11348 16680 11713 16708
rect 5353 16643 5411 16649
rect 4264 16612 5212 16640
rect 3510 16582 3516 16584
rect 3488 16576 3516 16582
rect 3488 16542 3500 16576
rect 3488 16536 3516 16542
rect 3510 16532 3516 16536
rect 3568 16532 3574 16584
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16572 3847 16575
rect 3835 16544 4016 16572
rect 3835 16541 3847 16544
rect 3789 16535 3847 16541
rect 2038 16464 2044 16516
rect 2096 16504 2102 16516
rect 3881 16507 3939 16513
rect 3881 16504 3893 16507
rect 2096 16476 3893 16504
rect 2096 16464 2102 16476
rect 3881 16473 3893 16476
rect 3927 16473 3939 16507
rect 3881 16467 3939 16473
rect 3988 16448 4016 16544
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4264 16581 4292 16612
rect 5184 16584 5212 16612
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 9674 16600 9680 16652
rect 9732 16600 9738 16652
rect 10778 16640 10784 16652
rect 9876 16612 10784 16640
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 4212 16544 4261 16572
rect 4212 16532 4218 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16572 4859 16575
rect 4890 16572 4896 16584
rect 4847 16544 4896 16572
rect 4847 16541 4859 16544
rect 4801 16535 4859 16541
rect 4890 16532 4896 16544
rect 4948 16532 4954 16584
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 5166 16532 5172 16584
rect 5224 16532 5230 16584
rect 5537 16575 5595 16581
rect 5537 16572 5549 16575
rect 5368 16544 5549 16572
rect 4617 16507 4675 16513
rect 4617 16473 4629 16507
rect 4663 16504 4675 16507
rect 5368 16504 5396 16544
rect 5537 16541 5549 16544
rect 5583 16541 5595 16575
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 5537 16535 5595 16541
rect 5736 16544 5917 16572
rect 4663 16476 5396 16504
rect 4663 16473 4675 16476
rect 4617 16467 4675 16473
rect 4816 16448 4844 16476
rect 3559 16439 3617 16445
rect 3559 16405 3571 16439
rect 3605 16436 3617 16439
rect 3786 16436 3792 16448
rect 3605 16408 3792 16436
rect 3605 16405 3617 16408
rect 3559 16399 3617 16405
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 3970 16396 3976 16448
rect 4028 16396 4034 16448
rect 4798 16396 4804 16448
rect 4856 16396 4862 16448
rect 5368 16436 5396 16476
rect 5445 16507 5503 16513
rect 5445 16473 5457 16507
rect 5491 16504 5503 16507
rect 5736 16504 5764 16544
rect 5905 16541 5917 16544
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 7374 16532 7380 16584
rect 7432 16532 7438 16584
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 7484 16544 9597 16572
rect 7484 16504 7512 16544
rect 9585 16541 9597 16544
rect 9631 16541 9643 16575
rect 9585 16535 9643 16541
rect 7650 16513 7656 16516
rect 5491 16476 5764 16504
rect 6748 16476 7512 16504
rect 5491 16473 5503 16476
rect 5445 16467 5503 16473
rect 6748 16448 6776 16476
rect 7644 16467 7656 16513
rect 7650 16464 7656 16467
rect 7708 16464 7714 16516
rect 8754 16464 8760 16516
rect 8812 16504 8818 16516
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8812 16476 9045 16504
rect 8812 16464 8818 16476
rect 9033 16473 9045 16476
rect 9079 16473 9091 16507
rect 9692 16504 9720 16600
rect 9876 16581 9904 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 9950 16532 9956 16584
rect 10008 16532 10014 16584
rect 11348 16572 11376 16680
rect 11701 16677 11713 16680
rect 11747 16708 11759 16711
rect 12066 16708 12072 16720
rect 11747 16680 12072 16708
rect 11747 16677 11759 16680
rect 11701 16671 11759 16677
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 12176 16640 12204 16748
rect 12360 16708 12388 16748
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 13173 16779 13231 16785
rect 13173 16776 13185 16779
rect 12584 16748 13185 16776
rect 12584 16736 12590 16748
rect 13173 16745 13185 16748
rect 13219 16745 13231 16779
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 13173 16739 13231 16745
rect 13260 16748 16405 16776
rect 13260 16708 13288 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 16850 16736 16856 16788
rect 16908 16736 16914 16788
rect 18046 16736 18052 16788
rect 18104 16736 18110 16788
rect 18782 16736 18788 16788
rect 18840 16736 18846 16788
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19475 16748 19932 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 12360 16680 13288 16708
rect 14182 16668 14188 16720
rect 14240 16708 14246 16720
rect 14642 16708 14648 16720
rect 14240 16680 14648 16708
rect 14240 16668 14246 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 18064 16708 18092 16736
rect 16776 16680 18092 16708
rect 18233 16711 18291 16717
rect 11532 16612 12204 16640
rect 11532 16581 11560 16612
rect 10796 16544 11376 16572
rect 11425 16575 11483 16581
rect 10796 16513 10824 16544
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 10781 16507 10839 16513
rect 10781 16504 10793 16507
rect 9692 16476 10793 16504
rect 9033 16467 9091 16473
rect 10781 16473 10793 16476
rect 10827 16473 10839 16507
rect 10781 16467 10839 16473
rect 10962 16464 10968 16516
rect 11020 16464 11026 16516
rect 6178 16436 6184 16448
rect 5368 16408 6184 16436
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6730 16396 6736 16448
rect 6788 16396 6794 16448
rect 7190 16396 7196 16448
rect 7248 16396 7254 16448
rect 9490 16396 9496 16448
rect 9548 16396 9554 16448
rect 11440 16436 11468 16535
rect 11808 16504 11836 16535
rect 11974 16532 11980 16584
rect 12032 16532 12038 16584
rect 12176 16581 12204 16612
rect 12250 16600 12256 16652
rect 12308 16600 12314 16652
rect 16776 16649 16804 16680
rect 18233 16677 18245 16711
rect 18279 16708 18291 16711
rect 18322 16708 18328 16720
rect 18279 16680 18328 16708
rect 18279 16677 18291 16680
rect 18233 16671 18291 16677
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 18874 16668 18880 16720
rect 18932 16708 18938 16720
rect 19245 16711 19303 16717
rect 19245 16708 19257 16711
rect 18932 16680 19257 16708
rect 18932 16668 18938 16680
rect 19245 16677 19257 16680
rect 19291 16677 19303 16711
rect 19245 16671 19303 16677
rect 16761 16643 16819 16649
rect 12452 16612 12756 16640
rect 12452 16581 12480 16612
rect 12728 16584 12756 16612
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 17819 16612 18460 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 12636 16504 12664 16535
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 16574 16532 16580 16584
rect 16632 16532 16638 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 16724 16544 17877 16572
rect 16724 16532 16730 16544
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 18230 16532 18236 16584
rect 18288 16532 18294 16584
rect 18432 16581 18460 16612
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19150 16640 19156 16652
rect 19024 16612 19156 16640
rect 19024 16600 19030 16612
rect 19150 16600 19156 16612
rect 19208 16640 19214 16652
rect 19518 16640 19524 16652
rect 19208 16612 19524 16640
rect 19208 16600 19214 16612
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 19904 16584 19932 16748
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 20036 16748 20085 16776
rect 20036 16736 20042 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 20533 16779 20591 16785
rect 20533 16745 20545 16779
rect 20579 16776 20591 16779
rect 21082 16776 21088 16788
rect 20579 16748 21088 16776
rect 20579 16745 20591 16748
rect 20533 16739 20591 16745
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 22462 16736 22468 16788
rect 22520 16776 22526 16788
rect 22833 16779 22891 16785
rect 22833 16776 22845 16779
rect 22520 16748 22845 16776
rect 22520 16736 22526 16748
rect 22833 16745 22845 16748
rect 22879 16745 22891 16779
rect 22833 16739 22891 16745
rect 23198 16736 23204 16788
rect 23256 16736 23262 16788
rect 23382 16736 23388 16788
rect 23440 16736 23446 16788
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 24029 16779 24087 16785
rect 24029 16776 24041 16779
rect 23808 16748 24041 16776
rect 23808 16736 23814 16748
rect 24029 16745 24041 16748
rect 24075 16745 24087 16779
rect 24029 16739 24087 16745
rect 25317 16779 25375 16785
rect 25317 16745 25329 16779
rect 25363 16776 25375 16779
rect 25590 16776 25596 16788
rect 25363 16748 25596 16776
rect 25363 16745 25375 16748
rect 25317 16739 25375 16745
rect 25590 16736 25596 16748
rect 25648 16736 25654 16788
rect 21358 16600 21364 16652
rect 21416 16600 21422 16652
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16572 18659 16575
rect 18690 16572 18696 16584
rect 18647 16544 18696 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 19628 16544 19840 16572
rect 11808 16476 12664 16504
rect 12452 16448 12480 16476
rect 12802 16464 12808 16516
rect 12860 16464 12866 16516
rect 12989 16507 13047 16513
rect 12989 16473 13001 16507
rect 13035 16473 13047 16507
rect 12989 16467 13047 16473
rect 11974 16436 11980 16448
rect 11440 16408 11980 16436
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 13004 16436 13032 16467
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 13320 16476 14688 16504
rect 13320 16464 13326 16476
rect 12492 16408 13032 16436
rect 12492 16396 12498 16408
rect 14182 16396 14188 16448
rect 14240 16396 14246 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14550 16436 14556 16448
rect 14332 16408 14556 16436
rect 14332 16396 14338 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 14660 16436 14688 16476
rect 16850 16464 16856 16516
rect 16908 16464 16914 16516
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16504 17463 16507
rect 17494 16504 17500 16516
rect 17451 16476 17500 16504
rect 17451 16473 17463 16476
rect 17405 16467 17463 16473
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 17589 16507 17647 16513
rect 17589 16473 17601 16507
rect 17635 16504 17647 16507
rect 17954 16504 17960 16516
rect 17635 16476 17960 16504
rect 17635 16473 17647 16476
rect 17589 16467 17647 16473
rect 17954 16464 17960 16476
rect 18012 16504 18018 16516
rect 18248 16504 18276 16532
rect 19444 16504 19472 16532
rect 19628 16513 19656 16544
rect 19812 16516 19840 16544
rect 19886 16532 19892 16584
rect 19944 16532 19950 16584
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 22094 16572 22100 16584
rect 21192 16544 22100 16572
rect 18012 16476 18276 16504
rect 19168 16476 19472 16504
rect 19613 16507 19671 16513
rect 18012 16464 18018 16476
rect 17218 16436 17224 16448
rect 14660 16408 17224 16436
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 17828 16408 18061 16436
rect 17828 16396 17834 16408
rect 18049 16405 18061 16408
rect 18095 16436 18107 16439
rect 18414 16436 18420 16448
rect 18095 16408 18420 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18414 16396 18420 16408
rect 18472 16436 18478 16448
rect 19168 16436 19196 16476
rect 19613 16473 19625 16507
rect 19659 16473 19671 16507
rect 19613 16467 19671 16473
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 19794 16464 19800 16516
rect 19852 16504 19858 16516
rect 20254 16504 20260 16516
rect 19852 16476 20260 16504
rect 19852 16464 19858 16476
rect 20254 16464 20260 16476
rect 20312 16504 20318 16516
rect 20717 16507 20775 16513
rect 20717 16504 20729 16507
rect 20312 16476 20729 16504
rect 20312 16464 20318 16476
rect 20717 16473 20729 16476
rect 20763 16473 20775 16507
rect 20717 16467 20775 16473
rect 19426 16445 19432 16448
rect 18472 16408 19196 16436
rect 19413 16439 19432 16445
rect 18472 16396 18478 16408
rect 19413 16405 19425 16439
rect 19413 16399 19432 16405
rect 19426 16396 19432 16399
rect 19484 16396 19490 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 20530 16445 20536 16448
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 19576 16408 20361 16436
rect 19576 16396 19582 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 20349 16399 20407 16405
rect 20512 16439 20536 16445
rect 20512 16405 20524 16439
rect 20588 16436 20594 16448
rect 21192 16436 21220 16544
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 23012 16575 23070 16581
rect 23012 16541 23024 16575
rect 23058 16572 23070 16575
rect 23216 16572 23244 16736
rect 23400 16708 23428 16736
rect 23058 16544 23244 16572
rect 23308 16680 23428 16708
rect 23058 16541 23070 16544
rect 23012 16535 23070 16541
rect 21606 16507 21664 16513
rect 21606 16504 21618 16507
rect 21284 16476 21618 16504
rect 21284 16445 21312 16476
rect 21606 16473 21618 16476
rect 21652 16473 21664 16507
rect 21606 16467 21664 16473
rect 23109 16507 23167 16513
rect 23109 16473 23121 16507
rect 23155 16473 23167 16507
rect 23109 16467 23167 16473
rect 23201 16507 23259 16513
rect 23201 16473 23213 16507
rect 23247 16504 23259 16507
rect 23308 16504 23336 16680
rect 23842 16668 23848 16720
rect 23900 16668 23906 16720
rect 25130 16668 25136 16720
rect 25188 16668 25194 16720
rect 23400 16612 23612 16640
rect 23400 16581 23428 16612
rect 23384 16575 23442 16581
rect 23384 16541 23396 16575
rect 23430 16541 23442 16575
rect 23384 16535 23442 16541
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 23584 16572 23612 16612
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 24636 16612 25881 16640
rect 24636 16600 24642 16612
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 25869 16603 25927 16609
rect 23584 16544 25820 16572
rect 23247 16476 23336 16504
rect 23247 16473 23259 16476
rect 23201 16467 23259 16473
rect 20588 16408 21220 16436
rect 21269 16439 21327 16445
rect 20512 16399 20536 16405
rect 20530 16396 20536 16399
rect 20588 16396 20594 16408
rect 21269 16405 21281 16439
rect 21315 16405 21327 16439
rect 21269 16399 21327 16405
rect 22741 16439 22799 16445
rect 22741 16405 22753 16439
rect 22787 16436 22799 16439
rect 23124 16436 23152 16467
rect 23566 16464 23572 16516
rect 23624 16464 23630 16516
rect 23842 16464 23848 16516
rect 23900 16464 23906 16516
rect 24854 16464 24860 16516
rect 24912 16464 24918 16516
rect 23860 16436 23888 16464
rect 22787 16408 23888 16436
rect 25792 16436 25820 16544
rect 27062 16532 27068 16584
rect 27120 16572 27126 16584
rect 27341 16575 27399 16581
rect 27341 16572 27353 16575
rect 27120 16544 27353 16572
rect 27120 16532 27126 16544
rect 27341 16541 27353 16544
rect 27387 16541 27399 16575
rect 27341 16535 27399 16541
rect 26136 16507 26194 16513
rect 26136 16473 26148 16507
rect 26182 16504 26194 16507
rect 26418 16504 26424 16516
rect 26182 16476 26424 16504
rect 26182 16473 26194 16476
rect 26136 16467 26194 16473
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 27154 16436 27160 16448
rect 25792 16408 27160 16436
rect 22787 16405 22799 16408
rect 22741 16399 22799 16405
rect 27154 16396 27160 16408
rect 27212 16436 27218 16448
rect 27249 16439 27307 16445
rect 27249 16436 27261 16439
rect 27212 16408 27261 16436
rect 27212 16396 27218 16408
rect 27249 16405 27261 16408
rect 27295 16405 27307 16439
rect 27249 16399 27307 16405
rect 27522 16396 27528 16448
rect 27580 16396 27586 16448
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 2924 16204 3617 16232
rect 2924 16192 2930 16204
rect 3605 16201 3617 16204
rect 3651 16201 3663 16235
rect 3605 16195 3663 16201
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 3973 16235 4031 16241
rect 3973 16232 3985 16235
rect 3844 16204 3985 16232
rect 3844 16192 3850 16204
rect 3973 16201 3985 16204
rect 4019 16201 4031 16235
rect 3973 16195 4031 16201
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 5810 16232 5816 16244
rect 4120 16204 5816 16232
rect 4120 16192 4126 16204
rect 1670 16124 1676 16176
rect 1728 16124 1734 16176
rect 2958 16124 2964 16176
rect 3016 16164 3022 16176
rect 3016 16136 4844 16164
rect 3016 16124 3022 16136
rect 3804 16108 3832 16136
rect 750 16056 756 16108
rect 808 16096 814 16108
rect 1489 16099 1547 16105
rect 1489 16096 1501 16099
rect 808 16068 1501 16096
rect 808 16056 814 16068
rect 1489 16065 1501 16068
rect 1535 16065 1547 16099
rect 1489 16059 1547 16065
rect 2216 16099 2274 16105
rect 2216 16065 2228 16099
rect 2262 16096 2274 16099
rect 3326 16096 3332 16108
rect 2262 16068 3332 16096
rect 2262 16065 2274 16068
rect 2216 16059 2274 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 3786 16056 3792 16108
rect 3844 16056 3850 16108
rect 4816 16105 4844 16136
rect 4890 16124 4896 16176
rect 4948 16164 4954 16176
rect 4948 16136 5396 16164
rect 4948 16124 4954 16136
rect 5368 16105 5396 16136
rect 5644 16105 5672 16204
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6178 16192 6184 16244
rect 6236 16232 6242 16244
rect 6236 16204 6500 16232
rect 6236 16192 6242 16204
rect 6472 16173 6500 16204
rect 7190 16192 7196 16244
rect 7248 16192 7254 16244
rect 7561 16235 7619 16241
rect 7561 16201 7573 16235
rect 7607 16232 7619 16235
rect 7650 16232 7656 16244
rect 7607 16204 7656 16232
rect 7607 16201 7619 16204
rect 7561 16195 7619 16201
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9398 16232 9404 16244
rect 9355 16204 9404 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11020 16204 11744 16232
rect 11020 16192 11026 16204
rect 6457 16167 6515 16173
rect 6457 16133 6469 16167
rect 6503 16133 6515 16167
rect 7208 16164 7236 16192
rect 8196 16167 8254 16173
rect 7208 16136 8156 16164
rect 6457 16127 6515 16133
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 3988 16068 4721 16096
rect 3988 16040 4016 16068
rect 4709 16065 4721 16068
rect 4755 16065 4767 16099
rect 4709 16059 4767 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6472 16096 6500 16127
rect 6227 16068 6500 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 7156 16068 7297 16096
rect 7156 16056 7162 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 8128 16096 8156 16136
rect 8196 16133 8208 16167
rect 8242 16164 8254 16167
rect 8662 16164 8668 16176
rect 8242 16136 8668 16164
rect 8242 16133 8254 16136
rect 8196 16127 8254 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 11716 16173 11744 16204
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12710 16232 12716 16244
rect 12124 16204 12716 16232
rect 12124 16192 12130 16204
rect 12710 16192 12716 16204
rect 12768 16232 12774 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 12768 16204 13093 16232
rect 12768 16192 12774 16204
rect 13081 16201 13093 16204
rect 13127 16201 13139 16235
rect 13998 16232 14004 16244
rect 13081 16195 13139 16201
rect 13832 16204 14004 16232
rect 11701 16167 11759 16173
rect 9692 16136 11652 16164
rect 9692 16096 9720 16136
rect 9858 16105 9864 16108
rect 8128 16068 9720 16096
rect 7377 16059 7435 16065
rect 9852 16059 9864 16105
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 15997 2007 16031
rect 1949 15991 2007 15997
rect 1964 15892 1992 15991
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3200 16000 3893 16028
rect 3200 15988 3206 16000
rect 3881 15997 3893 16000
rect 3927 16028 3939 16031
rect 3970 16028 3976 16040
rect 3927 16000 3976 16028
rect 3927 15997 3939 16000
rect 3881 15991 3939 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 16028 4307 16031
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 4295 16000 4353 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4341 15997 4353 16000
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 7392 16028 7420 16059
rect 9858 16056 9864 16059
rect 9916 16056 9922 16108
rect 11624 16096 11652 16136
rect 11701 16133 11713 16167
rect 11747 16133 11759 16167
rect 13832 16164 13860 16204
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 14182 16192 14188 16244
rect 14240 16192 14246 16244
rect 14734 16192 14740 16244
rect 14792 16232 14798 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 14792 16204 15301 16232
rect 14792 16192 14798 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16114 16232 16120 16244
rect 15988 16204 16120 16232
rect 15988 16192 15994 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 17034 16232 17040 16244
rect 16224 16204 17040 16232
rect 11701 16127 11759 16133
rect 11808 16136 13860 16164
rect 13900 16167 13958 16173
rect 11808 16096 11836 16136
rect 13900 16133 13912 16167
rect 13946 16164 13958 16167
rect 14200 16164 14228 16192
rect 13946 16136 14228 16164
rect 13946 16133 13958 16136
rect 13900 16127 13958 16133
rect 14274 16124 14280 16176
rect 14332 16164 14338 16176
rect 16224 16164 16252 16204
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 18064 16204 18368 16232
rect 14332 16136 16252 16164
rect 14332 16124 14338 16136
rect 11624 16068 11836 16096
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 12158 16096 12164 16108
rect 11931 16068 12164 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12158 16056 12164 16068
rect 12216 16096 12222 16108
rect 12802 16096 12808 16108
rect 12216 16068 12808 16096
rect 12216 16056 12222 16068
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 15102 16096 15108 16108
rect 13311 16068 15108 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 16114 16096 16120 16108
rect 15243 16068 16120 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16209 16099 16267 16105
rect 16209 16065 16221 16099
rect 16255 16096 16267 16099
rect 16298 16096 16304 16108
rect 16255 16068 16304 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 6963 16000 7420 16028
rect 7929 16031 7987 16037
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7929 15997 7941 16031
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 3329 15963 3387 15969
rect 3329 15929 3341 15963
rect 3375 15960 3387 15963
rect 4264 15960 4292 15991
rect 3375 15932 4292 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 5258 15920 5264 15972
rect 5316 15920 5322 15972
rect 6086 15920 6092 15972
rect 6144 15920 6150 15972
rect 6730 15920 6736 15972
rect 6788 15920 6794 15972
rect 7101 15963 7159 15969
rect 7101 15929 7113 15963
rect 7147 15960 7159 15963
rect 7374 15960 7380 15972
rect 7147 15932 7380 15960
rect 7147 15929 7159 15932
rect 7101 15923 7159 15929
rect 7374 15920 7380 15932
rect 7432 15960 7438 15972
rect 7944 15960 7972 15991
rect 7432 15932 7972 15960
rect 7432 15920 7438 15932
rect 2130 15892 2136 15904
rect 1964 15864 2136 15892
rect 2130 15852 2136 15864
rect 2188 15852 2194 15904
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4396 15864 4537 15892
rect 4396 15852 4402 15864
rect 4525 15861 4537 15864
rect 4571 15861 4583 15895
rect 5276 15892 5304 15920
rect 6748 15892 6776 15920
rect 5276 15864 6776 15892
rect 7944 15892 7972 15932
rect 9600 15892 9628 15991
rect 13188 15960 13216 16056
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 13648 15960 13676 15991
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 15470 16028 15476 16040
rect 14700 16000 15476 16028
rect 14700 15988 14706 16000
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 15565 16031 15623 16037
rect 15565 15997 15577 16031
rect 15611 16028 15623 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15611 16000 15669 16028
rect 15611 15997 15623 16000
rect 15565 15991 15623 15997
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 16224 16028 16252 16059
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 16390 16056 16396 16108
rect 16448 16056 16454 16108
rect 18064 16096 18092 16204
rect 18340 16176 18368 16204
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20346 16232 20352 16244
rect 19760 16204 20352 16232
rect 19760 16192 19766 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 20622 16192 20628 16244
rect 20680 16192 20686 16244
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 21082 16232 21088 16244
rect 20763 16204 21088 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 21358 16192 21364 16244
rect 21416 16232 21422 16244
rect 21634 16232 21640 16244
rect 21416 16204 21640 16232
rect 21416 16192 21422 16204
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 22830 16232 22836 16244
rect 21988 16204 22836 16232
rect 18322 16124 18328 16176
rect 18380 16124 18386 16176
rect 20640 16164 20668 16192
rect 21988 16173 22016 16204
rect 22830 16192 22836 16204
rect 22888 16192 22894 16244
rect 24762 16232 24768 16244
rect 24320 16204 24768 16232
rect 21973 16167 22031 16173
rect 21973 16164 21985 16167
rect 20640 16136 21985 16164
rect 21973 16133 21985 16136
rect 22019 16133 22031 16167
rect 21973 16127 22031 16133
rect 22189 16167 22247 16173
rect 22189 16133 22201 16167
rect 22235 16164 22247 16167
rect 22370 16164 22376 16176
rect 22235 16136 22376 16164
rect 22235 16133 22247 16136
rect 22189 16127 22247 16133
rect 22370 16124 22376 16136
rect 22428 16124 22434 16176
rect 24320 16108 24348 16204
rect 24762 16192 24768 16204
rect 24820 16232 24826 16244
rect 26142 16232 26148 16244
rect 24820 16204 26148 16232
rect 24820 16192 24826 16204
rect 25682 16164 25688 16176
rect 24412 16136 25688 16164
rect 18150 16099 18208 16105
rect 18150 16096 18162 16099
rect 18064 16068 18162 16096
rect 18150 16065 18162 16068
rect 18196 16065 18208 16099
rect 18150 16059 18208 16065
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 18506 16056 18512 16108
rect 18564 16096 18570 16108
rect 18564 16068 19656 16096
rect 18564 16056 18570 16068
rect 15657 15991 15715 15997
rect 16040 16000 16252 16028
rect 16040 15960 16068 16000
rect 19518 15988 19524 16040
rect 19576 15988 19582 16040
rect 19628 16028 19656 16068
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 20438 16056 20444 16108
rect 20496 16096 20502 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20496 16068 20545 16096
rect 20496 16056 20502 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 21048 16068 21097 16096
rect 21048 16056 21054 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 24302 16096 24308 16108
rect 21085 16059 21143 16065
rect 21192 16068 24308 16096
rect 21192 16028 21220 16068
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 24412 16028 24440 16136
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 25976 16173 26004 16204
rect 26142 16192 26148 16204
rect 26200 16192 26206 16244
rect 26418 16192 26424 16244
rect 26476 16192 26482 16244
rect 27522 16192 27528 16244
rect 27580 16192 27586 16244
rect 25961 16167 26019 16173
rect 25961 16133 25973 16167
rect 26007 16133 26019 16167
rect 25961 16127 26019 16133
rect 27424 16167 27482 16173
rect 27424 16133 27436 16167
rect 27470 16164 27482 16167
rect 27540 16164 27568 16192
rect 27470 16136 27568 16164
rect 27470 16133 27482 16136
rect 27424 16127 27482 16133
rect 24489 16099 24547 16105
rect 24489 16065 24501 16099
rect 24535 16096 24547 16099
rect 24578 16096 24584 16108
rect 24535 16068 24584 16096
rect 24535 16065 24547 16068
rect 24489 16059 24547 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 24762 16105 24768 16108
rect 24756 16059 24768 16105
rect 24762 16056 24768 16059
rect 24820 16056 24826 16108
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16096 26387 16099
rect 26605 16099 26663 16105
rect 26605 16096 26617 16099
rect 26375 16068 26617 16096
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 26605 16065 26617 16068
rect 26651 16065 26663 16099
rect 26605 16059 26663 16065
rect 26160 16028 26188 16059
rect 26970 16056 26976 16108
rect 27028 16096 27034 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 27028 16068 27169 16096
rect 27028 16056 27034 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 19628 16000 21220 16028
rect 22020 16000 24440 16028
rect 25792 16000 26188 16028
rect 10520 15932 13676 15960
rect 14844 15932 16068 15960
rect 16117 15963 16175 15969
rect 10520 15892 10548 15932
rect 7944 15864 10548 15892
rect 4525 15855 4583 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11296 15864 11529 15892
rect 11296 15852 11302 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 14844 15892 14872 15932
rect 16117 15929 16129 15963
rect 16163 15960 16175 15963
rect 16163 15932 17540 15960
rect 16163 15929 16175 15932
rect 16117 15923 16175 15929
rect 13136 15864 14872 15892
rect 13136 15852 13142 15864
rect 15010 15852 15016 15904
rect 15068 15852 15074 15904
rect 15378 15852 15384 15904
rect 15436 15852 15442 15904
rect 15470 15852 15476 15904
rect 15528 15852 15534 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 15933 15895 15991 15901
rect 15933 15892 15945 15895
rect 15620 15864 15945 15892
rect 15620 15852 15626 15864
rect 15933 15861 15945 15864
rect 15979 15861 15991 15895
rect 15933 15855 15991 15861
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 17402 15892 17408 15904
rect 16071 15864 17408 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17512 15892 17540 15932
rect 19536 15892 19564 15988
rect 17512 15864 19564 15892
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20772 15864 21005 15892
rect 20772 15852 20778 15864
rect 20993 15861 21005 15864
rect 21039 15892 21051 15895
rect 21082 15892 21088 15904
rect 21039 15864 21088 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 21818 15852 21824 15904
rect 21876 15852 21882 15904
rect 22020 15901 22048 16000
rect 23198 15920 23204 15972
rect 23256 15960 23262 15972
rect 24118 15960 24124 15972
rect 23256 15932 24124 15960
rect 23256 15920 23262 15932
rect 24118 15920 24124 15932
rect 24176 15920 24182 15972
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 25792 15892 25820 16000
rect 23164 15864 25820 15892
rect 23164 15852 23170 15864
rect 25866 15852 25872 15904
rect 25924 15852 25930 15904
rect 26160 15892 26188 16000
rect 28537 15895 28595 15901
rect 28537 15892 28549 15895
rect 26160 15864 28549 15892
rect 28537 15861 28549 15864
rect 28583 15861 28595 15895
rect 28537 15855 28595 15861
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 3384 15660 3893 15688
rect 3384 15648 3390 15660
rect 3881 15657 3893 15660
rect 3927 15657 3939 15691
rect 3881 15651 3939 15657
rect 4338 15648 4344 15700
rect 4396 15648 4402 15700
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 9490 15648 9496 15700
rect 9548 15648 9554 15700
rect 9769 15691 9827 15697
rect 9769 15657 9781 15691
rect 9815 15688 9827 15691
rect 9858 15688 9864 15700
rect 9815 15660 9864 15688
rect 9815 15657 9827 15660
rect 9769 15651 9827 15657
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10502 15648 10508 15700
rect 10560 15688 10566 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10560 15660 10793 15688
rect 10560 15648 10566 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 12434 15648 12440 15700
rect 12492 15648 12498 15700
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 13630 15688 13636 15700
rect 12768 15660 13636 15688
rect 12768 15648 12774 15660
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14424 15660 14657 15688
rect 14424 15648 14430 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 15749 15691 15807 15697
rect 15749 15688 15761 15691
rect 14645 15651 14703 15657
rect 15028 15660 15761 15688
rect 4154 15620 4160 15632
rect 2240 15592 4160 15620
rect 2240 15496 2268 15592
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 3559 15555 3617 15561
rect 3559 15521 3571 15555
rect 3605 15552 3617 15555
rect 3605 15524 4292 15552
rect 3605 15521 3617 15524
rect 3559 15515 3617 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1811 15456 1869 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 2222 15444 2228 15496
rect 2280 15444 2286 15496
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 3456 15484 3514 15487
rect 3292 15481 3514 15484
rect 3292 15456 3468 15481
rect 3292 15444 3298 15456
rect 3436 15450 3468 15456
rect 3456 15447 3468 15450
rect 3502 15447 3514 15481
rect 3456 15441 3514 15447
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4264 15493 4292 15524
rect 4356 15493 4384 15648
rect 4816 15620 4844 15648
rect 4540 15592 4844 15620
rect 4540 15493 4568 15592
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5718 15552 5724 15564
rect 4847 15524 5724 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5718 15512 5724 15524
rect 5776 15552 5782 15564
rect 5994 15552 6000 15564
rect 5776 15524 6000 15552
rect 5776 15512 5782 15524
rect 5994 15512 6000 15524
rect 6052 15552 6058 15564
rect 6089 15555 6147 15561
rect 6089 15552 6101 15555
rect 6052 15524 6101 15552
rect 6052 15512 6058 15524
rect 6089 15521 6101 15524
rect 6135 15521 6147 15555
rect 9306 15552 9312 15564
rect 6089 15515 6147 15521
rect 7668 15524 9312 15552
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 3844 15456 4077 15484
rect 3844 15444 3850 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4982 15444 4988 15496
rect 5040 15444 5046 15496
rect 7668 15493 7696 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 3970 15376 3976 15428
rect 4028 15416 4034 15428
rect 4154 15416 4160 15428
rect 4028 15388 4160 15416
rect 4028 15376 4034 15388
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 8404 15416 8432 15447
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9508 15484 9536 15648
rect 15028 15632 15056 15660
rect 15749 15657 15761 15660
rect 15795 15657 15807 15691
rect 15749 15651 15807 15657
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 16209 15691 16267 15697
rect 16209 15688 16221 15691
rect 15988 15660 16221 15688
rect 15988 15648 15994 15660
rect 16209 15657 16221 15660
rect 16255 15657 16267 15691
rect 16209 15651 16267 15657
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 17092 15660 17448 15688
rect 17092 15648 17098 15660
rect 13078 15580 13084 15632
rect 13136 15580 13142 15632
rect 15010 15620 15016 15632
rect 14384 15592 15016 15620
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13354 15552 13360 15564
rect 12952 15524 13360 15552
rect 12952 15512 12958 15524
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9508 15456 9597 15484
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 11072 15456 13461 15484
rect 11072 15416 11100 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 14274 15484 14280 15496
rect 13679 15456 14280 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 14384 15493 14412 15592
rect 15010 15580 15016 15592
rect 15068 15580 15074 15632
rect 15102 15580 15108 15632
rect 15160 15580 15166 15632
rect 16114 15580 16120 15632
rect 16172 15620 16178 15632
rect 17313 15623 17371 15629
rect 17313 15620 17325 15623
rect 16172 15592 17325 15620
rect 16172 15580 16178 15592
rect 17313 15589 17325 15592
rect 17359 15589 17371 15623
rect 17313 15583 17371 15589
rect 16298 15552 16304 15564
rect 15580 15524 16304 15552
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 14918 15484 14924 15496
rect 14875 15456 14924 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15286 15460 15292 15512
rect 15344 15500 15350 15512
rect 15344 15484 15424 15500
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15344 15472 15485 15484
rect 15344 15460 15350 15472
rect 15396 15456 15485 15472
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 8404 15388 11100 15416
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 11302 15419 11360 15425
rect 11302 15416 11314 15419
rect 11204 15388 11314 15416
rect 11204 15376 11210 15388
rect 11302 15385 11314 15388
rect 11348 15385 11360 15419
rect 11302 15379 11360 15385
rect 12406 15388 13308 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1670 15348 1676 15360
rect 1627 15320 1676 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 5718 15348 5724 15360
rect 5583 15320 5724 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 7432 15320 7481 15348
rect 7432 15308 7438 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8294 15348 8300 15360
rect 8251 15320 8300 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 12406 15348 12434 15388
rect 9364 15320 12434 15348
rect 9364 15308 9370 15320
rect 12894 15308 12900 15360
rect 12952 15308 12958 15360
rect 13280 15348 13308 15388
rect 13814 15376 13820 15428
rect 13872 15376 13878 15428
rect 14185 15419 14243 15425
rect 14185 15385 14197 15419
rect 14231 15385 14243 15419
rect 14185 15379 14243 15385
rect 14200 15348 14228 15379
rect 14550 15376 14556 15428
rect 14608 15416 14614 15428
rect 15013 15419 15071 15425
rect 15013 15416 15025 15419
rect 14608 15388 15025 15416
rect 14608 15376 14614 15388
rect 15013 15385 15025 15388
rect 15059 15385 15071 15419
rect 15013 15379 15071 15385
rect 15289 15419 15347 15425
rect 15289 15385 15301 15419
rect 15335 15416 15347 15419
rect 15580 15416 15608 15524
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 16942 15444 16948 15496
rect 17000 15444 17006 15496
rect 17420 15484 17448 15660
rect 17586 15648 17592 15700
rect 17644 15648 17650 15700
rect 17678 15648 17684 15700
rect 17736 15648 17742 15700
rect 17773 15691 17831 15697
rect 17773 15657 17785 15691
rect 17819 15688 17831 15691
rect 21818 15688 21824 15700
rect 17819 15660 21824 15688
rect 17819 15657 17831 15660
rect 17773 15651 17831 15657
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 23106 15648 23112 15700
rect 23164 15648 23170 15700
rect 23937 15691 23995 15697
rect 23937 15657 23949 15691
rect 23983 15657 23995 15691
rect 23937 15651 23995 15657
rect 18046 15620 18052 15632
rect 17972 15592 18052 15620
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17420 15456 17877 15484
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 15335 15388 15608 15416
rect 15335 15385 15347 15388
rect 15289 15379 15347 15385
rect 15930 15376 15936 15428
rect 15988 15376 15994 15428
rect 16025 15419 16083 15425
rect 16025 15385 16037 15419
rect 16071 15416 16083 15419
rect 16960 15416 16988 15444
rect 17218 15416 17224 15428
rect 16071 15388 17224 15416
rect 16071 15385 16083 15388
rect 16025 15379 16083 15385
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 17972 15416 18000 15592
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 20530 15580 20536 15632
rect 20588 15620 20594 15632
rect 22925 15623 22983 15629
rect 22925 15620 22937 15623
rect 20588 15592 22937 15620
rect 20588 15580 20594 15592
rect 22925 15589 22937 15592
rect 22971 15589 22983 15623
rect 22925 15583 22983 15589
rect 23750 15580 23756 15632
rect 23808 15580 23814 15632
rect 23952 15620 23980 15651
rect 24302 15648 24308 15700
rect 24360 15688 24366 15700
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 24360 15660 24593 15688
rect 24360 15648 24366 15660
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 24762 15648 24768 15700
rect 24820 15648 24826 15700
rect 25682 15648 25688 15700
rect 25740 15688 25746 15700
rect 27065 15691 27123 15697
rect 27065 15688 27077 15691
rect 25740 15660 27077 15688
rect 25740 15648 25746 15660
rect 27065 15657 27077 15660
rect 27111 15657 27123 15691
rect 27065 15651 27123 15657
rect 25130 15620 25136 15632
rect 23952 15592 25136 15620
rect 25130 15580 25136 15592
rect 25188 15620 25194 15632
rect 25866 15620 25872 15632
rect 25188 15592 25872 15620
rect 25188 15580 25194 15592
rect 25866 15580 25872 15592
rect 25924 15580 25930 15632
rect 18230 15552 18236 15564
rect 18064 15524 18236 15552
rect 18064 15493 18092 15524
rect 18230 15512 18236 15524
rect 18288 15552 18294 15564
rect 18288 15524 19104 15552
rect 18288 15512 18294 15524
rect 19076 15496 19104 15524
rect 20548 15524 24072 15552
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18555 15456 18613 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18601 15453 18613 15456
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 19058 15444 19064 15496
rect 19116 15444 19122 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19208 15456 19257 15484
rect 19208 15444 19214 15456
rect 19245 15453 19257 15456
rect 19291 15484 19303 15487
rect 20548 15484 20576 15524
rect 19291 15456 20576 15484
rect 19291 15453 19303 15456
rect 19245 15447 19303 15453
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 20680 15456 20944 15484
rect 20680 15444 20686 15456
rect 18141 15419 18199 15425
rect 18141 15416 18153 15419
rect 17644 15388 18153 15416
rect 17644 15376 17650 15388
rect 18141 15385 18153 15388
rect 18187 15385 18199 15419
rect 18141 15379 18199 15385
rect 18322 15376 18328 15428
rect 18380 15376 18386 15428
rect 20916 15425 20944 15456
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21177 15487 21235 15493
rect 21177 15484 21189 15487
rect 21140 15456 21189 15484
rect 21140 15444 21146 15456
rect 21177 15453 21189 15456
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 22756 15493 22784 15524
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 21324 15456 21373 15484
rect 21324 15444 21330 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 21591 15456 21741 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 24044 15428 24072 15524
rect 24397 15487 24455 15493
rect 24397 15453 24409 15487
rect 24443 15484 24455 15487
rect 24762 15484 24768 15496
rect 24443 15456 24768 15484
rect 24443 15453 24455 15456
rect 24397 15447 24455 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 24946 15444 24952 15496
rect 25004 15444 25010 15496
rect 28442 15444 28448 15496
rect 28500 15444 28506 15496
rect 19490 15419 19548 15425
rect 19490 15416 19502 15419
rect 18800 15388 19502 15416
rect 13280 15320 14228 15348
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 15733 15351 15791 15357
rect 15733 15317 15745 15351
rect 15779 15348 15791 15351
rect 16114 15348 16120 15360
rect 15779 15320 16120 15348
rect 15779 15317 15791 15320
rect 15733 15311 15791 15317
rect 16114 15308 16120 15320
rect 16172 15348 16178 15360
rect 16225 15351 16283 15357
rect 16225 15348 16237 15351
rect 16172 15320 16237 15348
rect 16172 15308 16178 15320
rect 16225 15317 16237 15320
rect 16271 15317 16283 15351
rect 16225 15311 16283 15317
rect 16393 15351 16451 15357
rect 16393 15317 16405 15351
rect 16439 15348 16451 15351
rect 16942 15348 16948 15360
rect 16439 15320 16948 15348
rect 16439 15317 16451 15320
rect 16393 15311 16451 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18598 15348 18604 15360
rect 17460 15320 18604 15348
rect 17460 15308 17466 15320
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 18800 15357 18828 15388
rect 19490 15385 19502 15388
rect 19536 15385 19548 15419
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 19490 15379 19548 15385
rect 20364 15388 20729 15416
rect 20364 15360 20392 15388
rect 20717 15385 20729 15388
rect 20763 15385 20775 15419
rect 20717 15379 20775 15385
rect 20901 15419 20959 15425
rect 20901 15385 20913 15419
rect 20947 15416 20959 15419
rect 20990 15416 20996 15428
rect 20947 15388 20996 15416
rect 20947 15385 20959 15388
rect 20901 15379 20959 15385
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22922 15416 22928 15428
rect 22244 15388 22928 15416
rect 22244 15376 22250 15388
rect 22922 15376 22928 15388
rect 22980 15416 22986 15428
rect 23293 15419 23351 15425
rect 23293 15416 23305 15419
rect 22980 15388 23305 15416
rect 22980 15376 22986 15388
rect 23293 15385 23305 15388
rect 23339 15385 23351 15419
rect 23293 15379 23351 15385
rect 24026 15376 24032 15428
rect 24084 15376 24090 15428
rect 24118 15376 24124 15428
rect 24176 15376 24182 15428
rect 27430 15376 27436 15428
rect 27488 15416 27494 15428
rect 28178 15419 28236 15425
rect 28178 15416 28190 15419
rect 27488 15388 28190 15416
rect 27488 15376 27494 15388
rect 28178 15385 28190 15388
rect 28224 15385 28236 15419
rect 28178 15379 28236 15385
rect 18785 15351 18843 15357
rect 18785 15317 18797 15351
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 20346 15308 20352 15360
rect 20404 15308 20410 15360
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 20496 15320 20637 15348
rect 20496 15308 20502 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 20625 15311 20683 15317
rect 21634 15308 21640 15360
rect 21692 15348 21698 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21692 15320 21925 15348
rect 21692 15308 21698 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 22554 15308 22560 15360
rect 22612 15348 22618 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22612 15320 22661 15348
rect 22612 15308 22618 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 22830 15308 22836 15360
rect 22888 15348 22894 15360
rect 23083 15351 23141 15357
rect 23083 15348 23095 15351
rect 22888 15320 23095 15348
rect 22888 15308 22894 15320
rect 23083 15317 23095 15320
rect 23129 15348 23141 15351
rect 23382 15348 23388 15360
rect 23129 15320 23388 15348
rect 23129 15317 23141 15320
rect 23083 15311 23141 15317
rect 23382 15308 23388 15320
rect 23440 15348 23446 15360
rect 23911 15351 23969 15357
rect 23911 15348 23923 15351
rect 23440 15320 23923 15348
rect 23440 15308 23446 15320
rect 23911 15317 23923 15320
rect 23957 15317 23969 15351
rect 23911 15311 23969 15317
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 5442 15144 5448 15156
rect 4172 15116 5448 15144
rect 1670 15085 1676 15088
rect 1664 15039 1676 15085
rect 1728 15076 1734 15088
rect 4172 15076 4200 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5626 15104 5632 15156
rect 5684 15104 5690 15156
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6089 15147 6147 15153
rect 6089 15144 6101 15147
rect 6052 15116 6101 15144
rect 6052 15104 6058 15116
rect 6089 15113 6101 15116
rect 6135 15113 6147 15147
rect 6089 15107 6147 15113
rect 7742 15104 7748 15156
rect 7800 15104 7806 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8352 15116 8432 15144
rect 8352 15104 8358 15116
rect 4798 15076 4804 15088
rect 1728 15048 1764 15076
rect 3068 15048 4200 15076
rect 1670 15036 1676 15039
rect 1728 15036 1734 15048
rect 3068 15017 3096 15048
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 14977 3295 15011
rect 3237 14971 3295 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 3252 14940 3280 14971
rect 3326 14968 3332 15020
rect 3384 14968 3390 15020
rect 4172 15017 4200 15048
rect 4724 15048 4804 15076
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4396 14980 4445 15008
rect 4396 14968 4402 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4614 14968 4620 15020
rect 4672 14968 4678 15020
rect 4724 15017 4752 15048
rect 4798 15036 4804 15048
rect 4856 15076 4862 15088
rect 5644 15076 5672 15104
rect 8404 15085 8432 15116
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 9456 15116 9597 15144
rect 9456 15104 9462 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 11146 15104 11152 15156
rect 11204 15104 11210 15156
rect 11238 15104 11244 15156
rect 11296 15104 11302 15156
rect 12434 15104 12440 15156
rect 12492 15104 12498 15156
rect 12894 15104 12900 15156
rect 12952 15104 12958 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14608 15116 14657 15144
rect 14608 15104 14614 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 15746 15104 15752 15156
rect 15804 15104 15810 15156
rect 17770 15144 17776 15156
rect 16592 15116 17776 15144
rect 4856 15048 5672 15076
rect 4856 15036 4862 15048
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 14977 4767 15011
rect 4965 15011 5023 15017
rect 4965 15008 4977 15011
rect 4709 14971 4767 14977
rect 4816 14980 4977 15008
rect 3510 14940 3516 14952
rect 3252 14912 3516 14940
rect 1397 14903 1455 14909
rect 1412 14804 1440 14903
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 4816 14940 4844 14980
rect 4965 14977 4977 14980
rect 5011 14977 5023 15011
rect 5644 15008 5672 15048
rect 8380 15079 8438 15085
rect 8380 15045 8392 15079
rect 8426 15045 8438 15079
rect 8380 15039 8438 15045
rect 5644 14980 5764 15008
rect 4965 14971 5023 14977
rect 4448 14912 4844 14940
rect 5736 14940 5764 14980
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6144 14980 6653 15008
rect 6144 14968 6150 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 11256 15008 11284 15104
rect 12253 15079 12311 15085
rect 12253 15076 12265 15079
rect 11716 15048 12265 15076
rect 11716 15020 11744 15048
rect 12253 15045 12265 15048
rect 12299 15045 12311 15079
rect 12253 15039 12311 15045
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 11256 14980 11345 15008
rect 11333 14977 11345 14980
rect 11379 14977 11391 15011
rect 11333 14971 11391 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 14977 12127 15011
rect 12912 15008 12940 15104
rect 13814 15036 13820 15088
rect 13872 15036 13878 15088
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12912 14980 13001 15008
rect 12069 14971 12127 14977
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5736 14912 6377 14940
rect 4448 14881 4476 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 8110 14940 8116 14952
rect 7156 14912 8116 14940
rect 7156 14900 7162 14912
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 12084 14940 12112 14971
rect 13832 14940 13860 15036
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 14056 14980 14841 15008
rect 14056 14968 14062 14980
rect 14829 14977 14841 14980
rect 14875 14977 14887 15011
rect 15764 15008 15792 15104
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 15764 14980 16313 15008
rect 14829 14971 14887 14977
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 11204 14912 13860 14940
rect 14844 14940 14872 14971
rect 16592 14940 16620 15116
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18322 15144 18328 15156
rect 18104 15116 18328 15144
rect 18104 15104 18110 15116
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 20272 15116 21128 15144
rect 20272 15088 20300 15116
rect 20254 15036 20260 15088
rect 20312 15036 20318 15088
rect 21100 15085 21128 15116
rect 21726 15104 21732 15156
rect 21784 15144 21790 15156
rect 21784 15116 24900 15144
rect 21784 15104 21790 15116
rect 24872 15088 24900 15116
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 27430 15104 27436 15156
rect 27488 15104 27494 15156
rect 20885 15079 20943 15085
rect 20885 15045 20897 15079
rect 20931 15076 20943 15079
rect 21085 15079 21143 15085
rect 20931 15045 20944 15076
rect 20885 15039 20944 15045
rect 21085 15045 21097 15079
rect 21131 15045 21143 15079
rect 21085 15039 21143 15045
rect 16925 15011 16983 15017
rect 16925 14977 16937 15011
rect 16971 15008 16983 15011
rect 17310 15008 17316 15020
rect 16971 14980 17316 15008
rect 16971 14977 16983 14980
rect 16925 14971 16983 14977
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 17696 15006 18000 15008
rect 18064 15006 20177 15008
rect 17696 14980 20177 15006
rect 14844 14912 16620 14940
rect 16669 14943 16727 14949
rect 11204 14900 11210 14912
rect 16669 14909 16681 14943
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 4433 14875 4491 14881
rect 4433 14841 4445 14875
rect 4479 14841 4491 14875
rect 9677 14875 9735 14881
rect 9677 14872 9689 14875
rect 4433 14835 4491 14841
rect 9508 14844 9689 14872
rect 2130 14804 2136 14816
rect 1412 14776 2136 14804
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 2777 14807 2835 14813
rect 2777 14804 2789 14807
rect 2740 14776 2789 14804
rect 2740 14764 2746 14776
rect 2777 14773 2789 14776
rect 2823 14773 2835 14807
rect 2777 14767 2835 14773
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9508 14813 9536 14844
rect 9677 14841 9689 14844
rect 9723 14841 9735 14875
rect 9677 14835 9735 14841
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 15746 14872 15752 14884
rect 12032 14844 15752 14872
rect 12032 14832 12038 14844
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 9493 14807 9551 14813
rect 9493 14804 9505 14807
rect 9364 14776 9505 14804
rect 9364 14764 9370 14776
rect 9493 14773 9505 14776
rect 9539 14773 9551 14807
rect 9493 14767 9551 14773
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 12802 14764 12808 14816
rect 12860 14764 12866 14816
rect 16485 14807 16543 14813
rect 16485 14773 16497 14807
rect 16531 14804 16543 14807
rect 16574 14804 16580 14816
rect 16531 14776 16580 14804
rect 16531 14773 16543 14776
rect 16485 14767 16543 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 16684 14804 16712 14903
rect 17696 14884 17724 14980
rect 17972 14978 18092 14980
rect 20165 14977 20177 14980
rect 20211 14977 20223 15011
rect 20272 15008 20300 15036
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20272 14980 20361 15008
rect 20165 14971 20223 14977
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20916 15008 20944 15039
rect 21634 15036 21640 15088
rect 21692 15076 21698 15088
rect 22158 15079 22216 15085
rect 22158 15076 22170 15079
rect 21692 15048 22170 15076
rect 21692 15036 21698 15048
rect 22158 15045 22170 15048
rect 22204 15045 22216 15079
rect 22158 15039 22216 15045
rect 23492 15048 24808 15076
rect 21358 15008 21364 15020
rect 20916 14980 21364 15008
rect 20349 14971 20407 14977
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 21913 15011 21971 15017
rect 21913 14977 21925 15011
rect 21959 15008 21971 15011
rect 22554 15008 22560 15020
rect 21959 14980 22560 15008
rect 21959 14977 21971 14980
rect 21913 14971 21971 14977
rect 22554 14968 22560 14980
rect 22612 15008 22618 15020
rect 23492 15017 23520 15048
rect 23750 15017 23756 15020
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 22612 14980 23489 15008
rect 22612 14968 22618 14980
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 23744 14971 23756 15017
rect 23750 14968 23756 14971
rect 23808 14968 23814 15020
rect 24780 15008 24808 15048
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 25409 15079 25467 15085
rect 25409 15076 25421 15079
rect 24912 15048 25421 15076
rect 24912 15036 24918 15048
rect 25409 15045 25421 15048
rect 25455 15045 25467 15079
rect 25409 15039 25467 15045
rect 26145 15011 26203 15017
rect 24780 14980 26004 15008
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 20254 14940 20260 14952
rect 17920 14912 20260 14940
rect 17920 14900 17926 14912
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 21634 14940 21640 14952
rect 20864 14912 21640 14940
rect 20864 14900 20870 14912
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 25590 14900 25596 14952
rect 25648 14900 25654 14952
rect 17678 14832 17684 14884
rect 17736 14832 17742 14884
rect 17770 14832 17776 14884
rect 17828 14872 17834 14884
rect 20622 14872 20628 14884
rect 17828 14844 20628 14872
rect 17828 14832 17834 14844
rect 20622 14832 20628 14844
rect 20680 14832 20686 14884
rect 20990 14832 20996 14884
rect 21048 14872 21054 14884
rect 21450 14872 21456 14884
rect 21048 14844 21456 14872
rect 21048 14832 21054 14844
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 25041 14875 25099 14881
rect 25041 14872 25053 14875
rect 24872 14844 25053 14872
rect 24872 14816 24900 14844
rect 25041 14841 25053 14844
rect 25087 14841 25099 14875
rect 25041 14835 25099 14841
rect 25682 14832 25688 14884
rect 25740 14872 25746 14884
rect 25869 14875 25927 14881
rect 25869 14872 25881 14875
rect 25740 14844 25881 14872
rect 25740 14832 25746 14844
rect 25869 14841 25881 14844
rect 25915 14841 25927 14875
rect 25976 14872 26004 14980
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26053 14943 26111 14949
rect 26053 14909 26065 14943
rect 26099 14940 26111 14943
rect 26160 14940 26188 14971
rect 27246 14968 27252 15020
rect 27304 14968 27310 15020
rect 26099 14912 26188 14940
rect 26099 14909 26111 14912
rect 26053 14903 26111 14909
rect 26970 14872 26976 14884
rect 25976 14844 26976 14872
rect 25869 14835 25927 14841
rect 26970 14832 26976 14844
rect 27028 14832 27034 14884
rect 19150 14804 19156 14816
rect 16684 14776 19156 14804
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 19978 14764 19984 14816
rect 20036 14764 20042 14816
rect 20714 14764 20720 14816
rect 20772 14764 20778 14816
rect 20901 14807 20959 14813
rect 20901 14773 20913 14807
rect 20947 14804 20959 14807
rect 21266 14804 21272 14816
rect 20947 14776 21272 14804
rect 20947 14773 20959 14776
rect 20901 14767 20959 14773
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 23293 14807 23351 14813
rect 23293 14773 23305 14807
rect 23339 14804 23351 14807
rect 23474 14804 23480 14816
rect 23339 14776 23480 14804
rect 23339 14773 23351 14776
rect 23293 14767 23351 14773
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 24854 14764 24860 14816
rect 24912 14764 24918 14816
rect 26326 14764 26332 14816
rect 26384 14764 26390 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1857 14603 1915 14609
rect 1857 14569 1869 14603
rect 1903 14600 1915 14603
rect 2498 14600 2504 14612
rect 1903 14572 2504 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 2498 14560 2504 14572
rect 2556 14600 2562 14612
rect 3142 14600 3148 14612
rect 2556 14572 3148 14600
rect 2556 14560 2562 14572
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3384 14572 3801 14600
rect 3384 14560 3390 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4801 14603 4859 14609
rect 4801 14600 4813 14603
rect 4396 14572 4813 14600
rect 4396 14560 4402 14572
rect 4801 14569 4813 14572
rect 4847 14569 4859 14603
rect 4801 14563 4859 14569
rect 5350 14560 5356 14612
rect 5408 14560 5414 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 15470 14600 15476 14612
rect 13596 14572 15476 14600
rect 13596 14560 13602 14572
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 17310 14600 17316 14612
rect 15795 14572 17316 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17405 14603 17463 14609
rect 17405 14569 17417 14603
rect 17451 14600 17463 14603
rect 18046 14600 18052 14612
rect 17451 14572 18052 14600
rect 17451 14569 17463 14572
rect 17405 14563 17463 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19702 14560 19708 14612
rect 19760 14600 19766 14612
rect 19981 14603 20039 14609
rect 19981 14600 19993 14603
rect 19760 14572 19993 14600
rect 19760 14560 19766 14572
rect 19981 14569 19993 14572
rect 20027 14600 20039 14603
rect 20162 14600 20168 14612
rect 20027 14572 20168 14600
rect 20027 14569 20039 14572
rect 19981 14563 20039 14569
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 22186 14600 22192 14612
rect 20364 14572 22192 14600
rect 4246 14532 4252 14544
rect 4089 14504 4252 14532
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 4089 14473 4117 14504
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 4982 14492 4988 14544
rect 5040 14492 5046 14544
rect 17586 14532 17592 14544
rect 14384 14504 17592 14532
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3476 14436 4077 14464
rect 3476 14424 3482 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 5000 14464 5028 14492
rect 14384 14476 14412 14504
rect 4816 14436 5028 14464
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 2866 14396 2872 14408
rect 2746 14368 2872 14396
rect 1949 14331 2007 14337
rect 1949 14297 1961 14331
rect 1995 14297 2007 14331
rect 1949 14291 2007 14297
rect 2400 14331 2458 14337
rect 2400 14297 2412 14331
rect 2446 14328 2458 14331
rect 2746 14328 2774 14368
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3970 14396 3976 14408
rect 3068 14368 3976 14396
rect 3068 14340 3096 14368
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4816 14405 4844 14436
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8941 14467 8999 14473
rect 8941 14464 8953 14467
rect 8168 14436 8953 14464
rect 8168 14424 8174 14436
rect 8941 14433 8953 14436
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 14366 14424 14372 14476
rect 14424 14424 14430 14476
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 2446 14300 2774 14328
rect 2446 14297 2458 14300
rect 2400 14291 2458 14297
rect 1964 14260 1992 14291
rect 3050 14288 3056 14340
rect 3108 14288 3114 14340
rect 4264 14328 4292 14359
rect 4890 14328 4896 14340
rect 3528 14300 4896 14328
rect 2682 14260 2688 14272
rect 1964 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 3528 14269 3556 14300
rect 4890 14288 4896 14300
rect 4948 14288 4954 14340
rect 5000 14328 5028 14359
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 5261 14399 5319 14405
rect 5261 14396 5273 14399
rect 5224 14368 5273 14396
rect 5224 14356 5230 14368
rect 5261 14365 5273 14368
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5718 14356 5724 14408
rect 5776 14356 5782 14408
rect 7098 14356 7104 14408
rect 7156 14356 7162 14408
rect 7374 14405 7380 14408
rect 7368 14396 7380 14405
rect 7335 14368 7380 14396
rect 7368 14359 7380 14368
rect 7374 14356 7380 14359
rect 7432 14356 7438 14408
rect 9214 14405 9220 14408
rect 9208 14396 9220 14405
rect 9175 14368 9220 14396
rect 9208 14359 9220 14368
rect 9214 14356 9220 14359
rect 9272 14356 9278 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10870 14405 10876 14408
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 9824 14368 10609 14396
rect 9824 14356 9830 14368
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10864 14396 10876 14405
rect 10831 14368 10876 14396
rect 10597 14359 10655 14365
rect 10864 14359 10876 14368
rect 5736 14328 5764 14356
rect 5000 14300 5764 14328
rect 10612 14328 10640 14359
rect 10870 14356 10876 14359
rect 10928 14356 10934 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12428 14399 12486 14405
rect 12428 14365 12440 14399
rect 12474 14396 12486 14399
rect 12802 14396 12808 14408
rect 12474 14368 12808 14396
rect 12474 14365 12486 14368
rect 12428 14359 12486 14365
rect 12176 14328 12204 14359
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14200 14368 14841 14396
rect 14200 14340 14228 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 15059 14368 15577 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 12986 14328 12992 14340
rect 10612 14300 12992 14328
rect 12986 14288 12992 14300
rect 13044 14288 13050 14340
rect 14182 14288 14188 14340
rect 14240 14288 14246 14340
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 14645 14331 14703 14337
rect 14645 14328 14657 14331
rect 14424 14300 14657 14328
rect 14424 14288 14430 14300
rect 14645 14297 14657 14300
rect 14691 14297 14703 14331
rect 15289 14331 15347 14337
rect 15289 14328 15301 14331
rect 14645 14291 14703 14297
rect 14752 14300 15301 14328
rect 3513 14263 3571 14269
rect 3513 14260 3525 14263
rect 3016 14232 3525 14260
rect 3016 14220 3022 14232
rect 3513 14229 3525 14232
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 10318 14220 10324 14272
rect 10376 14220 10382 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11756 14232 11989 14260
rect 11756 14220 11762 14232
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 11977 14223 12035 14229
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13541 14263 13599 14269
rect 13541 14260 13553 14263
rect 13228 14232 13553 14260
rect 13228 14220 13234 14232
rect 13541 14229 13553 14232
rect 13587 14229 13599 14263
rect 13541 14223 13599 14229
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14458 14260 14464 14272
rect 13872 14232 14464 14260
rect 13872 14220 13878 14232
rect 14458 14220 14464 14232
rect 14516 14260 14522 14272
rect 14752 14260 14780 14300
rect 15289 14297 15301 14300
rect 15335 14297 15347 14331
rect 15289 14291 15347 14297
rect 15473 14331 15531 14337
rect 15473 14297 15485 14331
rect 15519 14328 15531 14331
rect 15672 14328 15700 14504
rect 17586 14492 17592 14504
rect 17644 14532 17650 14544
rect 17644 14504 17816 14532
rect 17644 14492 17650 14504
rect 16390 14424 16396 14476
rect 16448 14424 16454 14476
rect 17678 14464 17684 14476
rect 17328 14436 17684 14464
rect 16408 14396 16436 14424
rect 17328 14396 17356 14436
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 17788 14464 17816 14504
rect 17862 14464 17868 14476
rect 17788 14436 17868 14464
rect 17788 14396 17816 14436
rect 17862 14424 17868 14436
rect 17920 14464 17926 14476
rect 19518 14464 19524 14476
rect 17920 14436 19524 14464
rect 17920 14424 17926 14436
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 20364 14464 20392 14572
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 23750 14560 23756 14612
rect 23808 14600 23814 14612
rect 23845 14603 23903 14609
rect 23845 14600 23857 14603
rect 23808 14572 23857 14600
rect 23808 14560 23814 14572
rect 23845 14569 23857 14572
rect 23891 14569 23903 14603
rect 23845 14563 23903 14569
rect 27246 14560 27252 14612
rect 27304 14600 27310 14612
rect 27617 14603 27675 14609
rect 27617 14600 27629 14603
rect 27304 14572 27629 14600
rect 27304 14560 27310 14572
rect 27617 14569 27629 14572
rect 27663 14569 27675 14603
rect 27617 14563 27675 14569
rect 23474 14492 23480 14544
rect 23532 14532 23538 14544
rect 23532 14504 23888 14532
rect 23532 14492 23538 14504
rect 19812 14436 20392 14464
rect 23569 14467 23627 14473
rect 16408 14368 17356 14396
rect 15519 14300 15700 14328
rect 17221 14331 17279 14337
rect 15519 14297 15531 14300
rect 15473 14291 15531 14297
rect 17221 14297 17233 14331
rect 17267 14297 17279 14331
rect 17328 14328 17356 14368
rect 17696 14368 17816 14396
rect 18049 14399 18107 14405
rect 17696 14337 17724 14368
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 18095 14368 18153 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 19334 14356 19340 14408
rect 19392 14356 19398 14408
rect 17421 14331 17479 14337
rect 17421 14328 17433 14331
rect 17328 14300 17433 14328
rect 17221 14291 17279 14297
rect 17421 14297 17433 14300
rect 17467 14297 17479 14331
rect 17421 14291 17479 14297
rect 17681 14331 17739 14337
rect 17681 14297 17693 14331
rect 17727 14297 17739 14331
rect 17865 14331 17923 14337
rect 17865 14328 17877 14331
rect 17681 14291 17739 14297
rect 17788 14300 17877 14328
rect 14516 14232 14780 14260
rect 15105 14263 15163 14269
rect 14516 14220 14522 14232
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 15194 14260 15200 14272
rect 15151 14232 15200 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 17236 14260 17264 14291
rect 17788 14272 17816 14300
rect 17865 14297 17877 14300
rect 17911 14297 17923 14331
rect 17865 14291 17923 14297
rect 17310 14260 17316 14272
rect 17236 14232 17316 14260
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17586 14220 17592 14272
rect 17644 14220 17650 14272
rect 17770 14220 17776 14272
rect 17828 14220 17834 14272
rect 18322 14220 18328 14272
rect 18380 14220 18386 14272
rect 19352 14260 19380 14356
rect 19812 14337 19840 14436
rect 23569 14433 23581 14467
rect 23615 14464 23627 14467
rect 23615 14436 23704 14464
rect 23615 14433 23627 14436
rect 23569 14427 23627 14433
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 20220 14368 20453 14396
rect 20220 14356 20226 14368
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 23676 14405 23704 14436
rect 23860 14408 23888 14504
rect 27522 14492 27528 14544
rect 27580 14492 27586 14544
rect 24946 14424 24952 14476
rect 25004 14424 25010 14476
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 23842 14356 23848 14408
rect 23900 14356 23906 14408
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 19797 14331 19855 14337
rect 19797 14297 19809 14331
rect 19843 14297 19855 14331
rect 19797 14291 19855 14297
rect 20257 14331 20315 14337
rect 20257 14297 20269 14331
rect 20303 14328 20315 14331
rect 20346 14328 20352 14340
rect 20303 14300 20352 14328
rect 20303 14297 20315 14300
rect 20257 14291 20315 14297
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 20898 14288 20904 14340
rect 20956 14328 20962 14340
rect 21054 14331 21112 14337
rect 21054 14328 21066 14331
rect 20956 14300 21066 14328
rect 20956 14288 20962 14300
rect 21054 14297 21066 14300
rect 21100 14297 21112 14331
rect 21054 14291 21112 14297
rect 23109 14331 23167 14337
rect 23109 14297 23121 14331
rect 23155 14328 23167 14331
rect 24964 14328 24992 14424
rect 26326 14356 26332 14408
rect 26384 14396 26390 14408
rect 26798 14399 26856 14405
rect 26798 14396 26810 14399
rect 26384 14368 26810 14396
rect 26384 14356 26390 14368
rect 26798 14365 26810 14368
rect 26844 14365 26856 14399
rect 26798 14359 26856 14365
rect 26970 14356 26976 14408
rect 27028 14396 27034 14408
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 27028 14368 27077 14396
rect 27028 14356 27034 14368
rect 27065 14365 27077 14368
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 27157 14331 27215 14337
rect 27157 14328 27169 14331
rect 23155 14300 24992 14328
rect 25608 14300 27169 14328
rect 23155 14297 23167 14300
rect 23109 14291 23167 14297
rect 25608 14272 25636 14300
rect 27157 14297 27169 14300
rect 27203 14328 27215 14331
rect 27338 14328 27344 14340
rect 27203 14300 27344 14328
rect 27203 14297 27215 14300
rect 27157 14291 27215 14297
rect 27338 14288 27344 14300
rect 27396 14288 27402 14340
rect 19997 14263 20055 14269
rect 19997 14260 20009 14263
rect 19352 14232 20009 14260
rect 19997 14229 20009 14232
rect 20043 14229 20055 14263
rect 19997 14223 20055 14229
rect 20162 14220 20168 14272
rect 20220 14220 20226 14272
rect 20622 14220 20628 14272
rect 20680 14220 20686 14272
rect 22186 14220 22192 14272
rect 22244 14220 22250 14272
rect 24857 14263 24915 14269
rect 24857 14229 24869 14263
rect 24903 14260 24915 14263
rect 25590 14260 25596 14272
rect 24903 14232 25596 14260
rect 24903 14229 24915 14232
rect 24857 14223 24915 14229
rect 25590 14220 25596 14232
rect 25648 14220 25654 14272
rect 25682 14220 25688 14272
rect 25740 14220 25746 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 1578 14016 1584 14068
rect 1636 14016 1642 14068
rect 2958 14016 2964 14068
rect 3016 14016 3022 14068
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 3510 14016 3516 14068
rect 3568 14016 3574 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4433 14059 4491 14065
rect 4433 14056 4445 14059
rect 4304 14028 4445 14056
rect 4304 14016 4310 14028
rect 4433 14025 4445 14028
rect 4479 14056 4491 14059
rect 4982 14056 4988 14068
rect 4479 14028 4988 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10686 14056 10692 14068
rect 10459 14028 10692 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12526 14056 12532 14068
rect 12207 14028 12532 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14025 14151 14059
rect 15930 14056 15936 14068
rect 14093 14019 14151 14025
rect 14476 14028 15936 14056
rect 2682 13948 2688 14000
rect 2740 13948 2746 14000
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 3436 13988 3464 14016
rect 4585 13991 4643 13997
rect 4585 13988 4597 13991
rect 2924 13960 3464 13988
rect 3620 13960 4597 13988
rect 2924 13948 2930 13960
rect 3620 13932 3648 13960
rect 4585 13957 4597 13960
rect 4631 13957 4643 13991
rect 4585 13951 4643 13957
rect 4801 13991 4859 13997
rect 4801 13957 4813 13991
rect 4847 13988 4859 13991
rect 6270 13988 6276 14000
rect 4847 13960 6276 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 7561 13991 7619 13997
rect 7561 13957 7573 13991
rect 7607 13988 7619 13991
rect 8754 13988 8760 14000
rect 7607 13960 8760 13988
rect 7607 13957 7619 13960
rect 7561 13951 7619 13957
rect 8754 13948 8760 13960
rect 8812 13988 8818 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8812 13960 8953 13988
rect 8812 13948 8818 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 8941 13951 8999 13957
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 11146 13988 11152 14000
rect 10827 13960 11152 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 750 13880 756 13932
rect 808 13920 814 13932
rect 1397 13923 1455 13929
rect 1397 13920 1409 13923
rect 808 13892 1409 13920
rect 808 13880 814 13892
rect 1397 13889 1409 13892
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 3602 13920 3608 13932
rect 3283 13892 3608 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 4982 13852 4988 13864
rect 4632 13824 4988 13852
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4632 13725 4660 13824
rect 4982 13812 4988 13824
rect 5040 13852 5046 13864
rect 6454 13852 6460 13864
rect 5040 13824 6460 13852
rect 5040 13812 5046 13824
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 8956 13852 8984 13951
rect 11146 13948 11152 13960
rect 11204 13948 11210 14000
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10318 13920 10324 13932
rect 9732 13892 10324 13920
rect 9732 13880 9738 13892
rect 10318 13880 10324 13892
rect 10376 13920 10382 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10376 13892 10609 13920
rect 10376 13880 10382 13892
rect 10597 13889 10609 13892
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 11974 13880 11980 13932
rect 12032 13880 12038 13932
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13596 13892 13645 13920
rect 13596 13880 13602 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13872 13892 13921 13920
rect 13872 13880 13878 13892
rect 13909 13889 13921 13892
rect 13955 13889 13967 13923
rect 13909 13883 13967 13889
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 14108 13920 14136 14019
rect 14182 13948 14188 14000
rect 14240 13988 14246 14000
rect 14476 13997 14504 14028
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16117 14059 16175 14065
rect 16117 14025 16129 14059
rect 16163 14056 16175 14059
rect 17313 14059 17371 14065
rect 17313 14056 17325 14059
rect 16163 14028 17325 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 17313 14025 17325 14028
rect 17359 14056 17371 14059
rect 17770 14056 17776 14068
rect 17359 14028 17776 14056
rect 17359 14025 17371 14028
rect 17313 14019 17371 14025
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 18012 14028 18153 14056
rect 18012 14016 18018 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 18322 14016 18328 14068
rect 18380 14056 18386 14068
rect 18380 14028 18460 14056
rect 18380 14016 18386 14028
rect 14369 13991 14427 13997
rect 14369 13988 14381 13991
rect 14240 13960 14381 13988
rect 14240 13948 14246 13960
rect 14369 13957 14381 13960
rect 14415 13957 14427 13991
rect 14369 13951 14427 13957
rect 14461 13991 14519 13997
rect 14461 13957 14473 13991
rect 14507 13957 14519 13991
rect 18432 13988 18460 14028
rect 19702 14016 19708 14068
rect 19760 14016 19766 14068
rect 20438 14016 20444 14068
rect 20496 14016 20502 14068
rect 20622 14016 20628 14068
rect 20680 14016 20686 14068
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14056 20867 14059
rect 20898 14056 20904 14068
rect 20855 14028 20904 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 22370 14056 22376 14068
rect 21508 14028 22376 14056
rect 21508 14016 21514 14028
rect 18570 13991 18628 13997
rect 18570 13988 18582 13991
rect 14461 13951 14519 13957
rect 14568 13960 18368 13988
rect 18432 13960 18582 13988
rect 14047 13892 14136 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14568 13920 14596 13960
rect 14332 13892 14596 13920
rect 14645 13923 14703 13929
rect 14332 13880 14338 13892
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 14826 13920 14832 13932
rect 14691 13892 14832 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 15010 13929 15016 13932
rect 15004 13883 15016 13929
rect 15010 13880 15016 13883
rect 15068 13880 15074 13932
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 16390 13920 16396 13932
rect 15528 13892 16396 13920
rect 15528 13880 15534 13892
rect 16390 13880 16396 13892
rect 16448 13920 16454 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16448 13892 17417 13920
rect 16448 13880 16454 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17644 13892 17785 13920
rect 17644 13880 17650 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 18230 13880 18236 13932
rect 18288 13880 18294 13932
rect 18340 13920 18368 13960
rect 18570 13957 18582 13960
rect 18616 13957 18628 13991
rect 18570 13951 18628 13957
rect 19978 13948 19984 14000
rect 20036 13988 20042 14000
rect 20036 13960 20576 13988
rect 20036 13948 20042 13960
rect 20088 13920 20116 13960
rect 18340 13892 20116 13920
rect 20162 13880 20168 13932
rect 20220 13880 20226 13932
rect 20548 13929 20576 13960
rect 20640 13929 20668 14016
rect 22296 13997 22324 14028
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 23937 14059 23995 14065
rect 23937 14025 23949 14059
rect 23983 14056 23995 14059
rect 24946 14056 24952 14068
rect 23983 14028 24952 14056
rect 23983 14025 23995 14028
rect 23937 14019 23995 14025
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 22281 13991 22339 13997
rect 22051 13957 22109 13963
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 21358 13920 21364 13932
rect 20956 13892 21364 13920
rect 20956 13880 20962 13892
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 22051 13923 22063 13957
rect 22097 13923 22109 13957
rect 22281 13957 22293 13991
rect 22327 13957 22339 13991
rect 28442 13988 28448 14000
rect 22281 13951 22339 13957
rect 22379 13960 22876 13988
rect 22051 13920 22109 13923
rect 22379 13920 22407 13960
rect 21468 13892 22407 13920
rect 22557 13923 22615 13929
rect 7852 13824 8432 13852
rect 8956 13824 13584 13852
rect 7852 13784 7880 13824
rect 6104 13756 7880 13784
rect 7929 13787 7987 13793
rect 6104 13728 6132 13756
rect 7929 13753 7941 13787
rect 7975 13784 7987 13787
rect 7975 13756 8340 13784
rect 7975 13753 7987 13756
rect 7929 13747 7987 13753
rect 8312 13728 8340 13756
rect 4617 13719 4675 13725
rect 4617 13716 4629 13719
rect 4028 13688 4629 13716
rect 4028 13676 4034 13688
rect 4617 13685 4629 13688
rect 4663 13685 4675 13719
rect 4617 13679 4675 13685
rect 6086 13676 6092 13728
rect 6144 13676 6150 13728
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 8021 13719 8079 13725
rect 8021 13716 8033 13719
rect 7800 13688 8033 13716
rect 7800 13676 7806 13688
rect 8021 13685 8033 13688
rect 8067 13685 8079 13719
rect 8021 13679 8079 13685
rect 8294 13676 8300 13728
rect 8352 13676 8358 13728
rect 8404 13716 8432 13824
rect 9214 13744 9220 13796
rect 9272 13744 9278 13796
rect 9766 13784 9772 13796
rect 9324 13756 9772 13784
rect 9324 13716 9352 13756
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 13446 13744 13452 13796
rect 13504 13744 13510 13796
rect 8404 13688 9352 13716
rect 9398 13676 9404 13728
rect 9456 13676 9462 13728
rect 13556 13716 13584 13824
rect 14734 13812 14740 13864
rect 14792 13812 14798 13864
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 17092 13824 17141 13852
rect 17092 13812 17098 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 18046 13812 18052 13864
rect 18104 13852 18110 13864
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 18104 13824 18337 13852
rect 18104 13812 18110 13824
rect 18325 13821 18337 13824
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 20346 13852 20352 13864
rect 19576 13824 20352 13852
rect 19576 13812 19582 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 21468 13852 21496 13892
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 20496 13824 21496 13852
rect 20496 13812 20502 13824
rect 22002 13812 22008 13864
rect 22060 13852 22066 13864
rect 22572 13852 22600 13883
rect 22848 13864 22876 13960
rect 26988 13960 28448 13988
rect 26988 13932 27016 13960
rect 28442 13948 28448 13960
rect 28500 13988 28506 14000
rect 28500 13960 28580 13988
rect 28500 13948 28506 13960
rect 23750 13880 23756 13932
rect 23808 13880 23814 13932
rect 26970 13880 26976 13932
rect 27028 13880 27034 13932
rect 28258 13880 28264 13932
rect 28316 13929 28322 13932
rect 28552 13929 28580 13960
rect 28316 13883 28328 13929
rect 28537 13923 28595 13929
rect 28537 13889 28549 13923
rect 28583 13889 28595 13923
rect 28537 13883 28595 13889
rect 28316 13880 28322 13883
rect 22060 13824 22600 13852
rect 22060 13812 22066 13824
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 25590 13812 25596 13864
rect 25648 13852 25654 13864
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 25648 13824 25697 13852
rect 25648 13812 25654 13824
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 16942 13744 16948 13796
rect 17000 13744 17006 13796
rect 17218 13784 17224 13796
rect 17052 13756 17224 13784
rect 14458 13716 14464 13728
rect 13556 13688 14464 13716
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 16666 13676 16672 13728
rect 16724 13676 16730 13728
rect 17052 13725 17080 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 20073 13787 20131 13793
rect 17368 13756 18092 13784
rect 17368 13744 17374 13756
rect 17037 13719 17095 13725
rect 17037 13685 17049 13719
rect 17083 13685 17095 13719
rect 17037 13679 17095 13685
rect 17494 13676 17500 13728
rect 17552 13676 17558 13728
rect 17862 13676 17868 13728
rect 17920 13676 17926 13728
rect 17954 13676 17960 13728
rect 18012 13676 18018 13728
rect 18064 13716 18092 13756
rect 19306 13756 19932 13784
rect 19306 13728 19334 13756
rect 18966 13716 18972 13728
rect 18064 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19242 13676 19248 13728
rect 19300 13688 19334 13728
rect 19300 13676 19306 13688
rect 19794 13676 19800 13728
rect 19852 13676 19858 13728
rect 19904 13716 19932 13756
rect 20073 13753 20085 13787
rect 20119 13784 20131 13787
rect 21913 13787 21971 13793
rect 21913 13784 21925 13787
rect 20119 13756 21925 13784
rect 20119 13753 20131 13756
rect 20073 13747 20131 13753
rect 21913 13753 21925 13756
rect 21959 13753 21971 13787
rect 25961 13787 26019 13793
rect 25961 13784 25973 13787
rect 21913 13747 21971 13753
rect 22112 13756 25973 13784
rect 22112 13725 22140 13756
rect 25961 13753 25973 13756
rect 26007 13784 26019 13787
rect 27157 13787 27215 13793
rect 27157 13784 27169 13787
rect 26007 13756 27169 13784
rect 26007 13753 26019 13756
rect 25961 13747 26019 13753
rect 27157 13753 27169 13756
rect 27203 13753 27215 13787
rect 27157 13747 27215 13753
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 19904 13688 20269 13716
rect 20257 13685 20269 13688
rect 20303 13685 20315 13719
rect 20257 13679 20315 13685
rect 22097 13719 22155 13725
rect 22097 13685 22109 13719
rect 22143 13685 22155 13719
rect 22097 13679 22155 13685
rect 22370 13676 22376 13728
rect 22428 13676 22434 13728
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 2038 13512 2044 13524
rect 1452 13484 2044 13512
rect 1452 13472 1458 13484
rect 2038 13472 2044 13484
rect 2096 13512 2102 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 2096 13484 2145 13512
rect 2096 13472 2102 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 2133 13475 2191 13481
rect 2498 13472 2504 13524
rect 2556 13472 2562 13524
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 3384 13484 4721 13512
rect 3384 13472 3390 13484
rect 4709 13481 4721 13484
rect 4755 13512 4767 13515
rect 5442 13512 5448 13524
rect 4755 13484 5448 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 6270 13512 6276 13524
rect 6227 13484 6276 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9214 13512 9220 13524
rect 8803 13484 9220 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2516 13308 2544 13472
rect 4157 13447 4215 13453
rect 4157 13413 4169 13447
rect 4203 13444 4215 13447
rect 4203 13416 4476 13444
rect 4203 13413 4215 13416
rect 4157 13407 4215 13413
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 2363 13280 2605 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2593 13277 2605 13280
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13308 2835 13311
rect 2866 13308 2872 13320
rect 2823 13280 2872 13308
rect 2823 13277 2835 13280
rect 2777 13271 2835 13277
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 2792 13240 2820 13271
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13277 3939 13311
rect 3881 13271 3939 13277
rect 2547 13212 2820 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 3602 13200 3608 13252
rect 3660 13240 3666 13252
rect 3896 13240 3924 13271
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4448 13317 4476 13416
rect 4798 13336 4804 13388
rect 4856 13336 4862 13388
rect 7098 13376 7104 13388
rect 6196 13348 7104 13376
rect 6196 13320 6224 13348
rect 7098 13336 7104 13348
rect 7156 13376 7162 13388
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 7156 13348 7389 13376
rect 7156 13336 7162 13348
rect 7377 13345 7389 13348
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 6178 13268 6184 13320
rect 6236 13268 6242 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 3660 13212 3924 13240
rect 4157 13243 4215 13249
rect 3660 13200 3666 13212
rect 4157 13209 4169 13243
rect 4203 13209 4215 13243
rect 5046 13243 5104 13249
rect 5046 13240 5058 13243
rect 4157 13203 4215 13209
rect 4540 13212 5058 13240
rect 2590 13132 2596 13184
rect 2648 13132 2654 13184
rect 4172 13172 4200 13203
rect 4430 13172 4436 13184
rect 4172 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 4540 13181 4568 13212
rect 5046 13209 5058 13212
rect 5092 13209 5104 13243
rect 5046 13203 5104 13209
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13141 4583 13175
rect 4525 13135 4583 13141
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 6840 13172 6868 13271
rect 8938 13268 8944 13320
rect 8996 13268 9002 13320
rect 9048 13317 9076 13484
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 13633 13515 13691 13521
rect 10980 13484 13288 13512
rect 9674 13444 9680 13456
rect 9324 13416 9680 13444
rect 9324 13317 9352 13416
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 9600 13348 9812 13376
rect 9490 13317 9496 13320
rect 9034 13311 9092 13317
rect 9034 13277 9046 13311
rect 9080 13277 9092 13311
rect 9034 13271 9092 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 9447 13311 9496 13317
rect 9447 13277 9459 13311
rect 9493 13277 9496 13311
rect 9447 13271 9496 13277
rect 9490 13268 9496 13271
rect 9548 13268 9554 13320
rect 7650 13249 7656 13252
rect 7644 13203 7656 13249
rect 7650 13200 7656 13203
rect 7708 13200 7714 13252
rect 9122 13200 9128 13252
rect 9180 13240 9186 13252
rect 9217 13243 9275 13249
rect 9217 13240 9229 13243
rect 9180 13212 9229 13240
rect 9180 13200 9186 13212
rect 9217 13209 9229 13212
rect 9263 13209 9275 13243
rect 9600 13240 9628 13348
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 9784 13308 9812 13348
rect 10980 13308 11008 13484
rect 11057 13447 11115 13453
rect 11057 13413 11069 13447
rect 11103 13413 11115 13447
rect 11057 13407 11115 13413
rect 11072 13376 11100 13407
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 11204 13416 12296 13444
rect 11204 13404 11210 13416
rect 12268 13388 12296 13416
rect 11072 13348 11468 13376
rect 11440 13320 11468 13348
rect 12250 13336 12256 13388
rect 12308 13336 12314 13388
rect 13260 13376 13288 13484
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 14182 13512 14188 13524
rect 13679 13484 14188 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 15010 13472 15016 13524
rect 15068 13472 15074 13524
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 15804 13484 16405 13512
rect 15804 13472 15810 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16393 13475 16451 13481
rect 16666 13472 16672 13524
rect 16724 13472 16730 13524
rect 17310 13472 17316 13524
rect 17368 13472 17374 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 19702 13512 19708 13524
rect 17644 13484 19708 13512
rect 17644 13472 17650 13484
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19852 13484 19901 13512
rect 19852 13472 19858 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 20036 13484 20085 13512
rect 20036 13472 20042 13484
rect 20073 13481 20085 13484
rect 20119 13481 20131 13515
rect 20073 13475 20131 13481
rect 20714 13472 20720 13524
rect 20772 13472 20778 13524
rect 20809 13515 20867 13521
rect 20809 13481 20821 13515
rect 20855 13512 20867 13515
rect 20990 13512 20996 13524
rect 20855 13484 20996 13512
rect 20855 13481 20867 13484
rect 20809 13475 20867 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 22002 13472 22008 13524
rect 22060 13472 22066 13524
rect 23750 13472 23756 13524
rect 23808 13512 23814 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23808 13484 24041 13512
rect 23808 13472 23814 13484
rect 24029 13481 24041 13484
rect 24075 13481 24087 13515
rect 24029 13475 24087 13481
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 28077 13515 28135 13521
rect 27028 13484 27292 13512
rect 27028 13472 27034 13484
rect 14458 13404 14464 13456
rect 14516 13444 14522 13456
rect 21913 13447 21971 13453
rect 14516 13416 21501 13444
rect 14516 13404 14522 13416
rect 17494 13376 17500 13388
rect 13260 13348 15884 13376
rect 9784 13280 11008 13308
rect 9677 13271 9735 13277
rect 9217 13203 9275 13209
rect 9508 13212 9628 13240
rect 9508 13172 9536 13212
rect 6840 13144 9536 13172
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 9692 13172 9720 13271
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11204 13280 11345 13308
rect 11204 13268 11210 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11422 13268 11428 13320
rect 11480 13268 11486 13320
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 11698 13268 11704 13320
rect 11756 13268 11762 13320
rect 12526 13317 12532 13320
rect 11839 13311 11897 13317
rect 11839 13308 11851 13311
rect 11813 13277 11851 13308
rect 11885 13308 11897 13311
rect 12509 13311 12532 13317
rect 11885 13280 12480 13308
rect 11885 13277 11897 13280
rect 11813 13271 11897 13277
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 9922 13243 9980 13249
rect 9922 13240 9934 13243
rect 9824 13212 9934 13240
rect 9824 13200 9830 13212
rect 9922 13209 9934 13212
rect 9968 13209 9980 13243
rect 11072 13240 11100 13268
rect 9922 13203 9980 13209
rect 10060 13212 11100 13240
rect 10060 13184 10088 13212
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 11624 13240 11652 13268
rect 11296 13212 11652 13240
rect 11296 13200 11302 13212
rect 10042 13172 10048 13184
rect 9692 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 11054 13172 11060 13184
rect 10468 13144 11060 13172
rect 10468 13132 10474 13144
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11330 13132 11336 13184
rect 11388 13172 11394 13184
rect 11813 13172 11841 13271
rect 12452 13240 12480 13280
rect 12509 13277 12521 13311
rect 12509 13271 12532 13277
rect 12526 13268 12532 13271
rect 12584 13268 12590 13320
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 14424 13280 14565 13308
rect 14424 13268 14430 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 13280 13240 13308 13268
rect 12452 13212 13308 13240
rect 14737 13243 14795 13249
rect 14737 13209 14749 13243
rect 14783 13240 14795 13243
rect 14826 13240 14832 13252
rect 14783 13212 14832 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 14826 13200 14832 13212
rect 14884 13240 14890 13252
rect 15856 13240 15884 13348
rect 16592 13348 17500 13376
rect 16592 13317 16620 13348
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 17604 13348 19257 13376
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 17604 13308 17632 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 19978 13336 19984 13388
rect 20036 13376 20042 13388
rect 20036 13348 20944 13376
rect 20036 13336 20042 13348
rect 16776 13280 17632 13308
rect 16776 13240 16804 13280
rect 17678 13268 17684 13320
rect 17736 13268 17742 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18138 13308 18144 13320
rect 18012 13280 18144 13308
rect 18012 13268 18018 13280
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 14884 13212 15792 13240
rect 15856 13212 16804 13240
rect 16853 13243 16911 13249
rect 14884 13200 14890 13212
rect 11388 13144 11841 13172
rect 11977 13175 12035 13181
rect 11388 13132 11394 13144
rect 11977 13141 11989 13175
rect 12023 13172 12035 13175
rect 12342 13172 12348 13184
rect 12023 13144 12348 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14700 13144 14933 13172
rect 14700 13132 14706 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 15764 13172 15792 13212
rect 16853 13209 16865 13243
rect 16899 13240 16911 13243
rect 16899 13212 17448 13240
rect 16899 13209 16911 13212
rect 16853 13203 16911 13209
rect 17420 13184 17448 13212
rect 17494 13200 17500 13252
rect 17552 13200 17558 13252
rect 17696 13240 17724 13268
rect 18800 13240 18828 13271
rect 18966 13268 18972 13320
rect 19024 13268 19030 13320
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19576 13280 19625 13308
rect 19576 13268 19582 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 20349 13311 20407 13317
rect 20349 13308 20361 13311
rect 19797 13271 19855 13277
rect 20012 13280 20361 13308
rect 19150 13240 19156 13252
rect 17696 13212 19156 13240
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 19426 13200 19432 13252
rect 19484 13200 19490 13252
rect 19702 13200 19708 13252
rect 19760 13200 19766 13252
rect 19812 13240 19840 13271
rect 20012 13240 20040 13280
rect 20349 13277 20361 13280
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 20916 13317 20944 13348
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21473 13308 21501 13416
rect 21913 13413 21925 13447
rect 21959 13444 21971 13447
rect 22094 13444 22100 13456
rect 21959 13416 22100 13444
rect 21959 13413 21971 13416
rect 21913 13407 21971 13413
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 23934 13404 23940 13456
rect 23992 13404 23998 13456
rect 27264 13385 27292 13484
rect 28077 13481 28089 13515
rect 28123 13512 28135 13515
rect 28258 13512 28264 13524
rect 28123 13484 28264 13512
rect 28123 13481 28135 13484
rect 28077 13475 28135 13481
rect 28258 13472 28264 13484
rect 28316 13472 28322 13524
rect 27614 13404 27620 13456
rect 27672 13404 27678 13456
rect 27249 13379 27307 13385
rect 27249 13345 27261 13379
rect 27295 13345 27307 13379
rect 27249 13339 27307 13345
rect 27338 13336 27344 13388
rect 27396 13336 27402 13388
rect 27801 13379 27859 13385
rect 27801 13345 27813 13379
rect 27847 13376 27859 13379
rect 27847 13348 27936 13376
rect 27847 13345 27859 13348
rect 27801 13339 27859 13345
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21473 13280 21557 13308
rect 21085 13271 21143 13277
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13308 22155 13311
rect 22143 13280 24900 13308
rect 22143 13277 22155 13280
rect 22097 13271 22155 13277
rect 19812 13212 20040 13240
rect 20070 13200 20076 13252
rect 20128 13200 20134 13252
rect 21100 13240 21128 13271
rect 21358 13240 21364 13252
rect 21100 13212 21364 13240
rect 16574 13172 16580 13184
rect 15764 13144 16580 13172
rect 14921 13135 14979 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 17126 13132 17132 13184
rect 17184 13132 17190 13184
rect 17310 13181 17316 13184
rect 17297 13175 17316 13181
rect 17297 13141 17309 13175
rect 17297 13135 17316 13141
rect 17310 13132 17316 13135
rect 17368 13132 17374 13184
rect 17402 13132 17408 13184
rect 17460 13132 17466 13184
rect 17678 13132 17684 13184
rect 17736 13172 17742 13184
rect 18601 13175 18659 13181
rect 18601 13172 18613 13175
rect 17736 13144 18613 13172
rect 17736 13132 17742 13144
rect 18601 13141 18613 13144
rect 18647 13172 18659 13175
rect 21100 13172 21128 13212
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 18647 13144 21128 13172
rect 21560 13172 21588 13271
rect 22370 13249 22376 13252
rect 22364 13240 22376 13249
rect 22331 13212 22376 13240
rect 22364 13203 22376 13212
rect 22370 13200 22376 13203
rect 22428 13200 22434 13252
rect 23569 13243 23627 13249
rect 23569 13240 23581 13243
rect 23032 13212 23581 13240
rect 23032 13184 23060 13212
rect 23569 13209 23581 13212
rect 23615 13209 23627 13243
rect 23569 13203 23627 13209
rect 24872 13240 24900 13280
rect 24946 13268 24952 13320
rect 25004 13308 25010 13320
rect 27908 13317 27936 13348
rect 25510 13311 25568 13317
rect 25510 13308 25522 13311
rect 25004 13280 25522 13308
rect 25004 13268 25010 13280
rect 25510 13277 25522 13280
rect 25556 13277 25568 13311
rect 25510 13271 25568 13277
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 27893 13311 27951 13317
rect 27893 13277 27905 13311
rect 27939 13277 27951 13311
rect 27893 13271 27951 13277
rect 25792 13240 25820 13271
rect 25958 13240 25964 13252
rect 24872 13212 25964 13240
rect 23014 13172 23020 13184
rect 21560 13144 23020 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 23382 13132 23388 13184
rect 23440 13172 23446 13184
rect 23477 13175 23535 13181
rect 23477 13172 23489 13175
rect 23440 13144 23489 13172
rect 23440 13132 23446 13144
rect 23477 13141 23489 13144
rect 23523 13141 23535 13175
rect 23477 13135 23535 13141
rect 24394 13132 24400 13184
rect 24452 13132 24458 13184
rect 24872 13172 24900 13212
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 26234 13200 26240 13252
rect 26292 13240 26298 13252
rect 26982 13243 27040 13249
rect 26982 13240 26994 13243
rect 26292 13212 26994 13240
rect 26292 13200 26298 13212
rect 26982 13209 26994 13212
rect 27028 13209 27040 13243
rect 26982 13203 27040 13209
rect 24946 13172 24952 13184
rect 24872 13144 24952 13172
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 25130 13132 25136 13184
rect 25188 13172 25194 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 25188 13144 25881 13172
rect 25188 13132 25194 13144
rect 25869 13141 25881 13144
rect 25915 13141 25927 13175
rect 25869 13135 25927 13141
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 2866 12968 2872 12980
rect 2823 12940 2872 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 3099 12940 3740 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 2130 12900 2136 12912
rect 1412 12872 2136 12900
rect 1412 12841 1440 12872
rect 2130 12860 2136 12872
rect 2188 12900 2194 12912
rect 3712 12900 3740 12940
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 5166 12968 5172 12980
rect 4488 12940 5172 12968
rect 4488 12928 4494 12940
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 7650 12928 7656 12980
rect 7708 12928 7714 12980
rect 7742 12928 7748 12980
rect 7800 12928 7806 12980
rect 9306 12968 9312 12980
rect 9232 12940 9312 12968
rect 6638 12909 6644 12912
rect 3850 12903 3908 12909
rect 3850 12900 3862 12903
rect 2188 12872 2774 12900
rect 2188 12860 2194 12872
rect 1670 12841 1676 12844
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 1664 12795 1676 12841
rect 1670 12792 1676 12795
rect 1728 12792 1734 12844
rect 2746 12764 2774 12872
rect 3436 12872 3648 12900
rect 3712 12872 3862 12900
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3326 12832 3332 12844
rect 3283 12804 3332 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3436 12841 3464 12872
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 3620 12832 3648 12872
rect 3850 12869 3862 12872
rect 3896 12869 3908 12903
rect 6621 12903 6644 12909
rect 3850 12863 3908 12869
rect 5828 12872 6316 12900
rect 4154 12832 4160 12844
rect 3620 12804 4160 12832
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 5828 12841 5856 12872
rect 6288 12844 6316 12872
rect 6621 12869 6633 12903
rect 6621 12863 6644 12869
rect 6638 12860 6644 12863
rect 6696 12860 6702 12912
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 2746 12736 3617 12764
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 6012 12764 6040 12795
rect 6270 12792 6276 12844
rect 6328 12792 6334 12844
rect 6086 12764 6092 12776
rect 6012 12736 6092 12764
rect 3605 12727 3663 12733
rect 3620 12628 3648 12727
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 4982 12656 4988 12708
rect 5040 12656 5046 12708
rect 7668 12696 7696 12928
rect 7760 12832 7788 12928
rect 9232 12909 9260 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 10962 12928 10968 12980
rect 11020 12928 11026 12980
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12345 12971 12403 12977
rect 12345 12968 12357 12971
rect 12084 12940 12357 12968
rect 9217 12903 9275 12909
rect 9217 12869 9229 12903
rect 9263 12869 9275 12903
rect 9217 12863 9275 12869
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7760 12804 8033 12832
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 7837 12699 7895 12705
rect 7837 12696 7849 12699
rect 7668 12668 7849 12696
rect 7837 12665 7849 12668
rect 7883 12665 7895 12699
rect 7837 12659 7895 12665
rect 4338 12628 4344 12640
rect 3620 12600 4344 12628
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 6178 12588 6184 12640
rect 6236 12588 6242 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8294 12628 8300 12640
rect 7791 12600 8300 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8294 12588 8300 12600
rect 8352 12628 8358 12640
rect 8956 12628 8984 12795
rect 9122 12792 9128 12844
rect 9180 12792 9186 12844
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12801 9367 12835
rect 9416 12832 9444 12928
rect 10980 12900 11008 12928
rect 12084 12900 12112 12940
rect 12345 12937 12357 12940
rect 12391 12937 12403 12971
rect 12345 12931 12403 12937
rect 14642 12928 14648 12980
rect 14700 12928 14706 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 10980 12872 12112 12900
rect 12250 12860 12256 12912
rect 12308 12900 12314 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 12308 12872 12449 12900
rect 12308 12860 12314 12872
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 12912 12872 13860 12900
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9416 12804 9597 12832
rect 9309 12795 9367 12801
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 9140 12696 9168 12792
rect 9324 12764 9352 12795
rect 11422 12792 11428 12844
rect 11480 12792 11486 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11790 12832 11796 12844
rect 11563 12804 11796 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12802 12832 12808 12844
rect 12207 12804 12808 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 9490 12764 9496 12776
rect 9324 12736 9496 12764
rect 9490 12724 9496 12736
rect 9548 12764 9554 12776
rect 11330 12764 11336 12776
rect 9548 12736 11336 12764
rect 9548 12724 9554 12736
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 11238 12696 11244 12708
rect 9140 12668 11244 12696
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 11440 12696 11468 12792
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12912 12764 12940 12872
rect 13832 12844 13860 12872
rect 12986 12792 12992 12844
rect 13044 12792 13050 12844
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13245 12835 13303 12841
rect 13245 12832 13257 12835
rect 13136 12804 13257 12832
rect 13136 12792 13142 12804
rect 13245 12801 13257 12804
rect 13291 12801 13303 12835
rect 13245 12795 13303 12801
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14660 12832 14688 12928
rect 15028 12900 15056 12931
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 19245 12971 19303 12977
rect 17368 12940 18276 12968
rect 17368 12928 17374 12940
rect 15350 12903 15408 12909
rect 15350 12900 15362 12903
rect 15028 12872 15362 12900
rect 15350 12869 15362 12872
rect 15396 12869 15408 12903
rect 17678 12900 17684 12912
rect 15350 12863 15408 12869
rect 15948 12872 17684 12900
rect 15948 12844 15976 12872
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14660 12804 14841 12832
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 12115 12736 12940 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 11440 12668 11805 12696
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 12084 12696 12112 12727
rect 11793 12659 11851 12665
rect 11900 12668 12112 12696
rect 8352 12600 8984 12628
rect 8352 12588 8358 12600
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9272 12600 9505 12628
rect 9272 12588 9278 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 10870 12588 10876 12640
rect 10928 12628 10934 12640
rect 11900 12628 11928 12668
rect 12434 12656 12440 12708
rect 12492 12656 12498 12708
rect 14734 12696 14740 12708
rect 14301 12668 14740 12696
rect 10928 12600 11928 12628
rect 10928 12588 10934 12600
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 12216 12600 12265 12628
rect 12216 12588 12222 12600
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12452 12628 12480 12656
rect 14301 12628 14329 12668
rect 14734 12656 14740 12668
rect 14792 12696 14798 12708
rect 15120 12696 15148 12795
rect 15930 12792 15936 12844
rect 15988 12792 15994 12844
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16540 12804 17049 12832
rect 16540 12792 16546 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17420 12841 17448 12872
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 18110 12903 18168 12909
rect 18110 12900 18122 12903
rect 17788 12872 18122 12900
rect 17267 12835 17325 12841
rect 17267 12801 17279 12835
rect 17313 12832 17325 12835
rect 17405 12835 17463 12841
rect 17313 12801 17330 12832
rect 17267 12795 17330 12801
rect 17405 12801 17417 12835
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17302 12764 17330 12795
rect 17586 12792 17592 12844
rect 17644 12792 17650 12844
rect 16500 12736 17330 12764
rect 16500 12708 16528 12736
rect 14792 12668 15148 12696
rect 14792 12656 14798 12668
rect 16482 12656 16488 12708
rect 16540 12656 16546 12708
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 16632 12668 17080 12696
rect 16632 12656 16638 12668
rect 12452 12600 14329 12628
rect 12253 12591 12311 12597
rect 14366 12588 14372 12640
rect 14424 12588 14430 12640
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 16942 12588 16948 12640
rect 17000 12588 17006 12640
rect 17052 12628 17080 12668
rect 17126 12656 17132 12708
rect 17184 12696 17190 12708
rect 17310 12696 17316 12708
rect 17184 12668 17316 12696
rect 17184 12656 17190 12668
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17788 12705 17816 12872
rect 18110 12869 18122 12872
rect 18156 12869 18168 12903
rect 18248 12900 18276 12940
rect 19245 12937 19257 12971
rect 19291 12968 19303 12971
rect 19426 12968 19432 12980
rect 19291 12940 19432 12968
rect 19291 12937 19303 12940
rect 19245 12931 19303 12937
rect 19426 12928 19432 12940
rect 19484 12968 19490 12980
rect 19978 12968 19984 12980
rect 19484 12940 19984 12968
rect 19484 12928 19490 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 20257 12971 20315 12977
rect 20257 12968 20269 12971
rect 20128 12940 20269 12968
rect 20128 12928 20134 12940
rect 20257 12937 20269 12940
rect 20303 12937 20315 12971
rect 20257 12931 20315 12937
rect 20901 12971 20959 12977
rect 20901 12937 20913 12971
rect 20947 12968 20959 12971
rect 21358 12968 21364 12980
rect 20947 12940 21364 12968
rect 20947 12937 20959 12940
rect 20901 12931 20959 12937
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 25590 12968 25596 12980
rect 25096 12940 25596 12968
rect 25096 12928 25102 12940
rect 25590 12928 25596 12940
rect 25648 12968 25654 12980
rect 25648 12940 25728 12968
rect 25648 12928 25654 12940
rect 20438 12900 20444 12912
rect 18248 12872 20444 12900
rect 18110 12863 18168 12869
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 22097 12903 22155 12909
rect 21692 12872 22048 12900
rect 21692 12860 21698 12872
rect 22020 12844 22048 12872
rect 22097 12869 22109 12903
rect 22143 12900 22155 12903
rect 22143 12872 22968 12900
rect 22143 12869 22155 12872
rect 22097 12863 22155 12869
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 17954 12832 17960 12844
rect 17911 12804 17960 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 19150 12792 19156 12844
rect 19208 12832 19214 12844
rect 19208 12804 20852 12832
rect 19208 12792 19214 12804
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20128 12736 20729 12764
rect 20128 12724 20134 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20824 12764 20852 12804
rect 20990 12792 20996 12844
rect 21048 12792 21054 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 21100 12764 21128 12795
rect 21174 12792 21180 12844
rect 21232 12792 21238 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 20824 12736 21128 12764
rect 20717 12727 20775 12733
rect 17773 12699 17831 12705
rect 17773 12665 17785 12699
rect 17819 12665 17831 12699
rect 17773 12659 17831 12665
rect 20530 12656 20536 12708
rect 20588 12656 20594 12708
rect 20625 12699 20683 12705
rect 20625 12665 20637 12699
rect 20671 12696 20683 12699
rect 21192 12696 21220 12792
rect 22204 12764 22232 12795
rect 22278 12792 22284 12844
rect 22336 12841 22342 12844
rect 22336 12835 22365 12841
rect 22353 12832 22365 12835
rect 22940 12832 22968 12872
rect 23014 12860 23020 12912
rect 23072 12860 23078 12912
rect 25130 12900 25136 12912
rect 23768 12872 25136 12900
rect 23768 12832 23796 12872
rect 25130 12860 25136 12872
rect 25188 12860 25194 12912
rect 25700 12909 25728 12940
rect 26142 12928 26148 12980
rect 26200 12928 26206 12980
rect 26234 12928 26240 12980
rect 26292 12928 26298 12980
rect 27614 12928 27620 12980
rect 27672 12968 27678 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 27672 12940 28549 12968
rect 27672 12928 27678 12940
rect 28537 12937 28549 12940
rect 28583 12937 28595 12971
rect 28537 12931 28595 12937
rect 25685 12903 25743 12909
rect 25685 12869 25697 12903
rect 25731 12869 25743 12903
rect 25685 12863 25743 12869
rect 22353 12804 22876 12832
rect 22940 12804 23796 12832
rect 22353 12801 22365 12804
rect 22336 12795 22365 12801
rect 22336 12792 22342 12795
rect 20671 12668 21220 12696
rect 22112 12736 22232 12764
rect 22465 12767 22523 12773
rect 20671 12665 20683 12668
rect 20625 12659 20683 12665
rect 20714 12628 20720 12640
rect 17052 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21266 12588 21272 12640
rect 21324 12588 21330 12640
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 21821 12631 21879 12637
rect 21821 12628 21833 12631
rect 21692 12600 21833 12628
rect 21692 12588 21698 12600
rect 21821 12597 21833 12600
rect 21867 12597 21879 12631
rect 22112 12628 22140 12736
rect 22465 12733 22477 12767
rect 22511 12733 22523 12767
rect 22848 12764 22876 12804
rect 23842 12792 23848 12844
rect 23900 12832 23906 12844
rect 24774 12835 24832 12841
rect 24774 12832 24786 12835
rect 23900 12804 24786 12832
rect 23900 12792 23906 12804
rect 24774 12801 24786 12804
rect 24820 12801 24832 12835
rect 24774 12795 24832 12801
rect 24946 12792 24952 12844
rect 25004 12832 25010 12844
rect 25041 12835 25099 12841
rect 25041 12832 25053 12835
rect 25004 12804 25053 12832
rect 25004 12792 25010 12804
rect 25041 12801 25053 12804
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 23014 12764 23020 12776
rect 22848 12736 23020 12764
rect 22465 12727 22523 12733
rect 22186 12656 22192 12708
rect 22244 12696 22250 12708
rect 22480 12696 22508 12727
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 23934 12724 23940 12776
rect 23992 12724 23998 12776
rect 22244 12668 22508 12696
rect 22244 12656 22250 12668
rect 23382 12656 23388 12708
rect 23440 12656 23446 12708
rect 23566 12656 23572 12708
rect 23624 12696 23630 12708
rect 23661 12699 23719 12705
rect 23661 12696 23673 12699
rect 23624 12668 23673 12696
rect 23624 12656 23630 12668
rect 23661 12665 23673 12668
rect 23707 12696 23719 12699
rect 23952 12696 23980 12724
rect 23707 12668 23980 12696
rect 25148 12696 25176 12860
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26160 12832 26188 12928
rect 26099 12804 26188 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 26970 12792 26976 12844
rect 27028 12832 27034 12844
rect 27430 12841 27436 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 27028 12804 27169 12832
rect 27028 12792 27034 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27424 12795 27436 12841
rect 27430 12792 27436 12795
rect 27488 12792 27494 12844
rect 25317 12699 25375 12705
rect 25317 12696 25329 12699
rect 25148 12668 25329 12696
rect 23707 12665 23719 12668
rect 23661 12659 23719 12665
rect 25317 12665 25329 12668
rect 25363 12665 25375 12699
rect 25317 12659 25375 12665
rect 24394 12628 24400 12640
rect 22112 12600 24400 12628
rect 21821 12591 21879 12597
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 25222 12588 25228 12640
rect 25280 12588 25286 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1728 12396 1869 12424
rect 1728 12384 1734 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 1857 12387 1915 12393
rect 2056 12396 2789 12424
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 1762 12356 1768 12368
rect 1627 12328 1768 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 1762 12316 1768 12328
rect 1820 12316 1826 12368
rect 750 12180 756 12232
rect 808 12220 814 12232
rect 2056 12229 2084 12396
rect 2777 12393 2789 12396
rect 2823 12424 2835 12427
rect 3326 12424 3332 12436
rect 2823 12396 3332 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13078 12424 13084 12436
rect 13035 12396 13084 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 14424 12396 15485 12424
rect 14424 12384 14430 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 15838 12424 15844 12436
rect 15703 12396 15844 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 16117 12427 16175 12433
rect 16117 12393 16129 12427
rect 16163 12393 16175 12427
rect 16117 12387 16175 12393
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 17034 12424 17040 12436
rect 16347 12396 17040 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 7745 12359 7803 12365
rect 7745 12325 7757 12359
rect 7791 12356 7803 12359
rect 12529 12359 12587 12365
rect 12529 12356 12541 12359
rect 7791 12328 12541 12356
rect 7791 12325 7803 12328
rect 7745 12319 7803 12325
rect 12529 12325 12541 12328
rect 12575 12356 12587 12359
rect 16132 12356 16160 12387
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 17405 12427 17463 12433
rect 17405 12393 17417 12427
rect 17451 12424 17463 12427
rect 17586 12424 17592 12436
rect 17451 12396 17592 12424
rect 17451 12393 17463 12396
rect 17405 12387 17463 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18230 12384 18236 12436
rect 18288 12384 18294 12436
rect 18874 12384 18880 12436
rect 18932 12384 18938 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 19702 12424 19708 12436
rect 19659 12396 19708 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 21358 12424 21364 12436
rect 20824 12396 21364 12424
rect 12575 12328 16160 12356
rect 12575 12325 12587 12328
rect 12529 12319 12587 12325
rect 16482 12316 16488 12368
rect 16540 12316 16546 12368
rect 18141 12359 18199 12365
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 18892 12356 18920 12384
rect 20824 12368 20852 12396
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 23842 12384 23848 12436
rect 23900 12384 23906 12436
rect 27430 12384 27436 12436
rect 27488 12424 27494 12436
rect 27525 12427 27583 12433
rect 27525 12424 27537 12427
rect 27488 12396 27537 12424
rect 27488 12384 27494 12396
rect 27525 12393 27537 12396
rect 27571 12393 27583 12427
rect 27525 12387 27583 12393
rect 18187 12328 18920 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 19978 12316 19984 12368
rect 20036 12316 20042 12368
rect 20806 12316 20812 12368
rect 20864 12316 20870 12368
rect 20990 12316 20996 12368
rect 21048 12356 21054 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 21048 12328 21281 12356
rect 21048 12316 21054 12328
rect 21269 12325 21281 12328
rect 21315 12356 21327 12359
rect 22554 12356 22560 12368
rect 21315 12328 22560 12356
rect 21315 12325 21327 12328
rect 21269 12319 21327 12325
rect 22554 12316 22560 12328
rect 22612 12316 22618 12368
rect 6362 12248 6368 12300
rect 6420 12248 6426 12300
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 11974 12288 11980 12300
rect 7432 12260 11980 12288
rect 7432 12248 7438 12260
rect 11974 12248 11980 12260
rect 12032 12288 12038 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 12032 12260 12173 12288
rect 12032 12248 12038 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 12667 12260 12848 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 808 12192 1409 12220
rect 808 12180 814 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2222 12180 2228 12232
rect 2280 12180 2286 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2590 12220 2596 12232
rect 2363 12192 2596 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 3789 12223 3847 12229
rect 3789 12220 3801 12223
rect 3292 12192 3801 12220
rect 3292 12180 3298 12192
rect 3789 12189 3801 12192
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 12820 12229 12848 12260
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 15286 12288 15292 12300
rect 13872 12260 14872 12288
rect 13872 12248 13878 12260
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14844 12229 14872 12260
rect 15028 12260 15292 12288
rect 15028 12229 15056 12260
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15013 12223 15071 12229
rect 14875 12192 14964 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 2240 12152 2268 12180
rect 2501 12155 2559 12161
rect 2501 12152 2513 12155
rect 2240 12124 2513 12152
rect 2501 12121 2513 12124
rect 2547 12121 2559 12155
rect 6610 12155 6668 12161
rect 6610 12152 6622 12155
rect 2501 12115 2559 12121
rect 6288 12124 6622 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 6288 12093 6316 12124
rect 6610 12121 6622 12124
rect 6656 12121 6668 12155
rect 14642 12152 14648 12164
rect 6610 12115 6668 12121
rect 9646 12124 14648 12152
rect 9646 12096 9674 12124
rect 14642 12112 14648 12124
rect 14700 12152 14706 12164
rect 14936 12152 14964 12192
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12220 15255 12223
rect 15470 12220 15476 12232
rect 15243 12192 15476 12220
rect 15243 12189 15255 12192
rect 15197 12183 15255 12189
rect 15102 12152 15108 12164
rect 14700 12124 14872 12152
rect 14936 12124 15108 12152
rect 14700 12112 14706 12124
rect 2225 12087 2283 12093
rect 2225 12084 2237 12087
rect 2096 12056 2237 12084
rect 2096 12044 2102 12056
rect 2225 12053 2237 12056
rect 2271 12053 2283 12087
rect 2225 12047 2283 12053
rect 6273 12087 6331 12093
rect 6273 12053 6285 12087
rect 6319 12053 6331 12087
rect 6273 12047 6331 12053
rect 9582 12044 9588 12096
rect 9640 12056 9674 12096
rect 9640 12044 9646 12056
rect 14182 12044 14188 12096
rect 14240 12044 14246 12096
rect 14844 12084 14872 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15212 12152 15240 12183
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 16500 12220 16528 12316
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17460 12260 17785 12288
rect 17460 12248 17466 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 18340 12260 19196 12288
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 15948 12192 16268 12220
rect 16500 12192 17233 12220
rect 15948 12161 15976 12192
rect 15289 12155 15347 12161
rect 15289 12152 15301 12155
rect 15212 12124 15301 12152
rect 15289 12121 15301 12124
rect 15335 12121 15347 12155
rect 15289 12115 15347 12121
rect 15933 12155 15991 12161
rect 15933 12121 15945 12155
rect 15979 12121 15991 12155
rect 15933 12115 15991 12121
rect 15489 12087 15547 12093
rect 15489 12084 15501 12087
rect 14844 12056 15501 12084
rect 15489 12053 15501 12056
rect 15535 12084 15547 12087
rect 16022 12084 16028 12096
rect 15535 12056 16028 12084
rect 15535 12053 15547 12056
rect 15489 12047 15547 12053
rect 16022 12044 16028 12056
rect 16080 12084 16086 12096
rect 16133 12087 16191 12093
rect 16133 12084 16145 12087
rect 16080 12056 16145 12084
rect 16080 12044 16086 12056
rect 16133 12053 16145 12056
rect 16179 12053 16191 12087
rect 16240 12084 16268 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 17310 12180 17316 12232
rect 17368 12220 17374 12232
rect 17368 12192 18000 12220
rect 17368 12180 17374 12192
rect 17037 12155 17095 12161
rect 17037 12121 17049 12155
rect 17083 12152 17095 12155
rect 17770 12152 17776 12164
rect 17083 12124 17776 12152
rect 17083 12121 17095 12124
rect 17037 12115 17095 12121
rect 17770 12112 17776 12124
rect 17828 12112 17834 12164
rect 17972 12152 18000 12192
rect 18046 12180 18052 12232
rect 18104 12180 18110 12232
rect 18340 12229 18368 12260
rect 19168 12232 19196 12260
rect 19610 12248 19616 12300
rect 19668 12288 19674 12300
rect 20073 12291 20131 12297
rect 20073 12288 20085 12291
rect 19668 12260 20085 12288
rect 19668 12248 19674 12260
rect 20073 12257 20085 12260
rect 20119 12257 20131 12291
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20073 12251 20131 12257
rect 20164 12260 20913 12288
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 18524 12152 18552 12183
rect 18598 12180 18604 12232
rect 18656 12180 18662 12232
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 17972 12124 18552 12152
rect 18791 12152 18819 12183
rect 19150 12180 19156 12232
rect 19208 12180 19214 12232
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20164 12220 20192 12260
rect 20901 12257 20913 12260
rect 20947 12288 20959 12291
rect 21450 12288 21456 12300
rect 20947 12260 21456 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 20036 12192 20192 12220
rect 20349 12223 20407 12229
rect 20036 12180 20042 12192
rect 20349 12189 20361 12223
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 21085 12223 21143 12229
rect 21085 12189 21097 12223
rect 21131 12220 21143 12223
rect 21174 12220 21180 12232
rect 21131 12192 21180 12220
rect 21131 12189 21143 12192
rect 21085 12183 21143 12189
rect 19242 12152 19248 12164
rect 18791 12124 19248 12152
rect 17494 12084 17500 12096
rect 16240 12056 17500 12084
rect 16133 12047 16191 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 18524 12084 18552 12124
rect 19242 12112 19248 12124
rect 19300 12152 19306 12164
rect 20162 12152 20168 12164
rect 19300 12124 20168 12152
rect 19300 12112 19306 12124
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 20364 12152 20392 12183
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 23661 12223 23719 12229
rect 23661 12220 23673 12223
rect 23532 12192 23673 12220
rect 23532 12180 23538 12192
rect 23661 12189 23673 12192
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 25038 12180 25044 12232
rect 25096 12180 25102 12232
rect 26694 12180 26700 12232
rect 26752 12180 26758 12232
rect 27338 12180 27344 12232
rect 27396 12180 27402 12232
rect 26430 12155 26488 12161
rect 26430 12152 26442 12155
rect 20364 12124 20944 12152
rect 20916 12096 20944 12124
rect 25240 12124 26442 12152
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18524 12056 18981 12084
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 18969 12047 19027 12053
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12084 20315 12087
rect 20438 12084 20444 12096
rect 20303 12056 20444 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20898 12044 20904 12096
rect 20956 12084 20962 12096
rect 22186 12084 22192 12096
rect 20956 12056 22192 12084
rect 20956 12044 20962 12056
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 25240 12093 25268 12124
rect 26430 12121 26442 12124
rect 26476 12121 26488 12155
rect 26430 12115 26488 12121
rect 25225 12087 25283 12093
rect 25225 12053 25237 12087
rect 25271 12053 25283 12087
rect 25225 12047 25283 12053
rect 25317 12087 25375 12093
rect 25317 12053 25329 12087
rect 25363 12084 25375 12087
rect 25406 12084 25412 12096
rect 25363 12056 25412 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 25406 12044 25412 12056
rect 25464 12044 25470 12096
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3568 11852 3801 11880
rect 3568 11840 3574 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4212 11852 4353 11880
rect 4212 11840 4218 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4341 11843 4399 11849
rect 6086 11840 6092 11892
rect 6144 11880 6150 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6144 11852 6377 11880
rect 6144 11840 6150 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11849 9643 11883
rect 9585 11843 9643 11849
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 6825 11815 6883 11821
rect 3660 11784 4200 11812
rect 3660 11772 3666 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2958 11744 2964 11756
rect 2271 11716 2964 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4172 11753 4200 11784
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 7374 11812 7380 11824
rect 6871 11784 7380 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 9600 11812 9628 11843
rect 10042 11840 10048 11892
rect 10100 11840 10106 11892
rect 12158 11840 12164 11892
rect 12216 11840 12222 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 18598 11880 18604 11892
rect 14240 11852 18604 11880
rect 14240 11840 14246 11852
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19242 11840 19248 11892
rect 19300 11889 19306 11892
rect 19300 11883 19319 11889
rect 19307 11849 19319 11883
rect 19300 11843 19319 11849
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 19886 11880 19892 11892
rect 19475 11852 19892 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 19300 11840 19306 11843
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 21284 11852 21588 11880
rect 9922 11815 9980 11821
rect 9922 11812 9934 11815
rect 9600 11784 9934 11812
rect 9922 11781 9934 11784
rect 9968 11781 9980 11815
rect 9922 11775 9980 11781
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 4203 11716 4261 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4479 11716 4721 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 10060 11744 10088 11840
rect 11701 11815 11759 11821
rect 11701 11781 11713 11815
rect 11747 11812 11759 11815
rect 11790 11812 11796 11824
rect 11747 11784 11796 11812
rect 11747 11781 11759 11784
rect 11701 11775 11759 11781
rect 9723 11716 10088 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 2590 11676 2596 11688
rect 2363 11648 2596 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 3988 11676 4016 11704
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 3988 11648 5273 11676
rect 5261 11645 5273 11648
rect 5307 11645 5319 11679
rect 8036 11676 8064 11707
rect 8113 11679 8171 11685
rect 8113 11676 8125 11679
rect 8036 11648 8125 11676
rect 5261 11639 5319 11645
rect 8113 11645 8125 11648
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8619 11648 8769 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 8757 11645 8769 11648
rect 8803 11676 8815 11679
rect 9217 11679 9275 11685
rect 8803 11648 9168 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 2130 11568 2136 11620
rect 2188 11608 2194 11620
rect 2685 11611 2743 11617
rect 2685 11608 2697 11611
rect 2188 11580 2697 11608
rect 2188 11568 2194 11580
rect 2685 11577 2697 11580
rect 2731 11577 2743 11611
rect 2685 11571 2743 11577
rect 6549 11611 6607 11617
rect 6549 11577 6561 11611
rect 6595 11608 6607 11611
rect 8297 11611 8355 11617
rect 6595 11580 6868 11608
rect 6595 11577 6607 11580
rect 6549 11571 6607 11577
rect 6840 11552 6868 11580
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 8662 11608 8668 11620
rect 8343 11580 8668 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 9030 11568 9036 11620
rect 9088 11568 9094 11620
rect 1946 11500 1952 11552
rect 2004 11500 2010 11552
rect 2498 11500 2504 11552
rect 2556 11500 2562 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5776 11512 5825 11540
rect 5776 11500 5782 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 5813 11503 5871 11509
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7708 11512 7849 11540
rect 7708 11500 7714 11512
rect 7837 11509 7849 11512
rect 7883 11509 7895 11543
rect 9140 11540 9168 11648
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9416 11676 9444 11707
rect 11716 11676 11744 11775
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 15286 11772 15292 11824
rect 15344 11812 15350 11824
rect 16114 11812 16120 11824
rect 15344 11784 16120 11812
rect 15344 11772 15350 11784
rect 16114 11772 16120 11784
rect 16172 11772 16178 11824
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 21284 11821 21312 11852
rect 19061 11815 19119 11821
rect 19061 11812 19073 11815
rect 16356 11784 19073 11812
rect 16356 11772 16362 11784
rect 19061 11781 19073 11784
rect 19107 11781 19119 11815
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 19061 11775 19119 11781
rect 19306 11784 21281 11812
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12158 11744 12164 11756
rect 11940 11716 12164 11744
rect 11940 11704 11946 11716
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12802 11704 12808 11756
rect 12860 11704 12866 11756
rect 9263 11648 9444 11676
rect 10980 11648 11744 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 10980 11540 11008 11648
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 17126 11676 17132 11688
rect 14424 11648 17132 11676
rect 14424 11636 14430 11648
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 19076 11676 19104 11775
rect 19306 11756 19334 11784
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 21269 11775 21327 11781
rect 19242 11704 19248 11756
rect 19300 11716 19334 11756
rect 19300 11704 19306 11716
rect 20162 11704 20168 11756
rect 20220 11704 20226 11756
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20404 11716 21005 11744
rect 20404 11704 20410 11716
rect 20993 11713 21005 11716
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 21082 11704 21088 11756
rect 21140 11704 21146 11756
rect 21358 11704 21364 11756
rect 21416 11704 21422 11756
rect 21458 11747 21516 11753
rect 21458 11713 21470 11747
rect 21504 11713 21516 11747
rect 21458 11707 21516 11713
rect 19978 11676 19984 11688
rect 19076 11648 19984 11676
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 20898 11636 20904 11688
rect 20956 11636 20962 11688
rect 21473 11676 21501 11707
rect 21468 11648 21501 11676
rect 21560 11676 21588 11852
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 22462 11880 22468 11892
rect 21968 11852 22468 11880
rect 21968 11840 21974 11852
rect 22462 11840 22468 11852
rect 22520 11840 22526 11892
rect 22002 11772 22008 11824
rect 22060 11812 22066 11824
rect 22557 11815 22615 11821
rect 22557 11812 22569 11815
rect 22060 11784 22569 11812
rect 22060 11772 22066 11784
rect 22557 11781 22569 11784
rect 22603 11781 22615 11815
rect 22557 11775 22615 11781
rect 23014 11772 23020 11824
rect 23072 11821 23078 11824
rect 23072 11815 23101 11821
rect 23089 11781 23101 11815
rect 23072 11775 23101 11781
rect 24857 11815 24915 11821
rect 24857 11781 24869 11815
rect 24903 11812 24915 11815
rect 24946 11812 24952 11824
rect 24903 11784 24952 11812
rect 24903 11781 24915 11784
rect 24857 11775 24915 11781
rect 23072 11772 23078 11775
rect 24946 11772 24952 11784
rect 25004 11772 25010 11824
rect 21634 11704 21640 11756
rect 21692 11748 21698 11756
rect 21821 11748 21879 11753
rect 21692 11747 21879 11748
rect 21692 11720 21833 11747
rect 21692 11704 21698 11720
rect 21821 11713 21833 11720
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 21910 11704 21916 11756
rect 21968 11704 21974 11756
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22112 11676 22140 11707
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22286 11747 22344 11753
rect 22286 11713 22298 11747
rect 22332 11713 22344 11747
rect 22286 11707 22344 11713
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11713 22799 11747
rect 22741 11707 22799 11713
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 21560 11648 22140 11676
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 11698 11608 11704 11620
rect 11103 11580 11704 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 11698 11568 11704 11580
rect 11756 11608 11762 11620
rect 11977 11611 12035 11617
rect 11977 11608 11989 11611
rect 11756 11580 11989 11608
rect 11756 11568 11762 11580
rect 11977 11577 11989 11580
rect 12023 11577 12035 11611
rect 11977 11571 12035 11577
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 20916 11608 20944 11636
rect 21468 11608 21496 11648
rect 13872 11580 20484 11608
rect 20916 11580 21496 11608
rect 13872 11568 13878 11580
rect 9140 11512 11008 11540
rect 7837 11503 7895 11509
rect 12986 11500 12992 11552
rect 13044 11500 13050 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 19245 11543 19303 11549
rect 19245 11540 19257 11543
rect 18840 11512 19257 11540
rect 18840 11500 18846 11512
rect 19245 11509 19257 11512
rect 19291 11509 19303 11543
rect 19245 11503 19303 11509
rect 20346 11500 20352 11552
rect 20404 11500 20410 11552
rect 20456 11540 20484 11580
rect 21634 11568 21640 11620
rect 21692 11568 21698 11620
rect 22094 11568 22100 11620
rect 22152 11608 22158 11620
rect 22296 11608 22324 11707
rect 22756 11676 22784 11707
rect 22388 11648 22784 11676
rect 22388 11620 22416 11648
rect 22152 11580 22324 11608
rect 22152 11568 22158 11580
rect 22370 11568 22376 11620
rect 22428 11568 22434 11620
rect 22848 11608 22876 11707
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11744 23259 11747
rect 23382 11744 23388 11756
rect 23247 11716 23388 11744
rect 23247 11713 23259 11716
rect 23201 11707 23259 11713
rect 23382 11704 23388 11716
rect 23440 11704 23446 11756
rect 27430 11753 27436 11756
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 25332 11716 25421 11744
rect 25332 11685 25360 11716
rect 25409 11713 25421 11716
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 27424 11707 27436 11753
rect 27430 11704 27436 11707
rect 27488 11704 27494 11756
rect 25317 11679 25375 11685
rect 25317 11645 25329 11679
rect 25363 11645 25375 11679
rect 25317 11639 25375 11645
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 26694 11676 26700 11688
rect 26292 11648 26700 11676
rect 26292 11636 26298 11648
rect 26694 11636 26700 11648
rect 26752 11676 26758 11688
rect 27157 11679 27215 11685
rect 27157 11676 27169 11679
rect 26752 11648 27169 11676
rect 26752 11636 26758 11648
rect 27157 11645 27169 11648
rect 27203 11645 27215 11679
rect 27157 11639 27215 11645
rect 25133 11611 25191 11617
rect 25133 11608 25145 11611
rect 22848 11580 25145 11608
rect 25133 11577 25145 11580
rect 25179 11608 25191 11611
rect 25406 11608 25412 11620
rect 25179 11580 25412 11608
rect 25179 11577 25191 11580
rect 25133 11571 25191 11577
rect 25406 11568 25412 11580
rect 25464 11568 25470 11620
rect 21358 11540 21364 11552
rect 20456 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 22465 11543 22523 11549
rect 22465 11540 22477 11543
rect 21600 11512 22477 11540
rect 21600 11500 21606 11512
rect 22465 11509 22477 11512
rect 22511 11509 22523 11543
rect 22465 11503 22523 11509
rect 23658 11500 23664 11552
rect 23716 11540 23722 11552
rect 23934 11540 23940 11552
rect 23716 11512 23940 11540
rect 23716 11500 23722 11512
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 25590 11500 25596 11552
rect 25648 11500 25654 11552
rect 28537 11543 28595 11549
rect 28537 11509 28549 11543
rect 28583 11540 28595 11543
rect 28583 11512 28948 11540
rect 28583 11509 28595 11512
rect 28537 11503 28595 11509
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 5353 11339 5411 11345
rect 2556 11308 2774 11336
rect 2556 11296 2562 11308
rect 2746 11132 2774 11308
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5626 11336 5632 11348
rect 5399 11308 5632 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 9766 11336 9772 11348
rect 6880 11308 9772 11336
rect 6880 11296 6886 11308
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 10134 11336 10140 11348
rect 10091 11308 10140 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 10686 11296 10692 11348
rect 10744 11296 10750 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 14277 11339 14335 11345
rect 12584 11308 13676 11336
rect 12584 11296 12590 11308
rect 5166 11228 5172 11280
rect 5224 11228 5230 11280
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 9674 11268 9680 11280
rect 8803 11240 9076 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 9048 11212 9076 11240
rect 9232 11240 9680 11268
rect 9030 11160 9036 11212
rect 9088 11160 9094 11212
rect 5718 11141 5724 11144
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 2746 11104 3249 11132
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3651 11104 3801 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11101 5503 11135
rect 5712 11132 5724 11141
rect 5679 11104 5724 11132
rect 5445 11095 5503 11101
rect 5712 11095 5724 11104
rect 3142 11024 3148 11076
rect 3200 11024 3206 11076
rect 3421 11067 3479 11073
rect 3421 11033 3433 11067
rect 3467 11064 3479 11067
rect 4890 11064 4896 11076
rect 3467 11036 4896 11064
rect 3467 11033 3479 11036
rect 3421 11027 3479 11033
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5460 11064 5488 11095
rect 5718 11092 5724 11095
rect 5776 11092 5782 11144
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 7650 11141 7656 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7644 11132 7656 11141
rect 7611 11104 7656 11132
rect 7377 11095 7435 11101
rect 7644 11095 7656 11104
rect 6472 11064 6500 11092
rect 7392 11064 7420 11095
rect 7650 11092 7656 11095
rect 7708 11092 7714 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9232 11141 9260 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 10704 11268 10732 11296
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 10704 11240 10793 11268
rect 10781 11237 10793 11240
rect 10827 11268 10839 11271
rect 11330 11268 11336 11280
rect 10827 11240 11336 11268
rect 10827 11237 10839 11240
rect 10781 11231 10839 11237
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 13648 11212 13676 11308
rect 14277 11305 14289 11339
rect 14323 11305 14335 11339
rect 14277 11299 14335 11305
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13780 11240 14105 11268
rect 13780 11228 13786 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14292 11268 14320 11299
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 14516 11308 14749 11336
rect 14516 11296 14522 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 14737 11299 14795 11305
rect 15948 11308 27200 11336
rect 15948 11268 15976 11308
rect 14292 11240 15976 11268
rect 18509 11271 18567 11277
rect 14093 11231 14151 11237
rect 18509 11237 18521 11271
rect 18555 11237 18567 11271
rect 18509 11231 18567 11237
rect 9306 11160 9312 11212
rect 9364 11200 9370 11212
rect 9364 11172 9444 11200
rect 9364 11160 9370 11172
rect 9416 11141 9444 11172
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 10594 11160 10600 11212
rect 10652 11200 10658 11212
rect 10652 11172 11008 11200
rect 10652 11160 10658 11172
rect 9191 11135 9260 11141
rect 9191 11132 9203 11135
rect 8904 11104 9203 11132
rect 8904 11092 8910 11104
rect 9191 11101 9203 11104
rect 9237 11104 9260 11135
rect 9401 11135 9459 11141
rect 9237 11101 9249 11104
rect 9191 11095 9249 11101
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9582 11132 9588 11144
rect 9539 11104 9588 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10980 11141 11008 11172
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 14240 11172 14504 11200
rect 14240 11160 14246 11172
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 9723 11104 10057 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10045 11101 10057 11104
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13366 11135 13424 11141
rect 13366 11132 13378 11135
rect 13044 11104 13378 11132
rect 13044 11092 13050 11104
rect 13366 11101 13378 11104
rect 13412 11101 13424 11135
rect 13366 11095 13424 11101
rect 5460 11036 7420 11064
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 9769 11067 9827 11073
rect 9769 11033 9781 11067
rect 9815 11033 9827 11067
rect 13814 11064 13820 11076
rect 9769 11027 9827 11033
rect 10152 11036 13820 11064
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 7098 10956 7104 11008
rect 7156 10956 7162 11008
rect 9324 10996 9352 11027
rect 9674 10996 9680 11008
rect 9324 10968 9680 10996
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 9784 10996 9812 11027
rect 10152 10996 10180 11036
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14261 11067 14319 11073
rect 14261 11033 14273 11067
rect 14307 11064 14319 11067
rect 14366 11064 14372 11076
rect 14307 11036 14372 11064
rect 14307 11033 14319 11036
rect 14261 11027 14319 11033
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 14476 11073 14504 11172
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14700 11172 14764 11200
rect 14700 11160 14706 11172
rect 14736 11073 14764 11172
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18524 11200 18552 11231
rect 20346 11228 20352 11280
rect 20404 11228 20410 11280
rect 23569 11271 23627 11277
rect 23569 11268 23581 11271
rect 22066 11240 23581 11268
rect 20364 11200 20392 11228
rect 18012 11172 18460 11200
rect 18524 11172 19380 11200
rect 20364 11172 20852 11200
rect 18012 11160 18018 11172
rect 15930 11092 15936 11144
rect 15988 11092 15994 11144
rect 16758 11132 16764 11144
rect 16132 11104 16764 11132
rect 14461 11067 14519 11073
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 14721 11067 14779 11073
rect 14507 11036 14688 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 9784 10968 10180 10996
rect 10226 10956 10232 11008
rect 10284 10956 10290 11008
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 11974 10996 11980 11008
rect 10560 10968 11980 10996
rect 10560 10956 10566 10968
rect 11974 10956 11980 10968
rect 12032 10996 12038 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 12032 10968 12265 10996
rect 12032 10956 12038 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 12253 10959 12311 10965
rect 14550 10956 14556 11008
rect 14608 10956 14614 11008
rect 14660 10996 14688 11036
rect 14721 11033 14733 11067
rect 14767 11033 14779 11067
rect 14721 11027 14779 11033
rect 14921 11067 14979 11073
rect 14921 11033 14933 11067
rect 14967 11033 14979 11067
rect 14921 11027 14979 11033
rect 15473 11067 15531 11073
rect 15473 11033 15485 11067
rect 15519 11033 15531 11067
rect 15473 11027 15531 11033
rect 15657 11067 15715 11073
rect 15657 11033 15669 11067
rect 15703 11064 15715 11067
rect 16022 11064 16028 11076
rect 15703 11036 16028 11064
rect 15703 11033 15715 11036
rect 15657 11027 15715 11033
rect 14936 10996 14964 11027
rect 14660 10968 14964 10996
rect 15488 10996 15516 11027
rect 16022 11024 16028 11036
rect 16080 11064 16086 11076
rect 16132 11064 16160 11104
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17552 11104 17877 11132
rect 17552 11092 17558 11104
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 16206 11073 16212 11076
rect 16080 11036 16160 11064
rect 16080 11024 16086 11036
rect 16200 11027 16212 11073
rect 16206 11024 16212 11027
rect 16264 11024 16270 11076
rect 18064 11064 18092 11095
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 18432 11132 18460 11172
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18432 11104 19257 11132
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19352 11132 19380 11172
rect 19501 11135 19559 11141
rect 19501 11132 19513 11135
rect 19352 11104 19513 11132
rect 19245 11095 19303 11101
rect 19501 11101 19513 11104
rect 19547 11101 19559 11135
rect 19501 11095 19559 11101
rect 17696 11036 18092 11064
rect 19260 11064 19288 11095
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 20824 11132 20852 11172
rect 20973 11135 21031 11141
rect 20973 11132 20985 11135
rect 20824 11104 20985 11132
rect 20973 11101 20985 11104
rect 21019 11101 21031 11135
rect 20973 11095 21031 11101
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 22066 11132 22094 11240
rect 23569 11237 23581 11240
rect 23615 11237 23627 11271
rect 23569 11231 23627 11237
rect 23658 11228 23664 11280
rect 23716 11268 23722 11280
rect 27172 11277 27200 11308
rect 27338 11296 27344 11348
rect 27396 11296 27402 11348
rect 27430 11296 27436 11348
rect 27488 11296 27494 11348
rect 24765 11271 24823 11277
rect 24765 11268 24777 11271
rect 23716 11240 24777 11268
rect 23716 11228 23722 11240
rect 24765 11237 24777 11240
rect 24811 11237 24823 11271
rect 24765 11231 24823 11237
rect 27157 11271 27215 11277
rect 27157 11237 27169 11271
rect 27203 11268 27215 11271
rect 28920 11268 28948 11512
rect 27203 11240 28948 11268
rect 27203 11237 27215 11240
rect 27157 11231 27215 11237
rect 23109 11203 23167 11209
rect 23109 11169 23121 11203
rect 23155 11200 23167 11203
rect 23198 11200 23204 11212
rect 23155 11172 23204 11200
rect 23155 11169 23167 11172
rect 23109 11163 23167 11169
rect 23198 11160 23204 11172
rect 23256 11160 23262 11212
rect 23477 11203 23535 11209
rect 23477 11169 23489 11203
rect 23523 11200 23535 11203
rect 23842 11200 23848 11212
rect 23523 11172 23848 11200
rect 23523 11169 23535 11172
rect 23477 11163 23535 11169
rect 23842 11160 23848 11172
rect 23900 11200 23906 11212
rect 24854 11200 24860 11212
rect 23900 11172 23980 11200
rect 23900 11160 23906 11172
rect 21416 11104 22094 11132
rect 21416 11092 21422 11104
rect 22554 11092 22560 11144
rect 22612 11092 22618 11144
rect 23290 11092 23296 11144
rect 23348 11092 23354 11144
rect 23952 11141 23980 11172
rect 24136 11172 24860 11200
rect 24136 11141 24164 11172
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 23707 11135 23765 11141
rect 23707 11101 23719 11135
rect 23753 11101 23765 11135
rect 23707 11095 23765 11101
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24120 11135 24178 11141
rect 24120 11101 24132 11135
rect 24166 11101 24178 11135
rect 24120 11095 24178 11101
rect 20732 11064 20760 11092
rect 21910 11064 21916 11076
rect 19260 11036 20760 11064
rect 20916 11036 21916 11064
rect 17696 11008 17724 11036
rect 15746 10996 15752 11008
rect 15488 10968 15752 10996
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17313 10999 17371 11005
rect 17313 10996 17325 10999
rect 17000 10968 17325 10996
rect 17000 10956 17006 10968
rect 17313 10965 17325 10968
rect 17359 10965 17371 10999
rect 17313 10959 17371 10965
rect 17678 10956 17684 11008
rect 17736 10956 17742 11008
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 18233 10999 18291 11005
rect 18233 10996 18245 10999
rect 17828 10968 18245 10996
rect 17828 10956 17834 10968
rect 18233 10965 18245 10968
rect 18279 10996 18291 10999
rect 19242 10996 19248 11008
rect 18279 10968 19248 10996
rect 18279 10965 18291 10968
rect 18233 10959 18291 10965
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 20530 10956 20536 11008
rect 20588 10996 20594 11008
rect 20625 10999 20683 11005
rect 20625 10996 20637 10999
rect 20588 10968 20637 10996
rect 20588 10956 20594 10968
rect 20625 10965 20637 10968
rect 20671 10996 20683 10999
rect 20916 10996 20944 11036
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 22572 11064 22600 11092
rect 23474 11064 23480 11076
rect 22572 11036 23480 11064
rect 23474 11024 23480 11036
rect 23532 11064 23538 11076
rect 23722 11064 23750 11095
rect 24210 11092 24216 11144
rect 24268 11092 24274 11144
rect 25590 11092 25596 11144
rect 25648 11132 25654 11144
rect 25878 11135 25936 11141
rect 25878 11132 25890 11135
rect 25648 11104 25890 11132
rect 25648 11092 25654 11104
rect 25878 11101 25890 11104
rect 25924 11101 25936 11135
rect 25878 11095 25936 11101
rect 26145 11135 26203 11141
rect 26145 11101 26157 11135
rect 26191 11132 26203 11135
rect 26234 11132 26240 11144
rect 26191 11104 26240 11132
rect 26191 11101 26203 11104
rect 26145 11095 26203 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 27430 11092 27436 11144
rect 27488 11132 27494 11144
rect 27617 11135 27675 11141
rect 27617 11132 27629 11135
rect 27488 11104 27629 11132
rect 27488 11092 27494 11104
rect 27617 11101 27629 11104
rect 27663 11101 27675 11135
rect 27617 11095 27675 11101
rect 23532 11036 23750 11064
rect 23845 11067 23903 11073
rect 23532 11024 23538 11036
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24394 11064 24400 11076
rect 23891 11036 24400 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 26878 11024 26884 11076
rect 26936 11024 26942 11076
rect 20671 10968 20944 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 22097 10999 22155 11005
rect 22097 10996 22109 10999
rect 21140 10968 22109 10996
rect 21140 10956 21146 10968
rect 22097 10965 22109 10968
rect 22143 10965 22155 10999
rect 22097 10959 22155 10965
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1946 10752 1952 10804
rect 2004 10792 2010 10804
rect 2004 10764 2636 10792
rect 2004 10752 2010 10764
rect 1854 10684 1860 10736
rect 1912 10724 1918 10736
rect 1912 10696 2452 10724
rect 1912 10684 1918 10696
rect 750 10616 756 10668
rect 808 10656 814 10668
rect 2424 10665 2452 10696
rect 2608 10665 2636 10764
rect 2958 10752 2964 10804
rect 3016 10752 3022 10804
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10761 6055 10795
rect 9030 10792 9036 10804
rect 5997 10755 6055 10761
rect 6104 10764 9036 10792
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4074 10727 4132 10733
rect 4074 10724 4086 10727
rect 4028 10696 4086 10724
rect 4028 10684 4034 10696
rect 4074 10693 4086 10696
rect 4120 10693 4132 10727
rect 4074 10687 4132 10693
rect 5074 10684 5080 10736
rect 5132 10684 5138 10736
rect 5660 10727 5718 10733
rect 5660 10693 5672 10727
rect 5706 10724 5718 10727
rect 6012 10724 6040 10755
rect 5706 10696 6040 10724
rect 5706 10693 5718 10696
rect 5660 10687 5718 10693
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 808 10628 1501 10656
rect 808 10616 814 10628
rect 1489 10625 1501 10628
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 4338 10616 4344 10668
rect 4396 10616 4402 10668
rect 5092 10656 5120 10684
rect 6104 10656 6132 10764
rect 7000 10727 7058 10733
rect 7000 10693 7012 10727
rect 7046 10724 7058 10727
rect 7098 10724 7104 10736
rect 7046 10696 7104 10724
rect 7046 10693 7058 10696
rect 7000 10687 7058 10693
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 8846 10733 8852 10736
rect 8823 10727 8852 10733
rect 8823 10693 8835 10727
rect 8823 10687 8852 10693
rect 8846 10684 8852 10687
rect 8904 10684 8910 10736
rect 8956 10733 8984 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9582 10792 9588 10804
rect 9140 10764 9588 10792
rect 8941 10727 8999 10733
rect 8941 10693 8953 10727
rect 8987 10693 8999 10727
rect 8941 10687 8999 10693
rect 5092 10628 6132 10656
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6512 10628 6745 10656
rect 6512 10616 6518 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 8662 10616 8668 10668
rect 8720 10616 8726 10668
rect 9140 10665 9168 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 9950 10792 9956 10804
rect 9907 10764 9956 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10502 10752 10508 10804
rect 10560 10752 10566 10804
rect 10689 10795 10747 10801
rect 10689 10761 10701 10795
rect 10735 10792 10747 10795
rect 10778 10792 10784 10804
rect 10735 10764 10784 10792
rect 10735 10761 10747 10764
rect 10689 10755 10747 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11882 10752 11888 10804
rect 11940 10752 11946 10804
rect 12250 10752 12256 10804
rect 12308 10752 12314 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16022 10792 16028 10804
rect 15979 10764 16028 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 11149 10727 11207 10733
rect 11149 10724 11161 10727
rect 9548 10696 11161 10724
rect 9548 10684 9554 10696
rect 11149 10693 11161 10696
rect 11195 10693 11207 10727
rect 11149 10687 11207 10693
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11793 10727 11851 10733
rect 11793 10724 11805 10727
rect 11388 10696 11805 10724
rect 11388 10684 11394 10696
rect 11793 10693 11805 10696
rect 11839 10693 11851 10727
rect 11900 10724 11928 10752
rect 14476 10724 14504 10755
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16908 10764 17049 10792
rect 16908 10752 16914 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 17954 10792 17960 10804
rect 17727 10764 17960 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 18322 10752 18328 10804
rect 18380 10752 18386 10804
rect 18769 10795 18827 10801
rect 18769 10761 18781 10795
rect 18815 10792 18827 10795
rect 19978 10792 19984 10804
rect 18815 10764 19984 10792
rect 18815 10761 18827 10764
rect 18769 10755 18827 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 20220 10764 20361 10792
rect 20220 10752 20226 10764
rect 20349 10761 20361 10764
rect 20395 10761 20407 10795
rect 22097 10795 22155 10801
rect 20349 10755 20407 10761
rect 20456 10764 20944 10792
rect 14798 10727 14856 10733
rect 14798 10724 14810 10727
rect 11900 10696 12020 10724
rect 14476 10696 14810 10724
rect 11793 10687 11851 10693
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6472 10588 6500 10616
rect 5960 10560 6500 10588
rect 5960 10548 5966 10560
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 9048 10520 9076 10619
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 10870 10616 10876 10668
rect 10928 10616 10934 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11698 10665 11704 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11296 10628 11529 10656
rect 11296 10616 11302 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11665 10659 11704 10665
rect 11665 10625 11677 10659
rect 11665 10619 11704 10625
rect 11698 10616 11704 10619
rect 11756 10616 11762 10668
rect 11992 10665 12020 10696
rect 14798 10693 14810 10696
rect 14844 10693 14856 10727
rect 14798 10687 14856 10693
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 15252 10696 16344 10724
rect 15252 10684 15258 10696
rect 16316 10668 16344 10696
rect 16942 10684 16948 10736
rect 17000 10724 17006 10736
rect 18969 10727 19027 10733
rect 17000 10696 18000 10724
rect 17000 10684 17006 10696
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11982 10659 12040 10665
rect 11982 10625 11994 10659
rect 12028 10625 12040 10659
rect 11982 10619 12040 10625
rect 9306 10588 9312 10600
rect 7800 10492 9076 10520
rect 9232 10560 9312 10588
rect 7800 10480 7806 10492
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5166 10452 5172 10464
rect 4571 10424 5172 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 5684 10424 8125 10452
rect 5684 10412 5690 10424
rect 8113 10421 8125 10424
rect 8159 10452 8171 10455
rect 9232 10452 9260 10560
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10888 10588 10916 10616
rect 10183 10560 10916 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 11054 10548 11060 10600
rect 11112 10548 11118 10600
rect 11900 10532 11928 10619
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12400 10628 12449 10656
rect 12400 10616 12406 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 12986 10656 12992 10668
rect 12759 10628 12992 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13170 10656 13176 10668
rect 13127 10628 13176 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13538 10656 13544 10668
rect 13403 10628 13544 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 13280 10588 13308 10619
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 14274 10616 14280 10668
rect 14332 10616 14338 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15896 10628 16037 10656
rect 15896 10616 15902 10628
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 16356 10628 17509 10656
rect 16356 10616 16362 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17710 10659 17768 10665
rect 17710 10656 17722 10659
rect 17644 10628 17722 10656
rect 17644 10616 17650 10628
rect 17710 10625 17722 10628
rect 17756 10625 17768 10659
rect 17710 10619 17768 10625
rect 13648 10588 13676 10616
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13280 10560 13584 10588
rect 13648 10560 14565 10588
rect 11882 10480 11888 10532
rect 11940 10480 11946 10532
rect 12161 10523 12219 10529
rect 12161 10489 12173 10523
rect 12207 10520 12219 10523
rect 12207 10492 12480 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 8159 10424 9260 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 10870 10412 10876 10464
rect 10928 10412 10934 10464
rect 12452 10461 12480 10492
rect 13556 10461 13584 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17184 10560 17877 10588
rect 17184 10548 17190 10560
rect 17865 10557 17877 10560
rect 17911 10557 17923 10591
rect 17865 10551 17923 10557
rect 15746 10480 15752 10532
rect 15804 10480 15810 10532
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 17972 10520 18000 10696
rect 18969 10693 18981 10727
rect 19015 10724 19027 10727
rect 19058 10724 19064 10736
rect 19015 10696 19064 10724
rect 19015 10693 19027 10696
rect 18969 10687 19027 10693
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 19610 10684 19616 10736
rect 19668 10724 19674 10736
rect 20456 10724 20484 10764
rect 19668 10696 20484 10724
rect 19668 10684 19674 10696
rect 20530 10684 20536 10736
rect 20588 10684 20594 10736
rect 20916 10733 20944 10764
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 22646 10792 22652 10804
rect 22143 10764 22652 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 22741 10795 22799 10801
rect 22741 10761 22753 10795
rect 22787 10792 22799 10795
rect 23382 10792 23388 10804
rect 22787 10764 23388 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23842 10752 23848 10804
rect 23900 10752 23906 10804
rect 27430 10752 27436 10804
rect 27488 10752 27494 10804
rect 20901 10727 20959 10733
rect 20901 10693 20913 10727
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 21082 10684 21088 10736
rect 21140 10684 21146 10736
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 23106 10724 23112 10736
rect 21324 10696 23112 10724
rect 21324 10684 21330 10696
rect 23106 10684 23112 10696
rect 23164 10684 23170 10736
rect 23661 10727 23719 10733
rect 23661 10693 23673 10727
rect 23707 10724 23719 10727
rect 23860 10724 23888 10752
rect 23707 10696 23888 10724
rect 24397 10727 24455 10733
rect 23707 10693 23719 10696
rect 23661 10687 23719 10693
rect 24397 10693 24409 10727
rect 24443 10724 24455 10727
rect 24670 10724 24676 10736
rect 24443 10696 24676 10724
rect 24443 10693 24455 10696
rect 24397 10687 24455 10693
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 24946 10684 24952 10736
rect 25004 10724 25010 10736
rect 25317 10727 25375 10733
rect 25317 10724 25329 10727
rect 25004 10696 25329 10724
rect 25004 10684 25010 10696
rect 25317 10693 25329 10696
rect 25363 10724 25375 10727
rect 26878 10724 26884 10736
rect 25363 10696 26884 10724
rect 25363 10693 25375 10696
rect 25317 10687 25375 10693
rect 26878 10684 26884 10696
rect 26936 10724 26942 10736
rect 26973 10727 27031 10733
rect 26973 10724 26985 10727
rect 26936 10696 26985 10724
rect 26936 10684 26942 10696
rect 26973 10693 26985 10696
rect 27019 10693 27031 10727
rect 26973 10687 27031 10693
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 19981 10659 20039 10665
rect 19981 10656 19993 10659
rect 18288 10628 19993 10656
rect 18288 10616 18294 10628
rect 19981 10625 19993 10628
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 20548 10656 20576 10684
rect 20211 10628 20576 10656
rect 22833 10659 22891 10665
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 22833 10625 22845 10659
rect 22879 10656 22891 10659
rect 23014 10656 23020 10668
rect 22879 10628 23020 10656
rect 22879 10625 22891 10628
rect 22833 10619 22891 10625
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23474 10665 23480 10668
rect 23472 10656 23480 10665
rect 23435 10628 23480 10656
rect 23472 10619 23480 10628
rect 23474 10616 23480 10619
rect 23532 10616 23538 10668
rect 23566 10616 23572 10668
rect 23624 10616 23630 10668
rect 23750 10616 23756 10668
rect 23808 10665 23814 10668
rect 23808 10659 23847 10665
rect 23835 10625 23847 10659
rect 23808 10619 23847 10625
rect 23937 10660 23995 10665
rect 24029 10660 24087 10665
rect 23937 10659 24087 10660
rect 23937 10625 23949 10659
rect 23983 10632 24041 10659
rect 23983 10625 23995 10632
rect 23937 10619 23995 10625
rect 24029 10625 24041 10632
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 23808 10616 23814 10619
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 18380 10560 23336 10588
rect 18380 10548 18386 10560
rect 18141 10523 18199 10529
rect 18141 10520 18153 10523
rect 17359 10492 17724 10520
rect 17972 10492 18153 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10421 12495 10455
rect 12437 10415 12495 10421
rect 13541 10455 13599 10461
rect 13541 10421 13553 10455
rect 13587 10452 13599 10455
rect 15764 10452 15792 10480
rect 13587 10424 15792 10452
rect 13587 10421 13599 10424
rect 13541 10415 13599 10421
rect 17402 10412 17408 10464
rect 17460 10412 17466 10464
rect 17696 10452 17724 10492
rect 18141 10489 18153 10492
rect 18187 10489 18199 10523
rect 23014 10520 23020 10532
rect 18141 10483 18199 10489
rect 18800 10492 23020 10520
rect 18800 10461 18828 10492
rect 23014 10480 23020 10492
rect 23072 10480 23078 10532
rect 23308 10529 23336 10560
rect 23382 10548 23388 10600
rect 23440 10588 23446 10600
rect 24228 10588 24256 10619
rect 24302 10616 24308 10668
rect 24360 10616 24366 10668
rect 24515 10659 24573 10665
rect 24515 10656 24527 10659
rect 24504 10625 24527 10656
rect 24561 10625 24573 10659
rect 24504 10619 24573 10625
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10625 26111 10659
rect 26053 10619 26111 10625
rect 23440 10560 24256 10588
rect 23440 10548 23446 10560
rect 24044 10532 24072 10560
rect 24504 10532 24532 10619
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 25777 10591 25835 10597
rect 25777 10557 25789 10591
rect 25823 10588 25835 10591
rect 26068 10588 26096 10619
rect 25823 10560 26096 10588
rect 25823 10557 25835 10560
rect 25777 10551 25835 10557
rect 23293 10523 23351 10529
rect 23293 10489 23305 10523
rect 23339 10489 23351 10523
rect 23293 10483 23351 10489
rect 24026 10480 24032 10532
rect 24084 10480 24090 10532
rect 24486 10480 24492 10532
rect 24544 10480 24550 10532
rect 24688 10520 24716 10551
rect 25682 10520 25688 10532
rect 24688 10492 25688 10520
rect 25682 10480 25688 10492
rect 25740 10480 25746 10532
rect 27249 10523 27307 10529
rect 27249 10520 27261 10523
rect 25792 10492 27261 10520
rect 18601 10455 18659 10461
rect 18601 10452 18613 10455
rect 17696 10424 18613 10452
rect 18601 10421 18613 10424
rect 18647 10421 18659 10455
rect 18601 10415 18659 10421
rect 18785 10455 18843 10461
rect 18785 10421 18797 10455
rect 18831 10421 18843 10455
rect 18785 10415 18843 10421
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 22373 10455 22431 10461
rect 22373 10452 22385 10455
rect 22244 10424 22385 10452
rect 22244 10412 22250 10424
rect 22373 10421 22385 10424
rect 22419 10421 22431 10455
rect 22373 10415 22431 10421
rect 22462 10412 22468 10464
rect 22520 10412 22526 10464
rect 22554 10412 22560 10464
rect 22612 10412 22618 10464
rect 23934 10412 23940 10464
rect 23992 10452 23998 10464
rect 25792 10452 25820 10492
rect 27249 10489 27261 10492
rect 27295 10520 27307 10523
rect 27295 10492 28948 10520
rect 27295 10489 27307 10492
rect 27249 10483 27307 10489
rect 23992 10424 25820 10452
rect 23992 10412 23998 10424
rect 25866 10412 25872 10464
rect 25924 10412 25930 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 5169 10251 5227 10257
rect 1636 10220 5120 10248
rect 1636 10208 1642 10220
rect 1854 10140 1860 10192
rect 1912 10140 1918 10192
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 2363 10152 2636 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 1872 10112 1900 10140
rect 1872 10084 1992 10112
rect 1578 10004 1584 10056
rect 1636 10004 1642 10056
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1964 10044 1992 10084
rect 2608 10053 2636 10152
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 2740 10084 3188 10112
rect 2740 10072 2746 10084
rect 2409 10047 2467 10053
rect 2409 10044 2421 10047
rect 1964 10016 2421 10044
rect 1857 10007 1915 10013
rect 2409 10013 2421 10016
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 1872 9976 1900 10007
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3160 10053 3188 10084
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10013 3203 10047
rect 3145 10007 3203 10013
rect 3786 10004 3792 10056
rect 3844 10004 3850 10056
rect 5092 10044 5120 10220
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5258 10248 5264 10260
rect 5215 10220 5264 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 6178 10248 6184 10260
rect 5767 10220 6184 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7340 10220 7573 10248
rect 7340 10208 7346 10220
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7561 10211 7619 10217
rect 9214 10208 9220 10260
rect 9272 10208 9278 10260
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 10965 10251 11023 10257
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11238 10248 11244 10260
rect 11011 10220 11244 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 5626 10140 5632 10192
rect 5684 10140 5690 10192
rect 5810 10140 5816 10192
rect 5868 10140 5874 10192
rect 7469 10183 7527 10189
rect 7469 10149 7481 10183
rect 7515 10180 7527 10183
rect 7650 10180 7656 10192
rect 7515 10152 7656 10180
rect 7515 10149 7527 10152
rect 7469 10143 7527 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5224 10084 9168 10112
rect 5224 10072 5230 10084
rect 5092 10016 5396 10044
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 1872 9948 2697 9976
rect 2685 9945 2697 9948
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 2869 9979 2927 9985
rect 2869 9976 2881 9979
rect 2832 9948 2881 9976
rect 2832 9936 2838 9948
rect 2869 9945 2881 9948
rect 2915 9945 2927 9979
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 2869 9939 2927 9945
rect 2976 9948 4046 9976
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2976 9908 3004 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 4034 9939 4092 9945
rect 4890 9936 4896 9988
rect 4948 9976 4954 9988
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 4948 9948 5273 9976
rect 4948 9936 4954 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 5368 9976 5396 10016
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5776 10016 6009 10044
rect 5776 10004 5782 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 8754 10044 8760 10056
rect 5997 10007 6055 10013
rect 6104 10016 8760 10044
rect 6104 9976 6132 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 5368 9948 6132 9976
rect 7101 9979 7159 9985
rect 5261 9939 5319 9945
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7374 9976 7380 9988
rect 7147 9948 7380 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 2087 9880 3004 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 3108 9880 3341 9908
rect 3108 9868 3114 9880
rect 3329 9877 3341 9880
rect 3375 9908 3387 9911
rect 4908 9908 4936 9936
rect 3375 9880 4936 9908
rect 5276 9908 5304 9939
rect 7116 9908 7144 9939
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 9030 9936 9036 9988
rect 9088 9936 9094 9988
rect 9140 9976 9168 10084
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9324 10053 9352 10208
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 10796 10044 10824 10211
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14332 10220 14657 10248
rect 14332 10208 14338 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15436 10220 15485 10248
rect 15436 10208 15442 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15620 10220 15761 10248
rect 15620 10208 15626 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 18230 10248 18236 10260
rect 15896 10220 18236 10248
rect 15896 10208 15902 10220
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 20346 10208 20352 10260
rect 20404 10248 20410 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 20404 10220 20453 10248
rect 20404 10208 20410 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 20441 10211 20499 10217
rect 20622 10208 20628 10260
rect 20680 10208 20686 10260
rect 22186 10208 22192 10260
rect 22244 10208 22250 10260
rect 22373 10251 22431 10257
rect 22373 10217 22385 10251
rect 22419 10248 22431 10251
rect 23198 10248 23204 10260
rect 22419 10220 23204 10248
rect 22419 10217 22431 10220
rect 22373 10211 22431 10217
rect 23198 10208 23204 10220
rect 23256 10248 23262 10260
rect 23658 10248 23664 10260
rect 23256 10220 23664 10248
rect 23256 10208 23262 10220
rect 23658 10208 23664 10220
rect 23716 10208 23722 10260
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 24268 10220 24409 10248
rect 24268 10208 24274 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 26234 10248 26240 10260
rect 24397 10211 24455 10217
rect 25608 10220 26240 10248
rect 11974 10140 11980 10192
rect 12032 10140 12038 10192
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10081 12219 10115
rect 13004 10112 13032 10208
rect 14458 10140 14464 10192
rect 14516 10140 14522 10192
rect 23569 10183 23627 10189
rect 16500 10152 17908 10180
rect 16500 10112 16528 10152
rect 13004 10084 16528 10112
rect 12161 10075 12219 10081
rect 9309 10007 9367 10013
rect 9416 10016 10824 10044
rect 12176 10044 12204 10075
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 16669 10115 16727 10121
rect 16669 10112 16681 10115
rect 16632 10084 16681 10112
rect 16632 10072 16638 10084
rect 16669 10081 16681 10084
rect 16715 10112 16727 10115
rect 17770 10112 17776 10124
rect 16715 10084 17776 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 17880 10112 17908 10152
rect 23569 10149 23581 10183
rect 23615 10180 23627 10183
rect 23750 10180 23756 10192
rect 23615 10152 23756 10180
rect 23615 10149 23627 10152
rect 23569 10143 23627 10149
rect 23750 10140 23756 10152
rect 23808 10140 23814 10192
rect 23860 10112 23888 10208
rect 24946 10140 24952 10192
rect 25004 10180 25010 10192
rect 25608 10180 25636 10220
rect 26234 10208 26240 10220
rect 26292 10248 26298 10260
rect 28537 10251 28595 10257
rect 26292 10220 27200 10248
rect 26292 10208 26298 10220
rect 25004 10152 25636 10180
rect 25004 10140 25010 10152
rect 24486 10112 24492 10124
rect 17880 10084 20852 10112
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12176 10016 12265 10044
rect 9416 9976 9444 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13412 10016 14197 10044
rect 13412 10004 13418 10016
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 9140 9948 9444 9976
rect 9582 9936 9588 9988
rect 9640 9936 9646 9988
rect 10597 9979 10655 9985
rect 10597 9945 10609 9979
rect 10643 9976 10655 9979
rect 10962 9976 10968 9988
rect 10643 9948 10968 9976
rect 10643 9945 10655 9948
rect 10597 9939 10655 9945
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9976 11759 9979
rect 12066 9976 12072 9988
rect 11747 9948 12072 9976
rect 11747 9945 11759 9948
rect 11701 9939 11759 9945
rect 12066 9936 12072 9948
rect 12124 9976 12130 9988
rect 13372 9976 13400 10004
rect 12124 9948 13400 9976
rect 14200 9976 14228 10007
rect 15838 10004 15844 10056
rect 15896 10004 15902 10056
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 16114 10004 16120 10056
rect 16172 10040 16178 10056
rect 16209 10047 16267 10053
rect 16209 10040 16221 10047
rect 16172 10013 16221 10040
rect 16255 10013 16267 10047
rect 17126 10044 17132 10056
rect 16172 10012 16267 10013
rect 16172 10004 16178 10012
rect 16209 10007 16267 10012
rect 16776 10016 17132 10044
rect 16776 9976 16804 10016
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 17218 10004 17224 10056
rect 17276 10004 17282 10056
rect 19444 10016 20668 10044
rect 14200 9948 16804 9976
rect 12124 9936 12130 9948
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 17678 9936 17684 9988
rect 17736 9976 17742 9988
rect 19334 9976 19340 9988
rect 17736 9948 19340 9976
rect 17736 9936 17742 9948
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 19444 9985 19472 10016
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9945 19487 9979
rect 19429 9939 19487 9945
rect 19610 9936 19616 9988
rect 19668 9936 19674 9988
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 20257 9979 20315 9985
rect 20257 9976 20269 9979
rect 19944 9948 20269 9976
rect 19944 9936 19950 9948
rect 20257 9945 20269 9948
rect 20303 9945 20315 9979
rect 20257 9939 20315 9945
rect 5276 9880 7144 9908
rect 9600 9908 9628 9936
rect 10797 9911 10855 9917
rect 10797 9908 10809 9911
rect 9600 9880 10809 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 10797 9877 10809 9880
rect 10843 9877 10855 9911
rect 10797 9871 10855 9877
rect 12434 9868 12440 9920
rect 12492 9868 12498 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16942 9908 16948 9920
rect 16163 9880 16948 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17034 9868 17040 9920
rect 17092 9868 17098 9920
rect 19242 9868 19248 9920
rect 19300 9868 19306 9920
rect 19352 9908 19380 9936
rect 20438 9908 20444 9920
rect 20496 9917 20502 9920
rect 20496 9911 20515 9917
rect 19352 9880 20444 9908
rect 20438 9868 20444 9880
rect 20503 9877 20515 9911
rect 20640 9908 20668 10016
rect 20714 10004 20720 10056
rect 20772 10004 20778 10056
rect 20824 10044 20852 10084
rect 22066 10084 23336 10112
rect 22066 10044 22094 10084
rect 23308 10053 23336 10084
rect 23768 10084 23888 10112
rect 24044 10084 24492 10112
rect 22833 10047 22891 10053
rect 22833 10044 22845 10047
rect 20824 10016 22094 10044
rect 22664 10016 22845 10044
rect 22664 9988 22692 10016
rect 22833 10013 22845 10016
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 23017 10047 23075 10053
rect 23017 10013 23029 10047
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10013 23351 10047
rect 23293 10007 23351 10013
rect 20984 9979 21042 9985
rect 20984 9945 20996 9979
rect 21030 9976 21042 9979
rect 21174 9976 21180 9988
rect 21030 9948 21180 9976
rect 21030 9945 21042 9948
rect 20984 9939 21042 9945
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 22557 9979 22615 9985
rect 22557 9945 22569 9979
rect 22603 9976 22615 9979
rect 22646 9976 22652 9988
rect 22603 9948 22652 9976
rect 22603 9945 22615 9948
rect 22557 9939 22615 9945
rect 22646 9936 22652 9948
rect 22704 9936 22710 9988
rect 21634 9908 21640 9920
rect 20640 9880 21640 9908
rect 20496 9871 20515 9877
rect 20496 9868 20502 9871
rect 21634 9868 21640 9880
rect 21692 9908 21698 9920
rect 22097 9911 22155 9917
rect 22097 9908 22109 9911
rect 21692 9880 22109 9908
rect 21692 9868 21698 9880
rect 22097 9877 22109 9880
rect 22143 9877 22155 9911
rect 22097 9871 22155 9877
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 22370 9917 22376 9920
rect 22347 9911 22376 9917
rect 22347 9908 22359 9911
rect 22244 9880 22359 9908
rect 22244 9868 22250 9880
rect 22347 9877 22359 9880
rect 22347 9871 22376 9877
rect 22370 9868 22376 9871
rect 22428 9868 22434 9920
rect 22830 9868 22836 9920
rect 22888 9908 22894 9920
rect 23032 9908 23060 10007
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23768 10053 23796 10084
rect 23753 10047 23811 10053
rect 23753 10013 23765 10047
rect 23799 10013 23811 10047
rect 23753 10007 23811 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 23934 10044 23940 10056
rect 23891 10016 23940 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 24044 10053 24072 10084
rect 24486 10072 24492 10084
rect 24544 10112 24550 10124
rect 25608 10121 25636 10152
rect 27172 10121 27200 10220
rect 28537 10217 28549 10251
rect 28583 10248 28595 10251
rect 28920 10248 28948 10492
rect 28583 10220 28948 10248
rect 28583 10217 28595 10220
rect 28537 10211 28595 10217
rect 25593 10115 25651 10121
rect 24544 10084 24716 10112
rect 24544 10072 24550 10084
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24029 10007 24087 10013
rect 24135 10016 24593 10044
rect 23201 9979 23259 9985
rect 23201 9945 23213 9979
rect 23247 9976 23259 9979
rect 24044 9976 24072 10007
rect 23247 9948 24072 9976
rect 23247 9945 23259 9948
rect 23201 9939 23259 9945
rect 22888 9880 23060 9908
rect 22888 9868 22894 9880
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24135 9908 24163 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24688 10044 24716 10084
rect 25593 10081 25605 10115
rect 25639 10081 25651 10115
rect 25593 10075 25651 10081
rect 27157 10115 27215 10121
rect 27157 10081 27169 10115
rect 27203 10081 27215 10115
rect 27157 10075 27215 10081
rect 25866 10053 25872 10056
rect 24883 10047 24941 10053
rect 24883 10044 24895 10047
rect 24688 10016 24895 10044
rect 24581 10007 24639 10013
rect 24883 10013 24895 10016
rect 24929 10013 24941 10047
rect 24883 10007 24941 10013
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10013 25099 10047
rect 25860 10044 25872 10053
rect 25827 10016 25872 10044
rect 25041 10007 25099 10013
rect 25860 10007 25872 10016
rect 24673 9979 24731 9985
rect 24673 9976 24685 9979
rect 24596 9948 24685 9976
rect 24596 9920 24624 9948
rect 24673 9945 24685 9948
rect 24719 9945 24731 9979
rect 24673 9939 24731 9945
rect 24762 9936 24768 9988
rect 24820 9936 24826 9988
rect 24084 9880 24163 9908
rect 24084 9868 24090 9880
rect 24578 9868 24584 9920
rect 24636 9868 24642 9920
rect 25056 9908 25084 10007
rect 25866 10004 25872 10007
rect 25924 10004 25930 10056
rect 27424 9979 27482 9985
rect 27424 9945 27436 9979
rect 27470 9976 27482 9979
rect 27522 9976 27528 9988
rect 27470 9948 27528 9976
rect 27470 9945 27482 9948
rect 27424 9939 27482 9945
rect 27522 9936 27528 9948
rect 27580 9936 27586 9988
rect 26973 9911 27031 9917
rect 26973 9908 26985 9911
rect 25056 9880 26985 9908
rect 26973 9877 26985 9880
rect 27019 9908 27031 9911
rect 27246 9908 27252 9920
rect 27019 9880 27252 9908
rect 27019 9877 27031 9880
rect 26973 9871 27031 9877
rect 27246 9868 27252 9880
rect 27304 9868 27310 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 1854 9664 1860 9716
rect 1912 9664 1918 9716
rect 10597 9707 10655 9713
rect 10597 9673 10609 9707
rect 10643 9704 10655 9707
rect 10870 9704 10876 9716
rect 10643 9676 10876 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14458 9704 14464 9716
rect 14231 9676 14464 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14458 9664 14464 9676
rect 14516 9704 14522 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14516 9676 14933 9704
rect 14516 9664 14522 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 16114 9704 16120 9716
rect 14921 9667 14979 9673
rect 15212 9676 16120 9704
rect 1486 9636 1492 9648
rect 1412 9608 1492 9636
rect 1412 9577 1440 9608
rect 1486 9596 1492 9608
rect 1544 9636 1550 9648
rect 1872 9636 1900 9664
rect 2038 9636 2044 9648
rect 1544 9608 2044 9636
rect 1544 9596 1550 9608
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1688 9577 1716 9608
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 5068 9639 5126 9645
rect 5068 9605 5080 9639
rect 5114 9636 5126 9639
rect 5810 9636 5816 9648
rect 5114 9608 5816 9636
rect 5114 9605 5126 9608
rect 5068 9599 5126 9605
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 10321 9639 10379 9645
rect 8812 9608 10088 9636
rect 8812 9596 8818 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2130 9568 2136 9580
rect 1903 9540 2136 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2682 9568 2688 9580
rect 2271 9540 2688 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2240 9500 2268 9531
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3651 9540 3709 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5902 9568 5908 9580
rect 4847 9540 5908 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 2148 9472 2268 9500
rect 2148 9376 2176 9472
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 2498 9432 2504 9444
rect 2455 9404 2504 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 2498 9392 2504 9404
rect 2556 9432 2562 9444
rect 2556 9404 3004 9432
rect 2556 9392 2562 9404
rect 1946 9324 1952 9376
rect 2004 9324 2010 9376
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 2590 9324 2596 9376
rect 2648 9324 2654 9376
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 2976 9364 3004 9404
rect 3602 9364 3608 9376
rect 2976 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 3712 9364 3740 9531
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 3881 9435 3939 9441
rect 3881 9432 3893 9435
rect 3844 9404 3893 9432
rect 3844 9392 3850 9404
rect 3881 9401 3893 9404
rect 3927 9432 3939 9435
rect 4816 9432 4844 9531
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7800 9540 8125 9568
rect 7800 9528 7806 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10060 9577 10088 9608
rect 10321 9605 10333 9639
rect 10367 9636 10379 9639
rect 13170 9636 13176 9648
rect 10367 9608 13176 9636
rect 10367 9605 10379 9608
rect 10321 9599 10379 9605
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 13446 9596 13452 9648
rect 13504 9636 13510 9648
rect 15212 9636 15240 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 16574 9704 16580 9716
rect 16408 9676 16580 9704
rect 15286 9645 15292 9648
rect 13504 9608 15240 9636
rect 13504 9596 13510 9608
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9916 9540 9965 9568
rect 9916 9528 9922 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10046 9571 10104 9577
rect 10046 9537 10058 9571
rect 10092 9537 10104 9571
rect 10046 9531 10104 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10459 9571 10517 9577
rect 10275 9540 10364 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 6086 9500 6092 9512
rect 3927 9404 4844 9432
rect 5828 9472 6092 9500
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 5828 9364 5856 9472
rect 6086 9460 6092 9472
rect 6144 9500 6150 9512
rect 10336 9500 10364 9540
rect 10459 9537 10471 9571
rect 10505 9568 10517 9571
rect 10594 9568 10600 9580
rect 10505 9540 10600 9568
rect 10505 9537 10517 9540
rect 10459 9531 10517 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 11238 9528 11244 9580
rect 11296 9528 11302 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 12526 9568 12532 9580
rect 11517 9531 11575 9537
rect 11716 9540 12532 9568
rect 11256 9500 11284 9528
rect 6144 9472 9720 9500
rect 10336 9472 11284 9500
rect 6144 9460 6150 9472
rect 6181 9435 6239 9441
rect 6181 9401 6193 9435
rect 6227 9432 6239 9435
rect 6638 9432 6644 9444
rect 6227 9404 6644 9432
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 6638 9392 6644 9404
rect 6696 9432 6702 9444
rect 9692 9432 9720 9472
rect 11532 9432 11560 9531
rect 11716 9441 11744 9540
rect 12526 9528 12532 9540
rect 12584 9568 12590 9580
rect 12802 9568 12808 9580
rect 12584 9540 12808 9568
rect 12584 9528 12590 9540
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13061 9571 13119 9577
rect 13061 9568 13073 9571
rect 12952 9540 13073 9568
rect 12952 9528 12958 9540
rect 13061 9537 13073 9540
rect 13107 9537 13119 9571
rect 13061 9531 13119 9537
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 14458 9568 14464 9580
rect 14240 9540 14464 9568
rect 14240 9528 14246 9540
rect 14458 9528 14464 9540
rect 14516 9568 14522 9580
rect 15013 9571 15071 9577
rect 14516 9540 14964 9568
rect 14516 9528 14522 9540
rect 12066 9460 12072 9512
rect 12124 9460 12130 9512
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 14642 9500 14648 9512
rect 14599 9472 14648 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14936 9500 14964 9540
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15212 9568 15240 9608
rect 15273 9639 15292 9645
rect 15273 9605 15285 9639
rect 15273 9599 15292 9605
rect 15286 9596 15292 9599
rect 15344 9596 15350 9648
rect 15473 9639 15531 9645
rect 15473 9605 15485 9639
rect 15519 9605 15531 9639
rect 16408 9636 16436 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 17218 9704 17224 9716
rect 16868 9676 17224 9704
rect 15473 9599 15531 9605
rect 16040 9608 16436 9636
rect 16485 9639 16543 9645
rect 15059 9540 15240 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15488 9500 15516 9599
rect 16040 9577 16068 9608
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 16868 9636 16896 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18049 9707 18107 9713
rect 18049 9704 18061 9707
rect 18012 9676 18061 9704
rect 18012 9664 18018 9676
rect 18049 9673 18061 9676
rect 18095 9673 18107 9707
rect 18049 9667 18107 9673
rect 20346 9664 20352 9716
rect 20404 9704 20410 9716
rect 20714 9704 20720 9716
rect 20404 9676 20720 9704
rect 20404 9664 20410 9676
rect 20714 9664 20720 9676
rect 20772 9704 20778 9716
rect 21085 9707 21143 9713
rect 21085 9704 21097 9707
rect 20772 9676 21097 9704
rect 20772 9664 20778 9676
rect 21085 9673 21097 9676
rect 21131 9673 21143 9707
rect 21085 9667 21143 9673
rect 21174 9664 21180 9716
rect 21232 9664 21238 9716
rect 21266 9664 21272 9716
rect 21324 9664 21330 9716
rect 22189 9707 22247 9713
rect 22189 9673 22201 9707
rect 22235 9704 22247 9707
rect 22462 9704 22468 9716
rect 22235 9676 22468 9704
rect 22235 9673 22247 9676
rect 22189 9667 22247 9673
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 23017 9707 23075 9713
rect 23017 9704 23029 9707
rect 22980 9676 23029 9704
rect 22980 9664 22986 9676
rect 23017 9673 23029 9676
rect 23063 9704 23075 9707
rect 24762 9704 24768 9716
rect 23063 9676 24768 9704
rect 23063 9673 23075 9676
rect 23017 9667 23075 9673
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 27522 9664 27528 9716
rect 27580 9664 27586 9716
rect 16531 9608 16896 9636
rect 16936 9639 16994 9645
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 16936 9605 16948 9639
rect 16982 9636 16994 9639
rect 17034 9636 17040 9648
rect 16982 9608 17040 9636
rect 16982 9605 16994 9608
rect 16936 9599 16994 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 17770 9596 17776 9648
rect 17828 9636 17834 9648
rect 17828 9608 20760 9636
rect 17828 9596 17834 9608
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16347 9540 18276 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16206 9500 16212 9512
rect 14936 9472 16212 9500
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 6696 9404 9628 9432
rect 9692 9404 11560 9432
rect 11701 9435 11759 9441
rect 6696 9392 6702 9404
rect 9600 9376 9628 9404
rect 11701 9401 11713 9435
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 11974 9392 11980 9444
rect 12032 9432 12038 9444
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 12032 9404 12357 9432
rect 12032 9392 12038 9404
rect 12345 9401 12357 9404
rect 12391 9401 12403 9435
rect 16316 9432 16344 9531
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 12345 9395 12403 9401
rect 12452 9404 12848 9432
rect 3712 9336 5856 9364
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 7926 9324 7932 9376
rect 7984 9324 7990 9376
rect 9582 9324 9588 9376
rect 9640 9324 9646 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 10686 9364 10692 9376
rect 9732 9336 10692 9364
rect 9732 9324 9738 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 12452 9364 12480 9404
rect 11020 9336 12480 9364
rect 11020 9324 11026 9336
rect 12526 9324 12532 9376
rect 12584 9324 12590 9376
rect 12820 9364 12848 9404
rect 15304 9404 16344 9432
rect 14182 9364 14188 9376
rect 12820 9336 14188 9364
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14274 9324 14280 9376
rect 14332 9324 14338 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 15304 9373 15332 9404
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 14608 9336 14657 9364
rect 14608 9324 14614 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14645 9327 14703 9333
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 14783 9336 15117 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16022 9364 16028 9376
rect 15887 9336 16028 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16022 9324 16028 9336
rect 16080 9364 16086 9376
rect 16684 9364 16712 9463
rect 18248 9441 18276 9540
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19346 9571 19404 9577
rect 19346 9568 19358 9571
rect 19024 9540 19358 9568
rect 19024 9528 19030 9540
rect 19346 9537 19358 9540
rect 19392 9537 19404 9571
rect 19346 9531 19404 9537
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 19961 9571 20019 9577
rect 19961 9568 19973 9571
rect 19576 9540 19973 9568
rect 19576 9528 19582 9540
rect 19961 9537 19973 9540
rect 20007 9537 20019 9571
rect 19961 9531 20019 9537
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19659 9472 19717 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 20732 9500 20760 9608
rect 21284 9568 21312 9664
rect 21726 9596 21732 9648
rect 21784 9636 21790 9648
rect 21821 9639 21879 9645
rect 21821 9636 21833 9639
rect 21784 9608 21833 9636
rect 21784 9596 21790 9608
rect 21821 9605 21833 9608
rect 21867 9605 21879 9639
rect 21821 9599 21879 9605
rect 22002 9596 22008 9648
rect 22060 9645 22066 9648
rect 22060 9639 22079 9645
rect 22067 9605 22079 9639
rect 22060 9599 22079 9605
rect 22060 9596 22066 9599
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 22940 9636 22968 9664
rect 22428 9608 22968 9636
rect 22428 9596 22434 9608
rect 24118 9596 24124 9648
rect 24176 9636 24182 9648
rect 24581 9639 24639 9645
rect 24581 9636 24593 9639
rect 24176 9608 24593 9636
rect 24176 9596 24182 9608
rect 24581 9605 24593 9608
rect 24627 9605 24639 9639
rect 24581 9599 24639 9605
rect 26878 9596 26884 9648
rect 26936 9636 26942 9648
rect 26973 9639 27031 9645
rect 26973 9636 26985 9639
rect 26936 9608 26985 9636
rect 26936 9596 26942 9608
rect 26973 9605 26985 9608
rect 27019 9605 27031 9639
rect 26973 9599 27031 9605
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21284 9540 21373 9568
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 22646 9528 22652 9580
rect 22704 9568 22710 9580
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 22704 9540 22937 9568
rect 22704 9528 22710 9540
rect 22925 9537 22937 9540
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 24136 9500 24164 9596
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 20732 9472 24164 9500
rect 27433 9503 27491 9509
rect 19705 9463 19763 9469
rect 27433 9469 27445 9503
rect 27479 9500 27491 9503
rect 27724 9500 27752 9531
rect 27479 9472 27752 9500
rect 27479 9469 27491 9472
rect 27433 9463 27491 9469
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 19720 9364 19748 9463
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 22830 9432 22836 9444
rect 21140 9404 22836 9432
rect 21140 9392 21146 9404
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 27246 9392 27252 9444
rect 27304 9392 27310 9444
rect 20622 9364 20628 9376
rect 16080 9336 20628 9364
rect 16080 9324 16086 9336
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 21174 9324 21180 9376
rect 21232 9364 21238 9376
rect 21450 9364 21456 9376
rect 21232 9336 21456 9364
rect 21232 9324 21238 9336
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 21634 9324 21640 9376
rect 21692 9364 21698 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21692 9336 22017 9364
rect 21692 9324 21698 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 24673 9367 24731 9373
rect 24673 9333 24685 9367
rect 24719 9364 24731 9367
rect 24946 9364 24952 9376
rect 24719 9336 24952 9364
rect 24719 9333 24731 9336
rect 24673 9327 24731 9333
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 1946 9120 1952 9172
rect 2004 9120 2010 9172
rect 2590 9120 2596 9172
rect 2648 9120 2654 9172
rect 2866 9160 2872 9172
rect 2746 9132 2872 9160
rect 1964 9024 1992 9120
rect 2608 9024 2636 9120
rect 1688 8996 1992 9024
rect 2240 8996 2636 9024
rect 1486 8916 1492 8968
rect 1544 8916 1550 8968
rect 1688 8965 1716 8996
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1765 8919 1823 8925
rect 1872 8928 1961 8956
rect 1504 8888 1532 8916
rect 1780 8888 1808 8919
rect 1504 8860 1808 8888
rect 1872 8820 1900 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2038 8916 2044 8968
rect 2096 8916 2102 8968
rect 2240 8965 2268 8996
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2547 8928 2605 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2593 8925 2605 8928
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2056 8888 2084 8916
rect 2332 8888 2360 8919
rect 2056 8860 2360 8888
rect 2746 8820 2774 9132
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3436 9132 5672 9160
rect 3436 8965 3464 9132
rect 5644 9092 5672 9132
rect 5718 9120 5724 9172
rect 5776 9120 5782 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 5920 9132 7297 9160
rect 5920 9092 5948 9132
rect 7285 9129 7297 9132
rect 7331 9160 7343 9163
rect 7331 9132 8708 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 5644 9064 5948 9092
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 3752 8996 3924 9024
rect 3752 8984 3758 8996
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3007 8928 3249 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8952 3663 8959
rect 3712 8952 3740 8984
rect 3651 8925 3740 8952
rect 3605 8924 3740 8925
rect 3605 8919 3663 8924
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 3896 8956 3924 8996
rect 5902 8984 5908 9036
rect 5960 8984 5966 9036
rect 8680 9024 8708 9132
rect 8754 9120 8760 9172
rect 8812 9120 8818 9172
rect 9582 9120 9588 9172
rect 9640 9120 9646 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9160 9827 9163
rect 9858 9160 9864 9172
rect 9815 9132 9864 9160
rect 9815 9129 9827 9132
rect 9769 9123 9827 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10376 9132 10609 9160
rect 10376 9120 10382 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 10226 9052 10232 9104
rect 10284 9052 10290 9104
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 10888 9092 10916 9123
rect 12250 9120 12256 9172
rect 12308 9160 12314 9172
rect 12308 9132 12848 9160
rect 12308 9120 12314 9132
rect 10560 9064 10916 9092
rect 10560 9052 10566 9064
rect 12526 9052 12532 9104
rect 12584 9052 12590 9104
rect 12820 9092 12848 9132
rect 12894 9120 12900 9172
rect 12952 9120 12958 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 14274 9160 14280 9172
rect 13403 9132 14280 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14734 9120 14740 9172
rect 14792 9120 14798 9172
rect 15194 9120 15200 9172
rect 15252 9120 15258 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15344 9132 15669 9160
rect 15344 9120 15350 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 15930 9160 15936 9172
rect 15887 9132 15936 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 16080 9132 16129 9160
rect 16080 9120 16086 9132
rect 16117 9129 16129 9132
rect 16163 9129 16175 9163
rect 16117 9123 16175 9129
rect 16206 9120 16212 9172
rect 16264 9120 16270 9172
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16724 9132 16957 9160
rect 16724 9120 16730 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 17129 9163 17187 9169
rect 17129 9129 17141 9163
rect 17175 9160 17187 9163
rect 18138 9160 18144 9172
rect 17175 9132 18144 9160
rect 17175 9129 17187 9132
rect 17129 9123 17187 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18966 9120 18972 9172
rect 19024 9120 19030 9172
rect 19518 9120 19524 9172
rect 19576 9120 19582 9172
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22833 9163 22891 9169
rect 22833 9160 22845 9163
rect 22520 9132 22845 9160
rect 22520 9120 22526 9132
rect 22833 9129 22845 9132
rect 22879 9129 22891 9163
rect 22833 9123 22891 9129
rect 23014 9120 23020 9172
rect 23072 9120 23078 9172
rect 23569 9163 23627 9169
rect 23569 9129 23581 9163
rect 23615 9129 23627 9163
rect 23569 9123 23627 9129
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 12820 9064 13553 9092
rect 13541 9061 13553 9064
rect 13587 9061 13599 9095
rect 13541 9055 13599 9061
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14550 9092 14556 9104
rect 14240 9064 14556 9092
rect 14240 9052 14246 9064
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 14752 9092 14780 9120
rect 15381 9095 15439 9101
rect 15381 9092 15393 9095
rect 14752 9064 15393 9092
rect 15381 9061 15393 9064
rect 15427 9061 15439 9095
rect 16224 9092 16252 9120
rect 17218 9092 17224 9104
rect 16224 9064 17224 9092
rect 15381 9055 15439 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 17954 9052 17960 9104
rect 18012 9052 18018 9104
rect 18693 9095 18751 9101
rect 18064 9064 18644 9092
rect 9858 9024 9864 9036
rect 8680 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 9950 8984 9956 9036
rect 10008 8984 10014 9036
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 3896 8928 5365 8956
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 4034 8891 4092 8897
rect 4034 8888 4046 8891
rect 3712 8860 4046 8888
rect 1872 8792 2774 8820
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3712 8820 3740 8860
rect 4034 8857 4046 8860
rect 4080 8857 4092 8891
rect 4034 8851 4092 8857
rect 5537 8891 5595 8897
rect 5537 8857 5549 8891
rect 5583 8888 5595 8891
rect 5810 8888 5816 8900
rect 5583 8860 5816 8888
rect 5583 8857 5595 8860
rect 5537 8851 5595 8857
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 5920 8888 5948 8984
rect 6172 8959 6230 8965
rect 6172 8925 6184 8959
rect 6218 8956 6230 8959
rect 6546 8956 6552 8968
rect 6218 8928 6552 8956
rect 6218 8925 6230 8928
rect 6172 8919 6230 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7644 8959 7702 8965
rect 7644 8925 7656 8959
rect 7690 8956 7702 8959
rect 7926 8956 7932 8968
rect 7690 8928 7932 8956
rect 7690 8925 7702 8928
rect 7644 8919 7702 8925
rect 7392 8888 7420 8919
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 10235 8965 10263 9052
rect 12544 9024 12572 9052
rect 10428 8996 11100 9024
rect 12544 8996 12756 9024
rect 10428 8965 10456 8996
rect 10091 8959 10149 8965
rect 10091 8934 10103 8959
rect 10060 8925 10103 8934
rect 10137 8925 10149 8959
rect 10060 8922 10149 8925
rect 9968 8919 10149 8922
rect 10204 8959 10263 8965
rect 10204 8925 10216 8959
rect 10250 8928 10263 8959
rect 10413 8959 10471 8965
rect 10250 8925 10262 8928
rect 10204 8919 10262 8925
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 9968 8906 10134 8919
rect 10594 8916 10600 8968
rect 10652 8916 10658 8968
rect 5920 8860 7420 8888
rect 9122 8848 9128 8900
rect 9180 8888 9186 8900
rect 9674 8897 9680 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 9180 8860 9413 8888
rect 9180 8848 9186 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9401 8851 9459 8857
rect 9617 8891 9680 8897
rect 9617 8857 9629 8891
rect 9663 8857 9680 8891
rect 9617 8851 9680 8857
rect 9674 8848 9680 8851
rect 9732 8848 9738 8900
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 9968 8894 10088 8906
rect 9968 8888 9996 8894
rect 9916 8860 9996 8888
rect 10321 8891 10379 8897
rect 9916 8848 9922 8860
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 10612 8888 10640 8916
rect 10367 8860 10640 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 10686 8848 10692 8900
rect 10744 8848 10750 8900
rect 10904 8897 10932 8996
rect 10889 8891 10947 8897
rect 10889 8857 10901 8891
rect 10935 8857 10947 8891
rect 11072 8888 11100 8996
rect 12273 8959 12331 8965
rect 12273 8925 12285 8959
rect 12319 8956 12331 8959
rect 12434 8956 12440 8968
rect 12319 8928 12440 8956
rect 12319 8925 12331 8928
rect 12273 8919 12331 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 12728 8965 12756 8996
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 18064 9024 18092 9064
rect 13320 8996 18092 9024
rect 18141 9027 18199 9033
rect 13320 8984 13326 8996
rect 18141 8993 18153 9027
rect 18187 9024 18199 9027
rect 18616 9024 18644 9064
rect 18693 9061 18705 9095
rect 18739 9092 18751 9095
rect 19536 9092 19564 9120
rect 22370 9092 22376 9104
rect 18739 9064 19564 9092
rect 19628 9064 22376 9092
rect 18739 9061 18751 9064
rect 18693 9055 18751 9061
rect 19628 9024 19656 9064
rect 22370 9052 22376 9064
rect 22428 9052 22434 9104
rect 23584 9092 23612 9123
rect 23750 9120 23756 9172
rect 23808 9120 23814 9172
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 24412 9132 25789 9160
rect 24412 9092 24440 9132
rect 25777 9129 25789 9132
rect 25823 9129 25835 9163
rect 25777 9123 25835 9129
rect 23584 9064 24440 9092
rect 25792 9092 25820 9123
rect 27614 9120 27620 9172
rect 27672 9160 27678 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 27672 9132 28273 9160
rect 27672 9120 27678 9132
rect 28261 9129 28273 9132
rect 28307 9129 28319 9163
rect 28261 9123 28319 9129
rect 25961 9095 26019 9101
rect 25961 9092 25973 9095
rect 25792 9064 25973 9092
rect 25961 9061 25973 9064
rect 26007 9061 26019 9095
rect 25961 9055 26019 9061
rect 26881 9027 26939 9033
rect 26881 9024 26893 9027
rect 18187 8996 18552 9024
rect 18616 8996 19656 9024
rect 26068 8996 26893 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 12544 8888 12572 8919
rect 12820 8888 12848 8984
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13964 8928 14289 8956
rect 13964 8916 13970 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 11072 8860 12480 8888
rect 12544 8860 12848 8888
rect 10889 8851 10947 8857
rect 3191 8792 3740 8820
rect 5169 8823 5227 8829
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5442 8820 5448 8832
rect 5215 8792 5448 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5442 8780 5448 8792
rect 5500 8820 5506 8832
rect 10502 8820 10508 8832
rect 5500 8792 10508 8820
rect 5500 8780 5506 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 10904 8820 10932 8851
rect 10652 8792 10932 8820
rect 10652 8780 10658 8792
rect 11054 8780 11060 8832
rect 11112 8780 11118 8832
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11974 8820 11980 8832
rect 11195 8792 11980 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 12452 8820 12480 8860
rect 13078 8848 13084 8900
rect 13136 8848 13142 8900
rect 14292 8888 14320 8919
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 15488 8956 15608 8958
rect 14936 8928 15148 8956
rect 14936 8888 14964 8928
rect 14292 8860 14964 8888
rect 15013 8891 15071 8897
rect 15013 8857 15025 8891
rect 15059 8857 15071 8891
rect 15013 8851 15071 8857
rect 12710 8820 12716 8832
rect 12452 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13412 8792 14105 8820
rect 13412 8780 13418 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15028 8820 15056 8851
rect 14792 8792 15056 8820
rect 15120 8820 15148 8928
rect 15488 8930 16344 8956
rect 15488 8900 15516 8930
rect 15580 8928 16344 8930
rect 15229 8891 15287 8897
rect 15229 8857 15241 8891
rect 15275 8888 15287 8891
rect 15378 8888 15384 8900
rect 15275 8860 15384 8888
rect 15275 8857 15287 8860
rect 15229 8851 15287 8857
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 15470 8848 15476 8900
rect 15528 8848 15534 8900
rect 16316 8897 16344 8928
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 18524 8965 18552 8996
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 17184 8928 17693 8956
rect 17184 8916 17190 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 19242 8956 19248 8968
rect 18831 8928 19248 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 20772 8928 20821 8956
rect 20772 8916 20778 8928
rect 20809 8925 20821 8928
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 20993 8959 21051 8965
rect 20993 8925 21005 8959
rect 21039 8956 21051 8959
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21039 8928 21373 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 22738 8916 22744 8968
rect 22796 8956 22802 8968
rect 23290 8956 23296 8968
rect 22796 8928 23296 8956
rect 22796 8916 22802 8928
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 24026 8916 24032 8968
rect 24084 8916 24090 8968
rect 24397 8959 24455 8965
rect 24397 8925 24409 8959
rect 24443 8956 24455 8959
rect 24946 8956 24952 8968
rect 24443 8928 24952 8956
rect 24443 8925 24455 8928
rect 24397 8919 24455 8925
rect 24946 8916 24952 8928
rect 25004 8956 25010 8968
rect 26068 8956 26096 8996
rect 26881 8993 26893 8996
rect 26927 8993 26939 9027
rect 26881 8987 26939 8993
rect 25004 8928 26096 8956
rect 25004 8916 25010 8928
rect 26602 8916 26608 8968
rect 26660 8916 26666 8968
rect 15673 8891 15731 8897
rect 15673 8888 15685 8891
rect 15672 8857 15685 8888
rect 15719 8888 15731 8891
rect 16301 8891 16359 8897
rect 15719 8860 16252 8888
rect 15719 8857 15731 8860
rect 15672 8851 15731 8857
rect 15672 8820 15700 8851
rect 15120 8792 15700 8820
rect 14792 8780 14798 8792
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 16114 8829 16120 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 15896 8792 15945 8820
rect 15896 8780 15902 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 16101 8823 16120 8829
rect 16101 8789 16113 8823
rect 16101 8783 16120 8789
rect 16114 8780 16120 8783
rect 16172 8780 16178 8832
rect 16224 8820 16252 8860
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 16574 8888 16580 8900
rect 16347 8860 16580 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 16758 8848 16764 8900
rect 16816 8888 16822 8900
rect 17494 8888 17500 8900
rect 16816 8860 17500 8888
rect 16816 8848 16822 8860
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 17770 8848 17776 8900
rect 17828 8888 17834 8900
rect 19610 8888 19616 8900
rect 17828 8860 19616 8888
rect 17828 8848 17834 8860
rect 19610 8848 19616 8860
rect 19668 8888 19674 8900
rect 20625 8891 20683 8897
rect 20625 8888 20637 8891
rect 19668 8860 20637 8888
rect 19668 8848 19674 8860
rect 20625 8857 20637 8860
rect 20671 8857 20683 8891
rect 20625 8851 20683 8857
rect 16961 8823 17019 8829
rect 16961 8820 16973 8823
rect 16224 8792 16973 8820
rect 16961 8789 16973 8792
rect 17007 8789 17019 8823
rect 16961 8783 17019 8789
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 19334 8820 19340 8832
rect 17184 8792 19340 8820
rect 17184 8780 17190 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 20640 8820 20668 8851
rect 21450 8848 21456 8900
rect 21508 8848 21514 8900
rect 22646 8848 22652 8900
rect 22704 8888 22710 8900
rect 23385 8891 23443 8897
rect 23385 8888 23397 8891
rect 22704 8860 23397 8888
rect 22704 8848 22710 8860
rect 23385 8857 23397 8860
rect 23431 8888 23443 8891
rect 23750 8888 23756 8900
rect 23431 8860 23756 8888
rect 23431 8857 23443 8860
rect 23385 8851 23443 8857
rect 23750 8848 23756 8860
rect 23808 8848 23814 8900
rect 24642 8891 24700 8897
rect 24642 8888 24654 8891
rect 24228 8860 24654 8888
rect 21468 8820 21496 8848
rect 20640 8792 21496 8820
rect 21542 8780 21548 8832
rect 21600 8780 21606 8832
rect 21634 8780 21640 8832
rect 21692 8820 21698 8832
rect 22664 8820 22692 8848
rect 21692 8792 22692 8820
rect 21692 8780 21698 8792
rect 22830 8780 22836 8832
rect 22888 8829 22894 8832
rect 22888 8823 22907 8829
rect 22895 8789 22907 8823
rect 22888 8783 22907 8789
rect 23595 8823 23653 8829
rect 23595 8789 23607 8823
rect 23641 8820 23653 8823
rect 23934 8820 23940 8832
rect 23641 8792 23940 8820
rect 23641 8789 23653 8792
rect 23595 8783 23653 8789
rect 22888 8780 22894 8783
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 24228 8829 24256 8860
rect 24642 8857 24654 8860
rect 24688 8857 24700 8891
rect 24642 8851 24700 8857
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 26326 8888 26332 8900
rect 24912 8860 26332 8888
rect 24912 8848 24918 8860
rect 26326 8848 26332 8860
rect 26384 8848 26390 8900
rect 27126 8891 27184 8897
rect 27126 8888 27138 8891
rect 26804 8860 27138 8888
rect 24213 8823 24271 8829
rect 24213 8789 24225 8823
rect 24259 8789 24271 8823
rect 24213 8783 24271 8789
rect 25866 8780 25872 8832
rect 25924 8780 25930 8832
rect 26804 8829 26832 8860
rect 27126 8857 27138 8860
rect 27172 8857 27184 8891
rect 27126 8851 27184 8857
rect 26789 8823 26847 8829
rect 26789 8789 26801 8823
rect 26835 8789 26847 8823
rect 26789 8783 26847 8789
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1486 8576 1492 8628
rect 1544 8576 1550 8628
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 2774 8616 2780 8628
rect 1627 8588 2780 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3142 8616 3148 8628
rect 2915 8588 3148 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7800 8588 8033 8616
rect 7800 8576 7806 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8754 8576 8760 8628
rect 8812 8576 8818 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9306 8616 9312 8628
rect 9180 8588 9312 8616
rect 9180 8576 9186 8588
rect 9306 8576 9312 8588
rect 9364 8616 9370 8628
rect 10226 8616 10232 8628
rect 9364 8588 10232 8616
rect 9364 8576 9370 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10870 8616 10876 8628
rect 10928 8625 10934 8628
rect 10928 8619 10947 8625
rect 10468 8588 10876 8616
rect 10468 8576 10474 8588
rect 10870 8576 10876 8588
rect 10935 8585 10947 8619
rect 10928 8579 10947 8585
rect 10928 8576 10934 8579
rect 14642 8576 14648 8628
rect 14700 8576 14706 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 16390 8616 16396 8628
rect 14792 8588 16396 8616
rect 14792 8576 14798 8588
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1504 8480 1532 8576
rect 4154 8508 4160 8560
rect 4212 8508 4218 8560
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1504 8452 1685 8480
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1903 8452 1961 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 3476 8452 5089 8480
rect 3476 8440 3482 8452
rect 5077 8449 5089 8452
rect 5123 8480 5135 8483
rect 5123 8452 5396 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 4798 8372 4804 8424
rect 4856 8372 4862 8424
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5184 8276 5212 8375
rect 5368 8356 5396 8452
rect 5350 8304 5356 8356
rect 5408 8304 5414 8356
rect 5460 8353 5488 8576
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5644 8452 5917 8480
rect 5644 8421 5672 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 5445 8347 5503 8353
rect 5445 8313 5457 8347
rect 5491 8313 5503 8347
rect 6380 8344 6408 8375
rect 6656 8353 6684 8576
rect 7837 8551 7895 8557
rect 7837 8517 7849 8551
rect 7883 8548 7895 8551
rect 8297 8551 8355 8557
rect 7883 8520 8248 8548
rect 7883 8517 7895 8520
rect 7837 8511 7895 8517
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8480 7711 8483
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7699 8452 8125 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8220 8480 8248 8520
rect 8297 8517 8309 8551
rect 8343 8548 8355 8551
rect 8772 8548 8800 8576
rect 8846 8557 8852 8560
rect 8343 8520 8800 8548
rect 8343 8517 8355 8520
rect 8297 8511 8355 8517
rect 8840 8511 8852 8557
rect 8846 8508 8852 8511
rect 8904 8508 8910 8560
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 10594 8548 10600 8560
rect 9732 8520 10600 8548
rect 9732 8508 9738 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8548 10747 8551
rect 10778 8548 10784 8560
rect 10735 8520 10784 8548
rect 10735 8517 10747 8520
rect 10689 8511 10747 8517
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 11885 8551 11943 8557
rect 11885 8517 11897 8551
rect 11931 8548 11943 8551
rect 12066 8548 12072 8560
rect 11931 8520 12072 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 15856 8557 15884 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 17129 8619 17187 8625
rect 16776 8588 17080 8616
rect 14277 8551 14335 8557
rect 14277 8548 14289 8551
rect 14200 8520 14289 8548
rect 10962 8480 10968 8492
rect 8220 8452 10968 8480
rect 8113 8443 8171 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11698 8489 11704 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11112 8452 11529 8480
rect 11112 8440 11118 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11665 8483 11704 8489
rect 11665 8449 11677 8483
rect 11665 8443 11704 8449
rect 11698 8440 11704 8443
rect 11756 8440 11762 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11982 8483 12040 8489
rect 11982 8449 11994 8483
rect 12028 8480 12040 8483
rect 13446 8480 13452 8492
rect 12028 8452 13452 8480
rect 12028 8449 12040 8452
rect 11982 8443 12040 8449
rect 8478 8372 8484 8424
rect 8536 8372 8542 8424
rect 8570 8372 8576 8424
rect 8628 8372 8634 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11238 8412 11244 8424
rect 9916 8384 11244 8412
rect 9916 8372 9922 8384
rect 11238 8372 11244 8384
rect 11296 8412 11302 8424
rect 11808 8412 11836 8443
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 14200 8480 14228 8520
rect 14277 8517 14289 8520
rect 14323 8517 14335 8551
rect 15841 8551 15899 8557
rect 14277 8511 14335 8517
rect 14507 8517 14565 8523
rect 14507 8514 14519 8517
rect 13648 8452 14228 8480
rect 14492 8483 14519 8514
rect 14553 8483 14565 8517
rect 15841 8517 15853 8551
rect 15887 8517 15899 8551
rect 15841 8511 15899 8517
rect 15930 8508 15936 8560
rect 15988 8548 15994 8560
rect 16057 8551 16115 8557
rect 16057 8548 16069 8551
rect 15988 8520 16069 8548
rect 15988 8508 15994 8520
rect 16057 8517 16069 8520
rect 16103 8548 16115 8551
rect 16482 8548 16488 8560
rect 16103 8520 16488 8548
rect 16103 8517 16115 8520
rect 16057 8511 16115 8517
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 16776 8557 16804 8588
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 16632 8520 16773 8548
rect 16632 8508 16638 8520
rect 16761 8517 16773 8520
rect 16807 8517 16819 8551
rect 16761 8511 16819 8517
rect 16942 8508 16948 8560
rect 17000 8557 17006 8560
rect 17000 8551 17019 8557
rect 17007 8517 17019 8551
rect 17052 8548 17080 8588
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17402 8616 17408 8628
rect 17175 8588 17408 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17644 8588 17908 8616
rect 17644 8576 17650 8588
rect 17604 8548 17632 8576
rect 17052 8520 17632 8548
rect 17000 8511 17019 8517
rect 17000 8508 17006 8511
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 17773 8551 17831 8557
rect 17773 8548 17785 8551
rect 17736 8520 17785 8548
rect 17736 8508 17742 8520
rect 17773 8517 17785 8520
rect 17819 8517 17831 8551
rect 17773 8511 17831 8517
rect 14492 8477 14565 8483
rect 13354 8412 13360 8424
rect 11296 8384 13360 8412
rect 11296 8372 11302 8384
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13648 8356 13676 8452
rect 14492 8412 14520 8477
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 14700 8452 17601 8480
rect 14700 8440 14706 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17880 8480 17908 8588
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18216 8588 19334 8616
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 18216 8557 18244 8588
rect 18201 8551 18259 8557
rect 18201 8548 18213 8551
rect 18012 8520 18213 8548
rect 18012 8508 18018 8520
rect 18201 8517 18213 8520
rect 18247 8517 18259 8551
rect 18201 8511 18259 8517
rect 18417 8551 18475 8557
rect 18417 8517 18429 8551
rect 18463 8548 18475 8551
rect 19058 8548 19064 8560
rect 18463 8520 19064 8548
rect 18463 8517 18475 8520
rect 18417 8511 18475 8517
rect 18432 8480 18460 8511
rect 19058 8508 19064 8520
rect 19116 8508 19122 8560
rect 19306 8548 19334 8588
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20599 8619 20657 8625
rect 20599 8616 20611 8619
rect 20036 8588 20611 8616
rect 20036 8576 20042 8588
rect 20599 8585 20611 8588
rect 20645 8585 20657 8619
rect 21174 8616 21180 8628
rect 21232 8625 21238 8628
rect 21232 8619 21251 8625
rect 20599 8579 20657 8585
rect 20732 8588 21180 8616
rect 20732 8548 20760 8588
rect 21174 8576 21180 8588
rect 21239 8585 21251 8619
rect 21232 8579 21251 8585
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 22646 8616 22652 8628
rect 21407 8588 22652 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21232 8576 21238 8579
rect 22646 8576 22652 8588
rect 22704 8576 22710 8628
rect 23201 8619 23259 8625
rect 23201 8585 23213 8619
rect 23247 8585 23259 8619
rect 23201 8579 23259 8585
rect 19306 8520 20760 8548
rect 20809 8551 20867 8557
rect 20809 8517 20821 8551
rect 20855 8517 20867 8551
rect 20809 8511 20867 8517
rect 17880 8452 18460 8480
rect 17589 8443 17647 8449
rect 14492 8384 16160 8412
rect 5445 8307 5503 8313
rect 5644 8316 6408 8344
rect 6641 8347 6699 8353
rect 5644 8288 5672 8316
rect 6641 8313 6653 8347
rect 6687 8313 6699 8347
rect 11057 8347 11115 8353
rect 6641 8307 6699 8313
rect 9876 8316 10456 8344
rect 5626 8276 5632 8288
rect 5184 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 5718 8236 5724 8288
rect 5776 8236 5782 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 9876 8276 9904 8316
rect 6880 8248 9904 8276
rect 6880 8236 6886 8248
rect 9950 8236 9956 8288
rect 10008 8236 10014 8288
rect 10428 8276 10456 8316
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11146 8344 11152 8356
rect 11103 8316 11152 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 12158 8304 12164 8356
rect 12216 8304 12222 8356
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12710 8344 12716 8356
rect 12308 8316 12716 8344
rect 12308 8304 12314 8316
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 13630 8304 13636 8356
rect 13688 8304 13694 8356
rect 16132 8344 16160 8384
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16390 8412 16396 8424
rect 16264 8384 16396 8412
rect 16264 8372 16270 8384
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17604 8412 17632 8443
rect 19794 8440 19800 8492
rect 19852 8440 19858 8492
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 20824 8480 20852 8511
rect 20990 8508 20996 8560
rect 21048 8557 21054 8560
rect 21048 8551 21077 8557
rect 21065 8517 21077 8551
rect 21048 8511 21077 8517
rect 21048 8508 21054 8511
rect 21542 8508 21548 8560
rect 21600 8548 21606 8560
rect 21726 8548 21732 8560
rect 21600 8520 21732 8548
rect 21600 8508 21606 8520
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 22002 8508 22008 8560
rect 22060 8548 22066 8560
rect 22060 8520 22140 8548
rect 22060 8508 22066 8520
rect 22112 8489 22140 8520
rect 20772 8452 20852 8480
rect 22088 8483 22146 8489
rect 20772 8440 20778 8452
rect 22088 8449 22100 8483
rect 22134 8449 22146 8483
rect 22088 8443 22146 8449
rect 20990 8412 20996 8424
rect 17604 8384 20996 8412
rect 20990 8372 20996 8384
rect 21048 8412 21054 8424
rect 21634 8412 21640 8424
rect 21048 8384 21640 8412
rect 21048 8372 21054 8384
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 21818 8372 21824 8424
rect 21876 8372 21882 8424
rect 23216 8412 23244 8579
rect 23290 8576 23296 8628
rect 23348 8576 23354 8628
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23624 8588 23980 8616
rect 23624 8576 23630 8588
rect 23474 8557 23480 8560
rect 23445 8551 23480 8557
rect 23445 8517 23457 8551
rect 23445 8511 23480 8517
rect 23474 8508 23480 8511
rect 23532 8508 23538 8560
rect 23584 8412 23612 8576
rect 23658 8508 23664 8560
rect 23716 8508 23722 8560
rect 23753 8551 23811 8557
rect 23753 8517 23765 8551
rect 23799 8548 23811 8551
rect 23842 8548 23848 8560
rect 23799 8520 23848 8548
rect 23799 8517 23811 8520
rect 23753 8511 23811 8517
rect 23842 8508 23848 8520
rect 23900 8508 23906 8560
rect 23952 8557 23980 8588
rect 24026 8576 24032 8628
rect 24084 8616 24090 8628
rect 24397 8619 24455 8625
rect 24397 8616 24409 8619
rect 24084 8588 24409 8616
rect 24084 8576 24090 8588
rect 24397 8585 24409 8588
rect 24443 8585 24455 8619
rect 24397 8579 24455 8585
rect 24854 8576 24860 8628
rect 24912 8576 24918 8628
rect 25317 8619 25375 8625
rect 25317 8585 25329 8619
rect 25363 8585 25375 8619
rect 25317 8579 25375 8585
rect 23937 8551 23995 8557
rect 23937 8517 23949 8551
rect 23983 8517 23995 8551
rect 23937 8511 23995 8517
rect 24872 8489 24900 8576
rect 25332 8548 25360 8579
rect 25866 8576 25872 8628
rect 25924 8576 25930 8628
rect 26602 8576 26608 8628
rect 26660 8616 26666 8628
rect 26973 8619 27031 8625
rect 26973 8616 26985 8619
rect 26660 8588 26985 8616
rect 26660 8576 26666 8588
rect 26973 8585 26985 8588
rect 27019 8585 27031 8619
rect 26973 8579 27031 8585
rect 25654 8551 25712 8557
rect 25654 8548 25666 8551
rect 25332 8520 25666 8548
rect 25654 8517 25666 8520
rect 25700 8517 25712 8551
rect 25654 8511 25712 8517
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8480 25191 8483
rect 25884 8480 25912 8576
rect 26326 8508 26332 8560
rect 26384 8548 26390 8560
rect 27433 8551 27491 8557
rect 27433 8548 27445 8551
rect 26384 8520 27445 8548
rect 26384 8508 26390 8520
rect 27433 8517 27445 8520
rect 27479 8517 27491 8551
rect 27433 8511 27491 8517
rect 25179 8452 25912 8480
rect 25179 8449 25191 8452
rect 25133 8443 25191 8449
rect 23216 8384 23612 8412
rect 24486 8372 24492 8424
rect 24544 8412 24550 8424
rect 25409 8415 25467 8421
rect 25409 8412 25421 8415
rect 24544 8384 25421 8412
rect 24544 8372 24550 8384
rect 25409 8381 25421 8384
rect 25455 8381 25467 8415
rect 25409 8375 25467 8381
rect 17954 8344 17960 8356
rect 14384 8316 14596 8344
rect 16132 8316 17960 8344
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 10428 8248 10885 8276
rect 10873 8245 10885 8248
rect 10919 8245 10931 8279
rect 10873 8239 10931 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 14384 8276 14412 8316
rect 11020 8248 14412 8276
rect 11020 8236 11026 8248
rect 14458 8236 14464 8288
rect 14516 8236 14522 8288
rect 14568 8276 14596 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 20438 8304 20444 8356
rect 20496 8304 20502 8356
rect 20640 8316 21864 8344
rect 15286 8276 15292 8288
rect 14568 8248 15292 8276
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 16022 8236 16028 8288
rect 16080 8236 16086 8288
rect 16206 8236 16212 8288
rect 16264 8236 16270 8288
rect 16942 8236 16948 8288
rect 17000 8236 17006 8288
rect 18230 8236 18236 8288
rect 18288 8236 18294 8288
rect 19978 8236 19984 8288
rect 20036 8236 20042 8288
rect 20640 8285 20668 8316
rect 20625 8279 20683 8285
rect 20625 8245 20637 8279
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 21836 8276 21864 8316
rect 23216 8316 24532 8344
rect 23216 8276 23244 8316
rect 21836 8248 23244 8276
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23658 8276 23664 8288
rect 23523 8248 23664 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 24118 8236 24124 8288
rect 24176 8236 24182 8288
rect 24504 8276 24532 8316
rect 24578 8304 24584 8356
rect 24636 8304 24642 8356
rect 27065 8347 27123 8353
rect 27065 8344 27077 8347
rect 26804 8316 27077 8344
rect 26804 8285 26832 8316
rect 27065 8313 27077 8316
rect 27111 8313 27123 8347
rect 27065 8307 27123 8313
rect 26789 8279 26847 8285
rect 26789 8276 26801 8279
rect 24504 8248 26801 8276
rect 26789 8245 26801 8248
rect 26835 8245 26847 8279
rect 26789 8239 26847 8245
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3418 8072 3424 8084
rect 3375 8044 3424 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4798 8072 4804 8084
rect 4540 8044 4804 8072
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 4387 7976 4476 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1627 7840 1716 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1688 7800 1716 7840
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2547 7840 2605 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2516 7800 2544 7831
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3068 7800 3096 7831
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 4448 7868 4476 7976
rect 4540 7945 4568 8044
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5828 8044 8340 8072
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 5828 7868 5856 8044
rect 5905 8007 5963 8013
rect 5905 7973 5917 8007
rect 5951 8004 5963 8007
rect 6365 8007 6423 8013
rect 6365 8004 6377 8007
rect 5951 7976 6377 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 6365 7973 6377 7976
rect 6411 8004 6423 8007
rect 8312 8004 8340 8044
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 8941 8035 8999 8041
rect 9048 8044 12265 8072
rect 9048 8004 9076 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 13078 8072 13084 8084
rect 12575 8044 13084 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 14516 8044 15792 8072
rect 14516 8032 14522 8044
rect 6411 7976 8248 8004
rect 8312 7976 9076 8004
rect 6411 7973 6423 7976
rect 6365 7967 6423 7973
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 3476 7840 5856 7868
rect 6472 7868 6500 7899
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 8220 7936 8248 7976
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 10008 7976 10333 8004
rect 10008 7964 10014 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 11054 8004 11060 8016
rect 10321 7967 10379 7973
rect 10704 7976 11060 8004
rect 10226 7936 10232 7948
rect 6696 7908 6776 7936
rect 8220 7908 10232 7936
rect 6696 7896 6702 7908
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6472 7840 6561 7868
rect 3476 7828 3482 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 1688 7772 3096 7800
rect 3237 7803 3295 7809
rect 1688 7744 1716 7772
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 3786 7800 3792 7812
rect 3283 7772 3792 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 3786 7760 3792 7772
rect 3844 7760 3850 7812
rect 3973 7803 4031 7809
rect 3973 7769 3985 7803
rect 4019 7800 4031 7803
rect 4792 7803 4850 7809
rect 4019 7772 4752 7800
rect 4019 7769 4031 7772
rect 3973 7763 4031 7769
rect 1670 7692 1676 7744
rect 1728 7692 1734 7744
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 4724 7732 4752 7772
rect 4792 7769 4804 7803
rect 4838 7800 4850 7803
rect 4890 7800 4896 7812
rect 4838 7772 4896 7800
rect 4838 7769 4850 7772
rect 4792 7763 4850 7769
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 5626 7760 5632 7812
rect 5684 7800 5690 7812
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 5684 7772 6009 7800
rect 5684 7760 5690 7772
rect 5997 7769 6009 7772
rect 6043 7800 6055 7803
rect 6638 7800 6644 7812
rect 6043 7772 6644 7800
rect 6043 7769 6055 7772
rect 5997 7763 6055 7769
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6748 7800 6776 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8536 7840 9137 7868
rect 8536 7828 8542 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10704 7868 10732 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 12437 8007 12495 8013
rect 12437 7973 12449 8007
rect 12483 8004 12495 8007
rect 12805 8007 12863 8013
rect 12805 8004 12817 8007
rect 12483 7976 12817 8004
rect 12483 7973 12495 7976
rect 12437 7967 12495 7973
rect 12805 7973 12817 7976
rect 12851 7973 12863 8007
rect 15764 8004 15792 8044
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16206 8072 16212 8084
rect 16163 8044 16212 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16298 8032 16304 8084
rect 16356 8032 16362 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 17788 8044 19441 8072
rect 17126 8004 17132 8016
rect 15764 7976 17132 8004
rect 12805 7967 12863 7973
rect 17126 7964 17132 7976
rect 17184 8004 17190 8016
rect 17681 8007 17739 8013
rect 17681 8004 17693 8007
rect 17184 7976 17693 8004
rect 17184 7964 17190 7976
rect 17681 7973 17693 7976
rect 17727 7973 17739 8007
rect 17681 7967 17739 7973
rect 12526 7936 12532 7948
rect 10888 7908 12532 7936
rect 10091 7840 10732 7868
rect 10781 7871 10839 7877
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10781 7837 10793 7871
rect 10827 7870 10839 7871
rect 10888 7870 10916 7908
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 17788 7936 17816 8044
rect 19429 8041 19441 8044
rect 19475 8041 19487 8075
rect 19429 8035 19487 8041
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 20070 8072 20076 8084
rect 19659 8044 20076 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 20070 8032 20076 8044
rect 20128 8032 20134 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 21174 8072 21180 8084
rect 21131 8044 21180 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 22465 8075 22523 8081
rect 22465 8041 22477 8075
rect 22511 8041 22523 8075
rect 22465 8035 22523 8041
rect 20714 7964 20720 8016
rect 20772 8004 20778 8016
rect 20990 8004 20996 8016
rect 20772 7976 20996 8004
rect 20772 7964 20778 7976
rect 20990 7964 20996 7976
rect 21048 7964 21054 8016
rect 12768 7908 14228 7936
rect 12768 7896 12774 7908
rect 10827 7842 10916 7870
rect 11517 7871 11575 7877
rect 10827 7837 10839 7842
rect 10781 7831 10839 7837
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11790 7868 11796 7880
rect 11563 7840 11796 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 10796 7800 10824 7831
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12434 7868 12440 7880
rect 12084 7840 12440 7868
rect 12084 7809 12112 7840
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13354 7868 13360 7880
rect 13311 7840 13360 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 14090 7868 14096 7880
rect 13740 7840 14096 7868
rect 12069 7803 12127 7809
rect 6748 7772 10824 7800
rect 10888 7772 12020 7800
rect 5644 7732 5672 7760
rect 4724 7704 5672 7732
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 10689 7735 10747 7741
rect 10689 7732 10701 7735
rect 10652 7704 10701 7732
rect 10652 7692 10658 7704
rect 10689 7701 10701 7704
rect 10735 7732 10747 7735
rect 10888 7732 10916 7772
rect 10735 7704 10916 7732
rect 10735 7701 10747 7704
rect 10689 7695 10747 7701
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 11992 7732 12020 7772
rect 12069 7769 12081 7803
rect 12115 7769 12127 7803
rect 12069 7763 12127 7769
rect 12250 7760 12256 7812
rect 12308 7809 12314 7812
rect 12308 7803 12327 7809
rect 12315 7769 12327 7803
rect 13740 7800 13768 7840
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14200 7868 14228 7908
rect 15120 7908 17816 7936
rect 15120 7868 15148 7908
rect 14200 7840 15148 7868
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 16298 7868 16304 7880
rect 16255 7840 16304 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16482 7828 16488 7880
rect 16540 7828 16546 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 16632 7840 16773 7868
rect 16632 7828 16638 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17034 7868 17040 7880
rect 16991 7840 17040 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 12308 7763 12327 7769
rect 12406 7772 13768 7800
rect 12308 7760 12314 7763
rect 12406 7732 12434 7772
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14338 7803 14396 7809
rect 14338 7800 14350 7803
rect 13872 7772 14350 7800
rect 13872 7760 13878 7772
rect 14338 7769 14350 7772
rect 14384 7769 14396 7803
rect 16500 7800 16528 7828
rect 14338 7763 14396 7769
rect 15488 7772 16528 7800
rect 17144 7800 17172 7831
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17313 7871 17371 7877
rect 17313 7868 17325 7871
rect 17276 7840 17325 7868
rect 17276 7828 17282 7840
rect 17313 7837 17325 7840
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 19061 7871 19119 7877
rect 19061 7837 19073 7871
rect 19107 7868 19119 7871
rect 19150 7868 19156 7880
rect 19107 7840 19156 7868
rect 19107 7837 19119 7840
rect 19061 7831 19119 7837
rect 19150 7828 19156 7840
rect 19208 7868 19214 7880
rect 19978 7877 19984 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19208 7840 19717 7868
rect 19208 7828 19214 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19972 7868 19984 7877
rect 19939 7840 19984 7868
rect 19705 7831 19763 7837
rect 19972 7831 19984 7840
rect 17420 7800 17448 7828
rect 17144 7772 17448 7800
rect 15488 7744 15516 7772
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 18794 7803 18852 7809
rect 18794 7800 18806 7803
rect 18748 7772 18806 7800
rect 18748 7760 18754 7772
rect 18794 7769 18806 7772
rect 18840 7769 18852 7803
rect 18794 7763 18852 7769
rect 19245 7803 19303 7809
rect 19245 7769 19257 7803
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 11992 7704 12434 7732
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12860 7704 13185 7732
rect 12860 7692 12866 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 16264 7704 16497 7732
rect 16264 7692 16270 7704
rect 16485 7701 16497 7704
rect 16531 7701 16543 7735
rect 16485 7695 16543 7701
rect 17497 7735 17555 7741
rect 17497 7701 17509 7735
rect 17543 7732 17555 7735
rect 19260 7732 19288 7763
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19445 7803 19503 7809
rect 19445 7800 19457 7803
rect 19392 7772 19457 7800
rect 19392 7760 19398 7772
rect 19445 7769 19457 7772
rect 19491 7769 19503 7803
rect 19720 7800 19748 7831
rect 19978 7828 19984 7831
rect 20036 7828 20042 7880
rect 20714 7828 20720 7880
rect 20772 7828 20778 7880
rect 21192 7868 21220 8032
rect 22480 8004 22508 8035
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 22649 8075 22707 8081
rect 22649 8072 22661 8075
rect 22612 8044 22661 8072
rect 22612 8032 22618 8044
rect 22649 8041 22661 8044
rect 22695 8041 22707 8075
rect 23474 8072 23480 8084
rect 22649 8035 22707 8041
rect 22848 8044 23480 8072
rect 22848 8004 22876 8044
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 24213 8075 24271 8081
rect 24213 8072 24225 8075
rect 23624 8044 24225 8072
rect 23624 8032 23630 8044
rect 24213 8041 24225 8044
rect 24259 8072 24271 8075
rect 24394 8072 24400 8084
rect 24259 8044 24400 8072
rect 24259 8041 24271 8044
rect 24213 8035 24271 8041
rect 24394 8032 24400 8044
rect 24452 8032 24458 8084
rect 22480 7976 22876 8004
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 21508 7908 22968 7936
rect 21508 7896 21514 7908
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21192 7840 21373 7868
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21468 7840 22094 7868
rect 20732 7800 20760 7828
rect 21468 7800 21496 7840
rect 19720 7772 20760 7800
rect 20824 7772 21496 7800
rect 19445 7763 19503 7769
rect 19886 7732 19892 7744
rect 17543 7704 19892 7732
rect 17543 7701 17555 7704
rect 17497 7695 17555 7701
rect 19886 7692 19892 7704
rect 19944 7732 19950 7744
rect 20824 7732 20852 7772
rect 21542 7760 21548 7812
rect 21600 7760 21606 7812
rect 22066 7800 22094 7840
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22738 7868 22744 7880
rect 22244 7840 22744 7868
rect 22244 7828 22250 7840
rect 22738 7828 22744 7840
rect 22796 7868 22802 7880
rect 22833 7871 22891 7877
rect 22833 7868 22845 7871
rect 22796 7840 22845 7868
rect 22796 7828 22802 7840
rect 22833 7837 22845 7840
rect 22879 7837 22891 7871
rect 22940 7868 22968 7908
rect 24578 7896 24584 7948
rect 24636 7936 24642 7948
rect 25774 7936 25780 7948
rect 24636 7908 25780 7936
rect 24636 7896 24642 7908
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 25866 7896 25872 7948
rect 25924 7896 25930 7948
rect 25884 7868 25912 7896
rect 22940 7840 25912 7868
rect 22833 7831 22891 7837
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 22281 7803 22339 7809
rect 22281 7800 22293 7803
rect 22066 7772 22293 7800
rect 22281 7769 22293 7772
rect 22327 7769 22339 7803
rect 22281 7763 22339 7769
rect 23100 7803 23158 7809
rect 23100 7769 23112 7803
rect 23146 7800 23158 7803
rect 23290 7800 23296 7812
rect 23146 7772 23296 7800
rect 23146 7769 23158 7772
rect 23100 7763 23158 7769
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 24302 7760 24308 7812
rect 24360 7800 24366 7812
rect 24360 7772 28396 7800
rect 24360 7760 24366 7772
rect 28368 7744 28396 7772
rect 19944 7704 20852 7732
rect 19944 7692 19950 7704
rect 21174 7692 21180 7744
rect 21232 7692 21238 7744
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 22481 7735 22539 7741
rect 22481 7732 22493 7735
rect 21416 7704 22493 7732
rect 21416 7692 21422 7704
rect 22481 7701 22493 7704
rect 22527 7701 22539 7735
rect 22481 7695 22539 7701
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 24762 7732 24768 7744
rect 23900 7704 24768 7732
rect 23900 7692 23906 7704
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 26970 7692 26976 7744
rect 27028 7692 27034 7744
rect 28350 7692 28356 7744
rect 28408 7692 28414 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 2314 7488 2320 7540
rect 2372 7488 2378 7540
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 2866 7488 2872 7540
rect 2924 7488 2930 7540
rect 3418 7488 3424 7540
rect 3476 7488 3482 7540
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 6546 7528 6552 7540
rect 5592 7500 6552 7528
rect 5592 7488 5598 7500
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 6730 7488 6736 7540
rect 6788 7488 6794 7540
rect 10962 7528 10968 7540
rect 8128 7500 10968 7528
rect 2332 7401 2360 7488
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1688 7364 1869 7392
rect 1688 7268 1716 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 1762 7284 1768 7336
rect 1820 7284 1826 7336
rect 2056 7324 2084 7355
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 2056 7296 2421 7324
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2792 7324 2820 7488
rect 2884 7401 2912 7488
rect 4448 7460 4476 7488
rect 4448 7432 5120 7460
rect 5092 7401 5120 7432
rect 5718 7420 5724 7472
rect 5776 7420 5782 7472
rect 6632 7463 6690 7469
rect 6632 7429 6644 7463
rect 6678 7460 6690 7463
rect 6748 7460 6776 7488
rect 6678 7432 6776 7460
rect 6678 7429 6690 7432
rect 6632 7423 6690 7429
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 4545 7395 4603 7401
rect 4545 7361 4557 7395
rect 4591 7392 4603 7395
rect 5077 7395 5135 7401
rect 4591 7364 5028 7392
rect 4591 7361 4603 7364
rect 4545 7355 4603 7361
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2792 7296 2973 7324
rect 2409 7287 2467 7293
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 5000 7324 5028 7364
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5736 7324 5764 7420
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7616 7364 7941 7392
rect 7616 7352 7622 7364
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 8018 7392 8024 7404
rect 7975 7364 8024 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8128 7401 8156 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11296 7500 11345 7528
rect 11296 7488 11302 7500
rect 11333 7497 11345 7500
rect 11379 7528 11391 7531
rect 11606 7528 11612 7540
rect 11379 7500 11612 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 12710 7528 12716 7540
rect 12406 7500 12716 7528
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 12406 7460 12434 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12860 7500 12909 7528
rect 12860 7488 12866 7500
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 12897 7491 12955 7497
rect 8260 7432 12434 7460
rect 8260 7420 8266 7432
rect 12526 7420 12532 7472
rect 12584 7420 12590 7472
rect 12912 7460 12940 7491
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 13044 7500 13093 7528
rect 13044 7488 13050 7500
rect 13081 7497 13093 7500
rect 13127 7497 13139 7531
rect 14369 7531 14427 7537
rect 13081 7491 13139 7497
rect 13188 7500 13768 7528
rect 13188 7460 13216 7500
rect 12912 7432 13216 7460
rect 13249 7463 13307 7469
rect 13249 7429 13261 7463
rect 13295 7460 13307 7463
rect 13354 7460 13360 7472
rect 13295 7432 13360 7460
rect 13295 7429 13307 7432
rect 13249 7423 13307 7429
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13740 7469 13768 7500
rect 14369 7497 14381 7531
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 13449 7463 13507 7469
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 13725 7463 13783 7469
rect 13495 7432 13676 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 10226 7401 10232 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 8343 7364 8585 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 10220 7355 10232 7401
rect 10226 7352 10232 7355
rect 10284 7352 10290 7404
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10652 7364 11529 7392
rect 10652 7352 10658 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11773 7395 11831 7401
rect 11773 7392 11785 7395
rect 11664 7364 11785 7392
rect 11664 7352 11670 7364
rect 11773 7361 11785 7364
rect 11819 7361 11831 7395
rect 11773 7355 11831 7361
rect 5000 7296 5764 7324
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 1670 7216 1676 7268
rect 1728 7216 1734 7268
rect 4816 7256 4844 7284
rect 6380 7256 6408 7287
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9916 7296 9965 7324
rect 9916 7284 9922 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 12544 7324 12572 7420
rect 13648 7404 13676 7432
rect 13725 7429 13737 7463
rect 13771 7429 13783 7463
rect 14384 7460 14412 7491
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15344 7500 15853 7528
rect 15344 7488 15350 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 16298 7488 16304 7540
rect 16356 7488 16362 7540
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 16448 7500 16712 7528
rect 16448 7488 16454 7500
rect 16684 7472 16712 7500
rect 17126 7488 17132 7540
rect 17184 7488 17190 7540
rect 17218 7488 17224 7540
rect 17276 7528 17282 7540
rect 17494 7528 17500 7540
rect 17276 7500 17500 7528
rect 17276 7488 17282 7500
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18046 7488 18052 7540
rect 18104 7488 18110 7540
rect 18690 7488 18696 7540
rect 18748 7488 18754 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 19889 7531 19947 7537
rect 19889 7528 19901 7531
rect 19852 7500 19901 7528
rect 19852 7488 19858 7500
rect 19889 7497 19901 7500
rect 19935 7497 19947 7531
rect 19889 7491 19947 7497
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 22094 7488 22100 7540
rect 22152 7488 22158 7540
rect 23290 7488 23296 7540
rect 23348 7488 23354 7540
rect 24118 7488 24124 7540
rect 24176 7488 24182 7540
rect 24305 7531 24363 7537
rect 24305 7497 24317 7531
rect 24351 7528 24363 7531
rect 24854 7528 24860 7540
rect 24351 7500 24860 7528
rect 24351 7497 24363 7500
rect 24305 7491 24363 7497
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 25774 7488 25780 7540
rect 25832 7488 25838 7540
rect 26786 7488 26792 7540
rect 26844 7488 26850 7540
rect 26970 7488 26976 7540
rect 27028 7488 27034 7540
rect 28350 7488 28356 7540
rect 28408 7488 28414 7540
rect 14706 7463 14764 7469
rect 14706 7460 14718 7463
rect 13725 7423 13783 7429
rect 14108 7432 14320 7460
rect 14384 7432 14718 7460
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 13044 7364 13553 7392
rect 13044 7352 13050 7364
rect 13541 7361 13553 7364
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13630 7352 13636 7404
rect 13688 7352 13694 7404
rect 14108 7324 14136 7432
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 14292 7392 14320 7432
rect 14706 7429 14718 7432
rect 14752 7429 14764 7463
rect 14706 7423 14764 7429
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 15933 7463 15991 7469
rect 15933 7460 15945 7463
rect 15620 7432 15945 7460
rect 15620 7420 15626 7432
rect 15933 7429 15945 7432
rect 15979 7429 15991 7463
rect 15933 7423 15991 7429
rect 16149 7463 16207 7469
rect 16149 7429 16161 7463
rect 16195 7460 16207 7463
rect 16482 7460 16488 7472
rect 16195 7432 16488 7460
rect 16195 7429 16207 7432
rect 16149 7423 16207 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 16945 7463 17003 7469
rect 16945 7460 16957 7463
rect 16724 7432 16957 7460
rect 16724 7420 16730 7432
rect 16945 7429 16957 7432
rect 16991 7429 17003 7463
rect 16945 7423 17003 7429
rect 16850 7392 16856 7404
rect 14292 7364 16856 7392
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17144 7401 17172 7488
rect 17788 7432 18460 7460
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 17129 7355 17187 7361
rect 17236 7364 17509 7392
rect 12544 7296 14136 7324
rect 9953 7287 10011 7293
rect 14274 7284 14280 7336
rect 14332 7324 14338 7336
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14332 7296 14473 7324
rect 14332 7284 14338 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 16868 7324 16896 7352
rect 17236 7324 17264 7364
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 17788 7401 17816 7432
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17736 7364 17785 7392
rect 17736 7352 17742 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 16868 7296 17264 7324
rect 17313 7327 17371 7333
rect 14461 7287 14519 7293
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 18248 7324 18276 7355
rect 17359 7296 18276 7324
rect 18432 7324 18460 7432
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 19429 7463 19487 7469
rect 19429 7460 19441 7463
rect 18656 7432 19441 7460
rect 18656 7420 18662 7432
rect 19429 7429 19441 7432
rect 19475 7429 19487 7463
rect 19429 7423 19487 7429
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7392 18567 7395
rect 21192 7392 21220 7488
rect 22112 7460 22140 7488
rect 23566 7460 23572 7472
rect 22112 7432 23572 7460
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 23842 7420 23848 7472
rect 23900 7420 23906 7472
rect 18555 7364 21220 7392
rect 18555 7361 18567 7364
rect 18509 7355 18567 7361
rect 22554 7352 22560 7404
rect 22612 7352 22618 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 24136 7392 24164 7488
rect 24394 7420 24400 7472
rect 24452 7460 24458 7472
rect 24642 7463 24700 7469
rect 24642 7460 24654 7463
rect 24452 7432 24654 7460
rect 24452 7420 24458 7432
rect 24642 7429 24654 7432
rect 24688 7429 24700 7463
rect 24642 7423 24700 7429
rect 26326 7420 26332 7472
rect 26384 7420 26390 7472
rect 26988 7460 27016 7488
rect 27218 7463 27276 7469
rect 27218 7460 27230 7463
rect 26988 7432 27230 7460
rect 27218 7429 27230 7432
rect 27264 7429 27276 7463
rect 27218 7423 27276 7429
rect 24486 7392 24492 7404
rect 23523 7364 24164 7392
rect 24412 7364 24492 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 24412 7333 24440 7364
rect 24486 7352 24492 7364
rect 24544 7392 24550 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 24544 7364 26985 7392
rect 24544 7352 24550 7364
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 24397 7327 24455 7333
rect 24397 7324 24409 7327
rect 18432 7296 19334 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 4816 7228 6408 7256
rect 7300 7228 8524 7256
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6086 7188 6092 7200
rect 5868 7160 6092 7188
rect 5868 7148 5874 7160
rect 6086 7148 6092 7160
rect 6144 7188 6150 7200
rect 7300 7188 7328 7228
rect 6144 7160 7328 7188
rect 6144 7148 6150 7160
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8202 7188 8208 7200
rect 7800 7160 8208 7188
rect 7800 7148 7806 7160
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 8496 7188 8524 7228
rect 12820 7228 14044 7256
rect 12820 7188 12848 7228
rect 8496 7160 12848 7188
rect 13262 7148 13268 7200
rect 13320 7148 13326 7200
rect 13906 7148 13912 7200
rect 13964 7148 13970 7200
rect 14016 7188 14044 7228
rect 15396 7228 16160 7256
rect 15396 7188 15424 7228
rect 16132 7197 16160 7228
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 16264 7228 17448 7256
rect 16264 7216 16270 7228
rect 14016 7160 15424 7188
rect 16117 7191 16175 7197
rect 16117 7157 16129 7191
rect 16163 7157 16175 7191
rect 17420 7188 17448 7228
rect 17678 7216 17684 7268
rect 17736 7216 17742 7268
rect 17957 7259 18015 7265
rect 17957 7225 17969 7259
rect 18003 7256 18015 7259
rect 18138 7256 18144 7268
rect 18003 7228 18144 7256
rect 18003 7225 18015 7228
rect 17957 7219 18015 7225
rect 18138 7216 18144 7228
rect 18196 7256 18202 7268
rect 18196 7228 19196 7256
rect 18196 7216 18202 7228
rect 19168 7200 19196 7228
rect 18966 7188 18972 7200
rect 17420 7160 18972 7188
rect 16117 7151 16175 7157
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 19150 7148 19156 7200
rect 19208 7148 19214 7200
rect 19306 7188 19334 7296
rect 22204 7296 24409 7324
rect 19797 7259 19855 7265
rect 19797 7225 19809 7259
rect 19843 7256 19855 7259
rect 22094 7256 22100 7268
rect 19843 7228 22100 7256
rect 19843 7225 19855 7228
rect 19797 7219 19855 7225
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 22204 7200 22232 7296
rect 24397 7293 24409 7296
rect 24443 7293 24455 7327
rect 24397 7287 24455 7293
rect 24213 7259 24271 7265
rect 24213 7225 24225 7259
rect 24259 7256 24271 7259
rect 24302 7256 24308 7268
rect 24259 7228 24308 7256
rect 24259 7225 24271 7228
rect 24213 7219 24271 7225
rect 24302 7216 24308 7228
rect 24360 7216 24366 7268
rect 26602 7216 26608 7268
rect 26660 7216 26666 7268
rect 22186 7188 22192 7200
rect 19306 7160 22192 7188
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 22370 7148 22376 7200
rect 22428 7148 22434 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 7006 6984 7012 6996
rect 3844 6956 7012 6984
rect 3844 6944 3850 6956
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7742 6984 7748 6996
rect 7392 6956 7748 6984
rect 6825 6919 6883 6925
rect 1688 6888 3924 6916
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 1688 6780 1716 6888
rect 3896 6797 3924 6888
rect 6825 6885 6837 6919
rect 6871 6916 6883 6919
rect 7392 6916 7420 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 8076 6956 9720 6984
rect 8076 6944 8082 6956
rect 6871 6888 7420 6916
rect 6871 6885 6883 6888
rect 6825 6879 6883 6885
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6380 6820 6653 6848
rect 1627 6752 1716 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1688 6724 1716 6752
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 2222 6780 2228 6792
rect 1811 6752 2228 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3896 6791 3964 6797
rect 3605 6783 3663 6789
rect 3605 6780 3617 6783
rect 3200 6752 3617 6780
rect 3200 6740 3206 6752
rect 3605 6749 3617 6752
rect 3651 6749 3663 6783
rect 3896 6760 3918 6791
rect 3906 6757 3918 6760
rect 3952 6757 3964 6791
rect 6380 6789 6408 6820
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7423 6820 7512 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 3906 6751 3964 6757
rect 6365 6783 6423 6789
rect 3605 6743 3663 6749
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 1857 6715 1915 6721
rect 1857 6712 1869 6715
rect 1728 6684 1869 6712
rect 1728 6672 1734 6684
rect 1857 6681 1869 6684
rect 1903 6681 1915 6715
rect 1857 6675 1915 6681
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 7101 6715 7159 6721
rect 7101 6712 7113 6715
rect 6696 6684 7113 6712
rect 6696 6672 6702 6684
rect 7101 6681 7113 6684
rect 7147 6681 7159 6715
rect 7484 6712 7512 6820
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9272 6820 9597 6848
rect 9272 6808 9278 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9692 6848 9720 6956
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10321 6987 10379 6993
rect 10321 6984 10333 6987
rect 10284 6956 10333 6984
rect 10284 6944 10290 6956
rect 10321 6953 10333 6956
rect 10367 6953 10379 6987
rect 10321 6947 10379 6953
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 11517 6987 11575 6993
rect 10468 6956 11468 6984
rect 10468 6944 10474 6956
rect 11238 6876 11244 6928
rect 11296 6916 11302 6928
rect 11333 6919 11391 6925
rect 11333 6916 11345 6919
rect 11296 6888 11345 6916
rect 11296 6876 11302 6888
rect 11333 6885 11345 6888
rect 11379 6885 11391 6919
rect 11440 6916 11468 6956
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 11790 6984 11796 6996
rect 11563 6956 11796 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14240 6956 14473 6984
rect 14240 6944 14246 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 16942 6984 16948 6996
rect 14461 6947 14519 6953
rect 14568 6956 16948 6984
rect 14568 6916 14596 6956
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17052 6956 18092 6984
rect 11440 6888 14596 6916
rect 14645 6919 14703 6925
rect 11333 6879 11391 6885
rect 14645 6885 14657 6919
rect 14691 6885 14703 6919
rect 14645 6879 14703 6885
rect 9692 6820 10088 6848
rect 9585 6811 9643 6817
rect 7644 6783 7702 6789
rect 7644 6749 7656 6783
rect 7690 6780 7702 6783
rect 8386 6780 8392 6792
rect 7690 6752 8392 6780
rect 7690 6749 7702 6752
rect 7644 6743 7702 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8536 6752 8953 6780
rect 8536 6740 8542 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9950 6780 9956 6792
rect 9447 6752 9956 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 10060 6724 10088 6820
rect 11054 6808 11060 6860
rect 11112 6808 11118 6860
rect 14660 6848 14688 6879
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 17052 6916 17080 6956
rect 14792 6888 17080 6916
rect 18064 6916 18092 6956
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18509 6987 18567 6993
rect 18509 6984 18521 6987
rect 18288 6956 18521 6984
rect 18288 6944 18294 6956
rect 18509 6953 18521 6956
rect 18555 6953 18567 6987
rect 21450 6984 21456 6996
rect 18509 6947 18567 6953
rect 18616 6956 21456 6984
rect 18616 6916 18644 6956
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 22186 6944 22192 6996
rect 22244 6944 22250 6996
rect 22554 6944 22560 6996
rect 22612 6984 22618 6996
rect 22649 6987 22707 6993
rect 22649 6984 22661 6987
rect 22612 6956 22661 6984
rect 22612 6944 22618 6956
rect 22649 6953 22661 6956
rect 22695 6953 22707 6987
rect 22649 6947 22707 6953
rect 24394 6944 24400 6996
rect 24452 6984 24458 6996
rect 24673 6987 24731 6993
rect 24673 6984 24685 6987
rect 24452 6956 24685 6984
rect 24452 6944 24458 6956
rect 24673 6953 24685 6956
rect 24719 6953 24731 6987
rect 24673 6947 24731 6953
rect 26694 6944 26700 6996
rect 26752 6984 26758 6996
rect 27157 6987 27215 6993
rect 27157 6984 27169 6987
rect 26752 6956 27169 6984
rect 26752 6944 26758 6956
rect 27157 6953 27169 6956
rect 27203 6953 27215 6987
rect 27157 6947 27215 6953
rect 18064 6888 18644 6916
rect 20993 6919 21051 6925
rect 14792 6876 14798 6888
rect 20993 6885 21005 6919
rect 21039 6885 21051 6919
rect 20993 6879 21051 6885
rect 15470 6848 15476 6860
rect 14660 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 18138 6808 18144 6860
rect 18196 6808 18202 6860
rect 21008 6848 21036 6879
rect 22204 6848 22232 6944
rect 22833 6919 22891 6925
rect 22833 6885 22845 6919
rect 22879 6916 22891 6919
rect 23106 6916 23112 6928
rect 22879 6888 23112 6916
rect 22879 6885 22891 6888
rect 22833 6879 22891 6885
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 21008 6820 21312 6848
rect 22204 6820 23244 6848
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13906 6780 13912 6792
rect 13219 6752 13912 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 17129 6783 17187 6789
rect 14148 6752 15056 6780
rect 14148 6740 14154 6752
rect 8570 6712 8576 6724
rect 7484 6684 8576 6712
rect 7101 6675 7159 6681
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 9122 6721 9128 6724
rect 9099 6715 9128 6721
rect 9099 6681 9111 6715
rect 9099 6675 9128 6681
rect 9122 6672 9128 6675
rect 9180 6672 9186 6724
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 9861 6715 9919 6721
rect 9861 6712 9873 6715
rect 9355 6684 9873 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 9861 6681 9873 6684
rect 9907 6681 9919 6715
rect 9861 6675 9919 6681
rect 3878 6653 3884 6656
rect 3835 6647 3884 6653
rect 3835 6613 3847 6647
rect 3881 6613 3884 6647
rect 3835 6607 3884 6613
rect 3878 6604 3884 6607
rect 3936 6604 3942 6656
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9324 6644 9352 6675
rect 10042 6672 10048 6724
rect 10100 6672 10106 6724
rect 13814 6712 13820 6724
rect 13372 6684 13820 6712
rect 8803 6616 9352 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 13372 6653 13400 6684
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 14921 6715 14979 6721
rect 14921 6681 14933 6715
rect 14967 6681 14979 6715
rect 15028 6712 15056 6752
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 18156 6780 18184 6808
rect 21284 6792 21312 6820
rect 17175 6752 18184 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 20772 6752 21189 6780
rect 20772 6740 20778 6752
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 22278 6780 22284 6792
rect 21324 6752 22284 6780
rect 21324 6740 21330 6752
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 23216 6789 23244 6820
rect 23201 6783 23259 6789
rect 23201 6749 23213 6783
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 24854 6740 24860 6792
rect 24912 6740 24918 6792
rect 25774 6740 25780 6792
rect 25832 6740 25838 6792
rect 17218 6712 17224 6724
rect 15028 6684 17224 6712
rect 14921 6675 14979 6681
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6613 13415 6647
rect 13357 6607 13415 6613
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 14936 6644 14964 6675
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17396 6715 17454 6721
rect 17396 6681 17408 6715
rect 17442 6712 17454 6715
rect 18046 6712 18052 6724
rect 17442 6684 18052 6712
rect 17442 6681 17454 6684
rect 17396 6675 17454 6681
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 18690 6672 18696 6724
rect 18748 6672 18754 6724
rect 20625 6715 20683 6721
rect 20625 6681 20637 6715
rect 20671 6712 20683 6715
rect 21444 6715 21502 6721
rect 20671 6684 21404 6712
rect 20671 6681 20683 6684
rect 20625 6675 20683 6681
rect 18708 6644 18736 6672
rect 14516 6616 18736 6644
rect 14516 6604 14522 6616
rect 21082 6604 21088 6656
rect 21140 6604 21146 6656
rect 21376 6644 21404 6684
rect 21444 6681 21456 6715
rect 21490 6712 21502 6715
rect 21634 6712 21640 6724
rect 21490 6684 21640 6712
rect 21490 6681 21502 6684
rect 21444 6675 21502 6681
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 23109 6715 23167 6721
rect 23109 6712 23121 6715
rect 22066 6684 23121 6712
rect 22066 6644 22094 6684
rect 23109 6681 23121 6684
rect 23155 6712 23167 6715
rect 23750 6712 23756 6724
rect 23155 6684 23756 6712
rect 23155 6681 23167 6684
rect 23109 6675 23167 6681
rect 23750 6672 23756 6684
rect 23808 6672 23814 6724
rect 26044 6715 26102 6721
rect 26044 6681 26056 6715
rect 26090 6712 26102 6715
rect 26142 6712 26148 6724
rect 26090 6684 26148 6712
rect 26090 6681 26102 6684
rect 26044 6675 26102 6681
rect 26142 6672 26148 6684
rect 26200 6672 26206 6724
rect 21376 6616 22094 6644
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6644 22615 6647
rect 23014 6644 23020 6656
rect 22603 6616 23020 6644
rect 22603 6613 22615 6616
rect 22557 6607 22615 6613
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 23385 6647 23443 6653
rect 23385 6644 23397 6647
rect 23348 6616 23397 6644
rect 23348 6604 23354 6616
rect 23385 6613 23397 6616
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 1854 6400 1860 6452
rect 1912 6400 1918 6452
rect 2222 6400 2228 6452
rect 2280 6400 2286 6452
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 750 6264 756 6316
rect 808 6304 814 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 808 6276 1409 6304
rect 808 6264 814 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1872 6313 1900 6400
rect 2240 6313 2268 6400
rect 4632 6372 4660 6403
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 4764 6412 5304 6440
rect 4764 6400 4770 6412
rect 4954 6375 5012 6381
rect 4954 6372 4966 6375
rect 4632 6344 4966 6372
rect 4954 6341 4966 6344
rect 5000 6341 5012 6375
rect 4954 6335 5012 6341
rect 3234 6313 3240 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 3212 6307 3240 6313
rect 3212 6273 3224 6307
rect 3212 6267 3240 6273
rect 3234 6264 3240 6267
rect 3292 6264 3298 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4798 6304 4804 6316
rect 4479 6276 4804 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 5276 6304 5304 6412
rect 6086 6400 6092 6452
rect 6144 6400 6150 6452
rect 6546 6400 6552 6452
rect 6604 6400 6610 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8478 6440 8484 6452
rect 8159 6412 8484 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 6564 6372 6592 6400
rect 6978 6375 7036 6381
rect 6978 6372 6990 6375
rect 6564 6344 6990 6372
rect 6978 6341 6990 6344
rect 7024 6341 7036 6375
rect 8956 6372 8984 6403
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10502 6440 10508 6452
rect 9916 6412 10508 6440
rect 9916 6400 9922 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 13630 6440 13636 6452
rect 12492 6412 13636 6440
rect 12492 6400 12498 6412
rect 9278 6375 9336 6381
rect 9278 6372 9290 6375
rect 8956 6344 9290 6372
rect 6978 6335 7036 6341
rect 9278 6341 9290 6344
rect 9324 6341 9336 6375
rect 9278 6335 9336 6341
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 5276 6276 6745 6304
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 9692 6304 9720 6400
rect 12544 6381 12572 6412
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 16040 6412 16436 6440
rect 12529 6375 12587 6381
rect 12529 6341 12541 6375
rect 12575 6341 12587 6375
rect 12529 6335 12587 6341
rect 12710 6332 12716 6384
rect 12768 6381 12774 6384
rect 12768 6375 12792 6381
rect 12780 6341 12792 6375
rect 12768 6335 12792 6341
rect 12768 6332 12774 6335
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 14458 6372 14464 6384
rect 14056 6344 14464 6372
rect 14056 6332 14062 6344
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 16040 6381 16068 6412
rect 16025 6375 16083 6381
rect 16025 6341 16037 6375
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 16114 6332 16120 6384
rect 16172 6372 16178 6384
rect 16225 6375 16283 6381
rect 16225 6372 16237 6375
rect 16172 6344 16237 6372
rect 16172 6332 16178 6344
rect 16225 6341 16237 6344
rect 16271 6341 16283 6375
rect 16408 6372 16436 6412
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17644 6412 17785 6440
rect 17644 6400 17650 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20254 6440 20260 6452
rect 20119 6412 20260 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 21082 6400 21088 6452
rect 21140 6400 21146 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21692 6412 21833 6440
rect 21692 6400 21698 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23532 6412 23673 6440
rect 23532 6400 23538 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 24762 6440 24768 6452
rect 23661 6403 23719 6409
rect 24596 6412 24768 6440
rect 16758 6372 16764 6384
rect 16408 6344 16764 6372
rect 16225 6335 16283 6341
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 19426 6372 19432 6384
rect 17512 6344 19432 6372
rect 8803 6276 9720 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 12342 6304 12348 6316
rect 9916 6276 12348 6304
rect 9916 6264 9922 6276
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12986 6304 12992 6316
rect 12492 6276 12992 6304
rect 12492 6264 12498 6276
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 17512 6304 17540 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 20898 6332 20904 6384
rect 20956 6332 20962 6384
rect 21100 6372 21128 6400
rect 21100 6344 22048 6372
rect 13219 6302 16252 6304
rect 16408 6302 17540 6304
rect 13219 6276 17540 6302
rect 17589 6307 17647 6313
rect 13219 6273 13231 6276
rect 16224 6274 16436 6276
rect 13173 6267 13231 6273
rect 17589 6273 17601 6307
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 18690 6304 18696 6316
rect 18371 6276 18696 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4706 6236 4712 6248
rect 4304 6208 4712 6236
rect 4304 6196 4310 6208
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 8588 6236 8616 6264
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8588 6208 9045 6236
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 14274 6236 14280 6248
rect 11940 6208 14280 6236
rect 11940 6196 11946 6208
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 17126 6236 17132 6248
rect 14660 6208 17132 6236
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 3786 6168 3792 6180
rect 1627 6140 3792 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 14660 6168 14688 6208
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17494 6236 17500 6248
rect 17276 6208 17500 6236
rect 17276 6196 17282 6208
rect 17494 6196 17500 6208
rect 17552 6236 17558 6248
rect 17604 6236 17632 6267
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18800 6276 18889 6304
rect 18800 6245 18828 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6304 20867 6307
rect 20916 6304 20944 6332
rect 21085 6307 21143 6313
rect 20855 6276 21036 6304
rect 20855 6273 20867 6276
rect 20809 6267 20867 6273
rect 17552 6208 17632 6236
rect 18785 6239 18843 6245
rect 17552 6196 17558 6208
rect 18785 6205 18797 6239
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6236 20499 6239
rect 20530 6236 20536 6248
rect 20487 6208 20536 6236
rect 20487 6205 20499 6208
rect 20441 6199 20499 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 20640 6236 20668 6267
rect 20640 6208 20852 6236
rect 9968 6140 14688 6168
rect 3283 6103 3341 6109
rect 3283 6069 3295 6103
rect 3329 6100 3341 6103
rect 4062 6100 4068 6112
rect 3329 6072 4068 6100
rect 3329 6069 3341 6072
rect 3283 6063 3341 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 9968 6100 9996 6140
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 14829 6171 14887 6177
rect 14829 6168 14841 6171
rect 14792 6140 14841 6168
rect 14792 6128 14798 6140
rect 14829 6137 14841 6140
rect 14875 6168 14887 6171
rect 14875 6140 15240 6168
rect 14875 6137 14887 6140
rect 14829 6131 14887 6137
rect 6788 6072 9996 6100
rect 6788 6060 6794 6072
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 12710 6060 12716 6112
rect 12768 6060 12774 6112
rect 12894 6060 12900 6112
rect 12952 6060 12958 6112
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 14700 6072 14933 6100
rect 14700 6060 14706 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 15212 6100 15240 6140
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 16172 6140 18184 6168
rect 16172 6128 16178 6140
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15212 6072 16221 6100
rect 14921 6063 14979 6069
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 16390 6060 16396 6112
rect 16448 6060 16454 6112
rect 18156 6100 18184 6140
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 18601 6171 18659 6177
rect 18601 6168 18613 6171
rect 18288 6140 18613 6168
rect 18288 6128 18294 6140
rect 18601 6137 18613 6140
rect 18647 6137 18659 6171
rect 20824 6168 20852 6208
rect 20898 6196 20904 6248
rect 20956 6196 20962 6248
rect 21008 6236 21036 6276
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21358 6304 21364 6316
rect 21131 6276 21364 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 22020 6313 22048 6344
rect 22370 6332 22376 6384
rect 22428 6372 22434 6384
rect 22526 6375 22584 6381
rect 22526 6372 22538 6375
rect 22428 6344 22538 6372
rect 22428 6332 22434 6344
rect 22526 6341 22538 6344
rect 22572 6341 22584 6375
rect 22526 6335 22584 6341
rect 22738 6332 22744 6384
rect 22796 6332 22802 6384
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 22756 6304 22784 6332
rect 23290 6304 23296 6316
rect 22005 6267 22063 6273
rect 22296 6276 23296 6304
rect 22296 6248 22324 6276
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 21269 6239 21327 6245
rect 21269 6236 21281 6239
rect 21008 6208 21281 6236
rect 21269 6205 21281 6208
rect 21315 6205 21327 6239
rect 21269 6199 21327 6205
rect 22278 6196 22284 6248
rect 22336 6196 22342 6248
rect 22186 6168 22192 6180
rect 18601 6131 18659 6137
rect 18984 6140 20760 6168
rect 20824 6140 22192 6168
rect 18984 6100 19012 6140
rect 20732 6112 20760 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 23676 6168 23704 6403
rect 23750 6332 23756 6384
rect 23808 6372 23814 6384
rect 24596 6381 24624 6412
rect 24762 6400 24768 6412
rect 24820 6440 24826 6452
rect 25317 6443 25375 6449
rect 25317 6440 25329 6443
rect 24820 6412 25329 6440
rect 24820 6400 24826 6412
rect 25317 6409 25329 6412
rect 25363 6440 25375 6443
rect 25363 6412 25636 6440
rect 25363 6409 25375 6412
rect 25317 6403 25375 6409
rect 25608 6381 25636 6412
rect 26142 6400 26148 6452
rect 26200 6400 26206 6452
rect 24581 6375 24639 6381
rect 24581 6372 24593 6375
rect 23808 6344 24593 6372
rect 23808 6332 23814 6344
rect 24581 6341 24593 6344
rect 24627 6341 24639 6375
rect 24581 6335 24639 6341
rect 25593 6375 25651 6381
rect 25593 6341 25605 6375
rect 25639 6341 25651 6375
rect 25593 6335 25651 6341
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 24213 6239 24271 6245
rect 24213 6205 24225 6239
rect 24259 6236 24271 6239
rect 24320 6236 24348 6267
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25225 6307 25283 6313
rect 25225 6304 25237 6307
rect 24912 6276 25237 6304
rect 24912 6264 24918 6276
rect 25225 6273 25237 6276
rect 25271 6273 25283 6307
rect 26329 6307 26387 6313
rect 26329 6304 26341 6307
rect 25225 6267 25283 6273
rect 26068 6276 26341 6304
rect 26068 6245 26096 6276
rect 26329 6273 26341 6276
rect 26375 6273 26387 6307
rect 26329 6267 26387 6273
rect 24259 6208 24348 6236
rect 26053 6239 26111 6245
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 26053 6205 26065 6239
rect 26099 6205 26111 6239
rect 26053 6199 26111 6205
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 23676 6140 24041 6168
rect 24029 6137 24041 6140
rect 24075 6137 24087 6171
rect 24857 6171 24915 6177
rect 24857 6168 24869 6171
rect 24029 6131 24087 6137
rect 24412 6140 24869 6168
rect 24412 6112 24440 6140
rect 24857 6137 24869 6140
rect 24903 6137 24915 6171
rect 24857 6131 24915 6137
rect 24946 6128 24952 6180
rect 25004 6168 25010 6180
rect 25869 6171 25927 6177
rect 25869 6168 25881 6171
rect 25004 6140 25881 6168
rect 25004 6128 25010 6140
rect 25869 6137 25881 6140
rect 25915 6137 25927 6171
rect 25869 6131 25927 6137
rect 18156 6072 19012 6100
rect 19061 6103 19119 6109
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 19334 6100 19340 6112
rect 19107 6072 19340 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 20346 6060 20352 6112
rect 20404 6060 20410 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 20496 6072 20545 6100
rect 20496 6060 20502 6072
rect 20533 6069 20545 6072
rect 20579 6069 20591 6103
rect 20533 6063 20591 6069
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 23382 6100 23388 6112
rect 20772 6072 23388 6100
rect 20772 6060 20778 6072
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 24394 6060 24400 6112
rect 24452 6060 24458 6112
rect 24486 6060 24492 6112
rect 24544 6060 24550 6112
rect 25038 6060 25044 6112
rect 25096 6060 25102 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6730 5896 6736 5908
rect 5684 5868 6736 5896
rect 5684 5856 5690 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 9950 5856 9956 5908
rect 10008 5896 10014 5908
rect 10008 5868 12572 5896
rect 10008 5856 10014 5868
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 8496 5828 8524 5856
rect 9766 5828 9772 5840
rect 7883 5800 8524 5828
rect 8588 5800 9772 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 4246 5720 4252 5772
rect 4304 5720 4310 5772
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7116 5732 8125 5760
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4154 5692 4160 5704
rect 4019 5664 4160 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4264 5692 4292 5720
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 4264 5664 6101 5692
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7116 5692 7144 5732
rect 8113 5729 8125 5732
rect 8159 5760 8171 5763
rect 8588 5760 8616 5800
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 8159 5732 8616 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9876 5760 9904 5856
rect 9732 5732 9904 5760
rect 9732 5720 9738 5732
rect 6696 5664 7144 5692
rect 6696 5652 6702 5664
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 9272 5664 9597 5692
rect 9272 5652 9278 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 4494 5627 4552 5633
rect 4494 5624 4506 5627
rect 4172 5596 4506 5624
rect 4172 5565 4200 5596
rect 4494 5593 4506 5596
rect 4540 5593 4552 5627
rect 4494 5587 4552 5593
rect 6356 5627 6414 5633
rect 6356 5593 6368 5627
rect 6402 5624 6414 5627
rect 7006 5624 7012 5636
rect 6402 5596 7012 5624
rect 6402 5593 6414 5596
rect 6356 5587 6414 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 9876 5633 9904 5732
rect 10061 5701 10089 5868
rect 12544 5840 12572 5868
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 12676 5868 12725 5896
rect 12676 5856 12682 5868
rect 12713 5865 12725 5868
rect 12759 5865 12771 5899
rect 12713 5859 12771 5865
rect 13170 5856 13176 5908
rect 13228 5856 13234 5908
rect 13354 5856 13360 5908
rect 13412 5856 13418 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13722 5896 13728 5908
rect 13587 5868 13728 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 16574 5896 16580 5908
rect 14332 5868 16580 5896
rect 14332 5856 14338 5868
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10229 5831 10287 5837
rect 10229 5828 10241 5831
rect 10192 5800 10241 5828
rect 10192 5788 10198 5800
rect 10229 5797 10241 5800
rect 10275 5797 10287 5831
rect 10229 5791 10287 5797
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 12032 5800 12480 5828
rect 12032 5788 12038 5800
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 10560 5732 10609 5760
rect 10560 5720 10566 5732
rect 10597 5729 10609 5732
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5652 10382 5704
rect 11882 5692 11888 5704
rect 10428 5664 11888 5692
rect 9743 5627 9801 5633
rect 9743 5624 9755 5627
rect 9180 5596 9755 5624
rect 9180 5584 9186 5596
rect 9743 5593 9755 5596
rect 9789 5624 9801 5627
rect 9861 5627 9919 5633
rect 9789 5593 9812 5624
rect 9743 5587 9812 5593
rect 9861 5593 9873 5627
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 9953 5627 10011 5633
rect 9953 5593 9965 5627
rect 9999 5624 10011 5627
rect 10244 5624 10272 5652
rect 9999 5596 10272 5624
rect 9999 5593 10011 5596
rect 9953 5587 10011 5593
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 7466 5516 7472 5568
rect 7524 5516 7530 5568
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 9784 5556 9812 5587
rect 10428 5556 10456 5664
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12066 5652 12072 5704
rect 12124 5652 12130 5704
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 12452 5701 12480 5800
rect 12526 5788 12532 5840
rect 12584 5788 12590 5840
rect 13372 5760 13400 5856
rect 13633 5831 13691 5837
rect 13633 5797 13645 5831
rect 13679 5828 13691 5831
rect 14366 5828 14372 5840
rect 13679 5800 14372 5828
rect 13679 5797 13691 5800
rect 13633 5791 13691 5797
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 15654 5788 15660 5840
rect 15712 5828 15718 5840
rect 15749 5831 15807 5837
rect 15749 5828 15761 5831
rect 15712 5800 15761 5828
rect 15712 5788 15718 5800
rect 15749 5797 15761 5800
rect 15795 5797 15807 5831
rect 15749 5791 15807 5797
rect 13372 5732 14320 5760
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 12894 5652 12900 5704
rect 12952 5692 12958 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 12952 5664 13461 5692
rect 12952 5652 12958 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5692 13967 5695
rect 14090 5692 14096 5704
rect 13955 5664 14096 5692
rect 13955 5661 13967 5664
rect 13909 5655 13967 5661
rect 10842 5627 10900 5633
rect 10842 5624 10854 5627
rect 10520 5596 10854 5624
rect 10520 5565 10548 5596
rect 10842 5593 10854 5596
rect 10888 5593 10900 5627
rect 10842 5587 10900 5593
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 12227 5627 12285 5633
rect 12227 5624 12239 5627
rect 11756 5596 12239 5624
rect 11756 5584 11762 5596
rect 12227 5593 12239 5596
rect 12273 5624 12285 5627
rect 13924 5624 13952 5655
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14292 5701 14320 5732
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 12273 5596 13952 5624
rect 12273 5593 12285 5596
rect 12227 5587 12285 5593
rect 9784 5528 10456 5556
rect 10505 5559 10563 5565
rect 10505 5525 10517 5559
rect 10551 5525 10563 5559
rect 10505 5519 10563 5525
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 14384 5556 14412 5655
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 16114 5692 16120 5704
rect 15436 5664 16120 5692
rect 15436 5652 15442 5664
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16224 5701 16252 5868
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16942 5856 16948 5908
rect 17000 5856 17006 5908
rect 17126 5856 17132 5908
rect 17184 5896 17190 5908
rect 17221 5899 17279 5905
rect 17221 5896 17233 5899
rect 17184 5868 17233 5896
rect 17184 5856 17190 5868
rect 17221 5865 17233 5868
rect 17267 5865 17279 5899
rect 17221 5859 17279 5865
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17368 5868 17693 5896
rect 17368 5856 17374 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 17862 5856 17868 5908
rect 17920 5856 17926 5908
rect 17954 5856 17960 5908
rect 18012 5856 18018 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 18104 5868 18153 5896
rect 18104 5856 18110 5868
rect 18141 5865 18153 5868
rect 18187 5865 18199 5899
rect 18141 5859 18199 5865
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5865 18659 5899
rect 18601 5859 18659 5865
rect 16485 5831 16543 5837
rect 16485 5797 16497 5831
rect 16531 5828 16543 5831
rect 17037 5831 17095 5837
rect 17037 5828 17049 5831
rect 16531 5800 17049 5828
rect 16531 5797 16543 5800
rect 16485 5791 16543 5797
rect 17037 5797 17049 5800
rect 17083 5797 17095 5831
rect 17037 5791 17095 5797
rect 18417 5831 18475 5837
rect 18417 5797 18429 5831
rect 18463 5797 18475 5831
rect 18417 5791 18475 5797
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 18432 5760 18460 5791
rect 16623 5732 18460 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 16209 5695 16267 5701
rect 16209 5661 16221 5695
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 16666 5652 16672 5704
rect 16724 5652 16730 5704
rect 17862 5692 17868 5704
rect 17717 5664 17868 5692
rect 17717 5661 17785 5664
rect 14636 5627 14694 5633
rect 14636 5593 14648 5627
rect 14682 5624 14694 5627
rect 14734 5624 14740 5636
rect 14682 5596 14740 5624
rect 14682 5593 14694 5596
rect 14636 5587 14694 5593
rect 14734 5584 14740 5596
rect 14792 5584 14798 5636
rect 16850 5584 16856 5636
rect 16908 5624 16914 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16908 5596 17417 5624
rect 16908 5584 16914 5596
rect 17405 5593 17417 5596
rect 17451 5624 17463 5627
rect 17494 5624 17500 5636
rect 17451 5596 17500 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 17717 5630 17739 5661
rect 17727 5627 17739 5630
rect 17773 5627 17785 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18616 5692 18644 5859
rect 19150 5856 19156 5908
rect 19208 5856 19214 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 19484 5868 20300 5896
rect 19484 5856 19490 5868
rect 19168 5828 19196 5856
rect 19168 5800 19288 5828
rect 19260 5701 19288 5800
rect 20272 5760 20300 5868
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20717 5899 20775 5905
rect 20717 5896 20729 5899
rect 20404 5868 20729 5896
rect 20404 5856 20410 5868
rect 20717 5865 20729 5868
rect 20763 5865 20775 5899
rect 20717 5859 20775 5865
rect 20806 5856 20812 5908
rect 20864 5856 20870 5908
rect 20901 5899 20959 5905
rect 20901 5865 20913 5899
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 20625 5831 20683 5837
rect 20625 5797 20637 5831
rect 20671 5828 20683 5831
rect 20824 5828 20852 5856
rect 20671 5800 20852 5828
rect 20671 5797 20683 5800
rect 20625 5791 20683 5797
rect 20438 5760 20444 5772
rect 20272 5732 20444 5760
rect 20438 5720 20444 5732
rect 20496 5760 20502 5772
rect 20916 5760 20944 5859
rect 22186 5856 22192 5908
rect 22244 5896 22250 5908
rect 24394 5896 24400 5908
rect 22244 5868 24400 5896
rect 22244 5856 22250 5868
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 24486 5856 24492 5908
rect 24544 5856 24550 5908
rect 25038 5856 25044 5908
rect 25096 5896 25102 5908
rect 25096 5868 25912 5896
rect 25096 5856 25102 5868
rect 20496 5732 20944 5760
rect 20496 5720 20502 5732
rect 19245 5695 19303 5701
rect 18616 5664 19196 5692
rect 17727 5621 17785 5627
rect 18325 5627 18383 5633
rect 18325 5624 18337 5627
rect 17880 5596 18337 5624
rect 14332 5528 14412 5556
rect 14332 5516 14338 5528
rect 16298 5516 16304 5568
rect 16356 5516 16362 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 17195 5559 17253 5565
rect 17195 5556 17207 5559
rect 16540 5528 17207 5556
rect 16540 5516 16546 5528
rect 17195 5525 17207 5528
rect 17241 5525 17253 5559
rect 17512 5556 17540 5584
rect 17880 5556 17908 5596
rect 18325 5593 18337 5596
rect 18371 5624 18383 5627
rect 18785 5627 18843 5633
rect 18785 5624 18797 5627
rect 18371 5596 18797 5624
rect 18371 5593 18383 5596
rect 18325 5587 18383 5593
rect 18785 5593 18797 5596
rect 18831 5593 18843 5627
rect 19168 5624 19196 5664
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19501 5695 19559 5701
rect 19501 5692 19513 5695
rect 19392 5664 19513 5692
rect 19392 5652 19398 5664
rect 19501 5661 19513 5664
rect 19547 5661 19559 5695
rect 24504 5692 24532 5856
rect 25510 5695 25568 5701
rect 25510 5692 25522 5695
rect 19501 5655 19559 5661
rect 20364 5664 24440 5692
rect 24504 5664 25522 5692
rect 20364 5624 20392 5664
rect 19168 5596 20392 5624
rect 20640 5596 21016 5624
rect 18785 5587 18843 5593
rect 17512 5528 17908 5556
rect 18125 5559 18183 5565
rect 17195 5519 17253 5525
rect 18125 5525 18137 5559
rect 18171 5556 18183 5559
rect 18414 5556 18420 5568
rect 18171 5528 18420 5556
rect 18171 5525 18183 5528
rect 18125 5519 18183 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 18585 5559 18643 5565
rect 18585 5525 18597 5559
rect 18631 5556 18643 5559
rect 20640 5556 20668 5596
rect 18631 5528 20668 5556
rect 18631 5525 18643 5528
rect 18585 5519 18643 5525
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 20875 5559 20933 5565
rect 20875 5556 20887 5559
rect 20772 5528 20887 5556
rect 20772 5516 20778 5528
rect 20875 5525 20887 5528
rect 20921 5525 20933 5559
rect 20988 5556 21016 5596
rect 21082 5584 21088 5636
rect 21140 5584 21146 5636
rect 21358 5584 21364 5636
rect 21416 5584 21422 5636
rect 24412 5624 24440 5664
rect 25510 5661 25522 5664
rect 25556 5661 25568 5695
rect 25510 5655 25568 5661
rect 25774 5652 25780 5704
rect 25832 5652 25838 5704
rect 25884 5701 25912 5868
rect 25869 5695 25927 5701
rect 25869 5661 25881 5695
rect 25915 5661 25927 5695
rect 25869 5655 25927 5661
rect 24946 5624 24952 5636
rect 24412 5596 24952 5624
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 25792 5624 25820 5652
rect 25056 5596 25820 5624
rect 21376 5556 21404 5584
rect 25056 5568 25084 5596
rect 20988 5528 21404 5556
rect 20875 5519 20933 5525
rect 23014 5516 23020 5568
rect 23072 5556 23078 5568
rect 23750 5556 23756 5568
rect 23072 5528 23756 5556
rect 23072 5516 23078 5528
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 26050 5516 26056 5568
rect 26108 5516 26114 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 4172 5284 4200 5312
rect 5276 5284 5304 5315
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 7650 5312 7656 5364
rect 7708 5312 7714 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 4172 5256 5304 5284
rect 5721 5287 5779 5293
rect 5721 5253 5733 5287
rect 5767 5284 5779 5287
rect 6638 5284 6644 5296
rect 5767 5256 6644 5284
rect 5767 5253 5779 5256
rect 5721 5247 5779 5253
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5258 5216 5264 5228
rect 5215 5188 5264 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5258 5176 5264 5188
rect 5316 5216 5322 5228
rect 5736 5216 5764 5247
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 6822 5284 6828 5296
rect 6779 5256 6828 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 6917 5287 6975 5293
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 6963 5256 7328 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 7300 5228 7328 5256
rect 5316 5188 5764 5216
rect 7193 5219 7251 5225
rect 5316 5176 5322 5188
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 5626 5148 5632 5160
rect 5368 5120 5632 5148
rect 4893 5083 4951 5089
rect 4893 5049 4905 5083
rect 4939 5080 4951 5083
rect 5368 5080 5396 5120
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 7208 5148 7236 5179
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7668 5216 7696 5312
rect 7760 5284 7788 5315
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10376 5324 10609 5352
rect 10376 5312 10382 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 12342 5352 12348 5364
rect 10597 5315 10655 5321
rect 11624 5324 12348 5352
rect 8082 5287 8140 5293
rect 8082 5284 8094 5287
rect 7760 5256 8094 5284
rect 8082 5253 8094 5256
rect 8128 5253 8140 5287
rect 8082 5247 8140 5253
rect 10410 5244 10416 5296
rect 10468 5244 10474 5296
rect 11624 5293 11652 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 13464 5324 14320 5352
rect 11609 5287 11667 5293
rect 11609 5253 11621 5287
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 11793 5287 11851 5293
rect 11793 5253 11805 5287
rect 11839 5284 11851 5287
rect 11974 5284 11980 5296
rect 11839 5256 11980 5284
rect 11839 5253 11851 5256
rect 11793 5247 11851 5253
rect 7607 5188 7696 5216
rect 7837 5219 7895 5225
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7837 5185 7849 5219
rect 7883 5216 7895 5219
rect 8570 5216 8576 5228
rect 7883 5188 8576 5216
rect 7883 5185 7895 5188
rect 7837 5179 7895 5185
rect 6595 5120 7236 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 7852 5148 7880 5179
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10100 5188 10241 5216
rect 10100 5176 10106 5188
rect 10229 5185 10241 5188
rect 10275 5216 10287 5219
rect 11624 5216 11652 5247
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 12529 5287 12587 5293
rect 12529 5253 12541 5287
rect 12575 5284 12587 5287
rect 12618 5284 12624 5296
rect 12575 5256 12624 5284
rect 12575 5253 12587 5256
rect 12529 5247 12587 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 12745 5287 12803 5293
rect 12745 5284 12757 5287
rect 12728 5253 12757 5284
rect 12791 5284 12803 5287
rect 13464 5284 13492 5324
rect 12791 5256 13492 5284
rect 13532 5287 13590 5293
rect 12791 5253 12803 5256
rect 12728 5247 12803 5253
rect 13532 5253 13544 5287
rect 13578 5284 13590 5287
rect 14090 5284 14096 5296
rect 13578 5256 14096 5284
rect 13578 5253 13590 5256
rect 13532 5247 13590 5253
rect 10275 5188 11652 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 7708 5120 7880 5148
rect 7708 5108 7714 5120
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10870 5148 10876 5160
rect 9824 5120 10876 5148
rect 9824 5108 9830 5120
rect 10870 5108 10876 5120
rect 10928 5148 10934 5160
rect 12728 5148 12756 5247
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 14292 5284 14320 5324
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14608 5324 14657 5352
rect 14608 5312 14614 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 14645 5315 14703 5321
rect 14734 5312 14740 5364
rect 14792 5312 14798 5364
rect 15378 5312 15384 5364
rect 15436 5312 15442 5364
rect 15825 5355 15883 5361
rect 15825 5321 15837 5355
rect 15871 5352 15883 5355
rect 15930 5352 15936 5364
rect 15871 5324 15936 5352
rect 15871 5321 15883 5324
rect 15825 5315 15883 5321
rect 15930 5312 15936 5324
rect 15988 5352 15994 5364
rect 16317 5355 16375 5361
rect 16317 5352 16329 5355
rect 15988 5324 16329 5352
rect 15988 5312 15994 5324
rect 16317 5321 16329 5324
rect 16363 5321 16375 5355
rect 16317 5315 16375 5321
rect 16485 5355 16543 5361
rect 16485 5321 16497 5355
rect 16531 5352 16543 5355
rect 16666 5352 16672 5364
rect 16531 5324 16672 5352
rect 16531 5321 16543 5324
rect 16485 5315 16543 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 17678 5352 17684 5364
rect 16908 5324 17684 5352
rect 16908 5312 16914 5324
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 18506 5361 18512 5364
rect 18488 5355 18512 5361
rect 18488 5321 18500 5355
rect 18564 5352 18570 5364
rect 18564 5324 20300 5352
rect 18488 5315 18512 5321
rect 18506 5312 18512 5315
rect 18564 5312 18570 5324
rect 15396 5284 15424 5312
rect 14292 5256 15424 5284
rect 16025 5287 16083 5293
rect 16025 5253 16037 5287
rect 16071 5253 16083 5287
rect 16025 5247 16083 5253
rect 16117 5287 16175 5293
rect 16117 5253 16129 5287
rect 16163 5284 16175 5287
rect 17586 5284 17592 5296
rect 16163 5256 17592 5284
rect 16163 5253 16175 5256
rect 16117 5247 16175 5253
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 14274 5216 14280 5228
rect 13311 5188 14280 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14700 5188 14933 5216
rect 14700 5176 14706 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 16040 5216 16068 5247
rect 17586 5244 17592 5256
rect 17644 5284 17650 5296
rect 18693 5287 18751 5293
rect 18693 5284 18705 5287
rect 17644 5256 18705 5284
rect 17644 5244 17650 5256
rect 18693 5253 18705 5256
rect 18739 5253 18751 5287
rect 18693 5247 18751 5253
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5253 20223 5287
rect 20272 5284 20300 5324
rect 20530 5312 20536 5364
rect 20588 5312 20594 5364
rect 22633 5355 22691 5361
rect 22633 5321 22645 5355
rect 22679 5352 22691 5355
rect 22679 5324 23152 5352
rect 22679 5321 22691 5324
rect 22633 5315 22691 5321
rect 20381 5287 20439 5293
rect 20381 5284 20393 5287
rect 20272 5256 20393 5284
rect 20165 5247 20223 5253
rect 20381 5253 20393 5256
rect 20427 5284 20439 5287
rect 22738 5284 22744 5296
rect 20427 5256 22744 5284
rect 20427 5253 20439 5256
rect 20381 5247 20439 5253
rect 17218 5216 17224 5228
rect 16040 5188 17224 5216
rect 14921 5179 14979 5185
rect 17218 5176 17224 5188
rect 17276 5216 17282 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17276 5188 17785 5216
rect 17276 5176 17282 5188
rect 17773 5185 17785 5188
rect 17819 5216 17831 5219
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17819 5188 18061 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 10928 5120 12756 5148
rect 10928 5108 10934 5120
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14424 5120 15700 5148
rect 14424 5108 14430 5120
rect 4939 5052 5396 5080
rect 5445 5083 5503 5089
rect 4939 5049 4951 5052
rect 4893 5043 4951 5049
rect 5445 5049 5457 5083
rect 5491 5080 5503 5083
rect 5491 5052 7512 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 7484 5024 7512 5052
rect 8772 5052 12434 5080
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8772 5012 8800 5052
rect 7524 4984 8800 5012
rect 7524 4972 7530 4984
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 11974 4972 11980 5024
rect 12032 4972 12038 5024
rect 12406 5012 12434 5052
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 15672 5089 15700 5120
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17552 5120 17877 5148
rect 17552 5108 17558 5120
rect 17865 5117 17877 5120
rect 17911 5117 17923 5151
rect 20180 5148 20208 5247
rect 20254 5176 20260 5228
rect 20312 5216 20318 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20312 5188 20637 5216
rect 20312 5176 20318 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 20806 5176 20812 5228
rect 20864 5176 20870 5228
rect 20990 5176 20996 5228
rect 21048 5176 21054 5228
rect 22204 5225 22232 5256
rect 22738 5244 22744 5256
rect 22796 5244 22802 5296
rect 22833 5287 22891 5293
rect 22833 5253 22845 5287
rect 22879 5284 22891 5287
rect 23014 5284 23020 5296
rect 22879 5256 23020 5284
rect 22879 5253 22891 5256
rect 22833 5247 22891 5253
rect 22189 5219 22247 5225
rect 21836 5188 22048 5216
rect 21008 5148 21036 5176
rect 17865 5111 17923 5117
rect 17972 5120 21036 5148
rect 15657 5083 15715 5089
rect 12676 5052 12848 5080
rect 12676 5040 12682 5052
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 12406 4984 12725 5012
rect 12713 4981 12725 4984
rect 12759 4981 12771 5015
rect 12820 5012 12848 5052
rect 15657 5049 15669 5083
rect 15703 5049 15715 5083
rect 17402 5080 17408 5092
rect 15657 5043 15715 5049
rect 15764 5052 17408 5080
rect 13630 5012 13636 5024
rect 12820 4984 13636 5012
rect 12713 4975 12771 4981
rect 13630 4972 13636 4984
rect 13688 5012 13694 5024
rect 15764 5012 15792 5052
rect 17402 5040 17408 5052
rect 17460 5080 17466 5092
rect 17589 5083 17647 5089
rect 17589 5080 17601 5083
rect 17460 5052 17601 5080
rect 17460 5040 17466 5052
rect 17589 5049 17601 5052
rect 17635 5080 17647 5083
rect 17972 5080 18000 5120
rect 17635 5052 18000 5080
rect 18325 5083 18383 5089
rect 17635 5049 17647 5052
rect 17589 5043 17647 5049
rect 18325 5049 18337 5083
rect 18371 5080 18383 5083
rect 18874 5080 18880 5092
rect 18371 5052 18880 5080
rect 18371 5049 18383 5052
rect 18325 5043 18383 5049
rect 18874 5040 18880 5052
rect 18932 5040 18938 5092
rect 19150 5040 19156 5092
rect 19208 5080 19214 5092
rect 19208 5052 21128 5080
rect 19208 5040 19214 5052
rect 13688 4984 15792 5012
rect 13688 4972 13694 4984
rect 15838 4972 15844 5024
rect 15896 4972 15902 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16482 5012 16488 5024
rect 16347 4984 16488 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 17770 5012 17776 5024
rect 16632 4984 17776 5012
rect 16632 4972 16638 4984
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 19058 5012 19064 5024
rect 18555 4984 19064 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 20346 4972 20352 5024
rect 20404 4972 20410 5024
rect 20806 4972 20812 5024
rect 20864 5012 20870 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20864 4984 21005 5012
rect 20864 4972 20870 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 21100 5012 21128 5052
rect 21836 5012 21864 5188
rect 22020 5157 22048 5188
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22646 5216 22652 5228
rect 22235 5188 22269 5216
rect 22388 5188 22652 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 21913 5151 21971 5157
rect 21913 5117 21925 5151
rect 21959 5117 21971 5151
rect 21913 5111 21971 5117
rect 22005 5151 22063 5157
rect 22005 5117 22017 5151
rect 22051 5117 22063 5151
rect 22005 5111 22063 5117
rect 21928 5080 21956 5111
rect 22094 5108 22100 5160
rect 22152 5108 22158 5160
rect 22388 5157 22416 5188
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 22373 5151 22431 5157
rect 22373 5117 22385 5151
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 22738 5108 22744 5160
rect 22796 5148 22802 5160
rect 22848 5148 22876 5247
rect 23014 5244 23020 5256
rect 23072 5244 23078 5296
rect 23124 5284 23152 5324
rect 23382 5312 23388 5364
rect 23440 5312 23446 5364
rect 24121 5355 24179 5361
rect 24121 5321 24133 5355
rect 24167 5352 24179 5355
rect 24670 5352 24676 5364
rect 24167 5324 24676 5352
rect 24167 5321 24179 5324
rect 24121 5315 24179 5321
rect 23400 5284 23428 5312
rect 23124 5256 23428 5284
rect 23124 5225 23152 5256
rect 23109 5219 23167 5225
rect 23109 5185 23121 5219
rect 23155 5185 23167 5219
rect 23109 5179 23167 5185
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5216 23259 5219
rect 23474 5216 23480 5228
rect 23247 5188 23480 5216
rect 23247 5185 23259 5188
rect 23201 5179 23259 5185
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23808 5188 23857 5216
rect 23808 5176 23814 5188
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 23293 5151 23351 5157
rect 23293 5148 23305 5151
rect 22796 5120 22876 5148
rect 23124 5120 23305 5148
rect 22796 5108 22802 5120
rect 22465 5083 22523 5089
rect 22465 5080 22477 5083
rect 21928 5052 22477 5080
rect 22465 5049 22477 5052
rect 22511 5049 22523 5083
rect 22465 5043 22523 5049
rect 22572 5052 22784 5080
rect 22572 5012 22600 5052
rect 21100 4984 22600 5012
rect 20993 4975 21051 4981
rect 22646 4972 22652 5024
rect 22704 4972 22710 5024
rect 22756 5012 22784 5052
rect 22922 5040 22928 5092
rect 22980 5040 22986 5092
rect 23124 5012 23152 5120
rect 23293 5117 23305 5120
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 23382 5108 23388 5160
rect 23440 5108 23446 5160
rect 24136 5012 24164 5315
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 24946 5312 24952 5364
rect 25004 5312 25010 5364
rect 26050 5244 26056 5296
rect 26108 5293 26114 5296
rect 26108 5284 26120 5293
rect 26108 5256 26153 5284
rect 26108 5247 26120 5256
rect 26108 5244 26114 5247
rect 25774 5176 25780 5228
rect 25832 5216 25838 5228
rect 26329 5219 26387 5225
rect 26329 5216 26341 5219
rect 25832 5188 26341 5216
rect 25832 5176 25838 5188
rect 26329 5185 26341 5188
rect 26375 5185 26387 5219
rect 26329 5179 26387 5185
rect 22756 4984 24164 5012
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 4856 4780 5365 4808
rect 4856 4768 4862 4780
rect 5353 4777 5365 4780
rect 5399 4808 5411 4811
rect 7650 4808 7656 4820
rect 5399 4780 7656 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8996 4780 9321 4808
rect 8996 4768 9002 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 10042 4768 10048 4820
rect 10100 4768 10106 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 16574 4808 16580 4820
rect 13679 4780 16580 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 17494 4808 17500 4820
rect 16715 4780 17500 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 17770 4768 17776 4820
rect 17828 4768 17834 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 18690 4808 18696 4820
rect 18095 4780 18696 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 20254 4808 20260 4820
rect 18800 4780 20260 4808
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 7377 4743 7435 4749
rect 7377 4740 7389 4743
rect 7340 4712 7389 4740
rect 7340 4700 7346 4712
rect 7377 4709 7389 4712
rect 7423 4740 7435 4743
rect 10060 4740 10088 4768
rect 11698 4740 11704 4752
rect 7423 4712 10088 4740
rect 10152 4712 11704 4740
rect 7423 4709 7435 4712
rect 7377 4703 7435 4709
rect 9766 4672 9772 4684
rect 9600 4644 9772 4672
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 8478 4604 8484 4616
rect 7147 4576 8484 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9416 4576 9505 4604
rect 9416 4548 9444 4576
rect 9493 4573 9505 4576
rect 9539 4604 9551 4607
rect 9600 4604 9628 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10152 4672 10180 4712
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 12710 4700 12716 4752
rect 12768 4700 12774 4752
rect 17129 4743 17187 4749
rect 17129 4709 17141 4743
rect 17175 4709 17187 4743
rect 17788 4740 17816 4768
rect 18800 4740 18828 4780
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20496 4780 20637 4808
rect 20496 4768 20502 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 22646 4768 22652 4820
rect 22704 4768 22710 4820
rect 23014 4768 23020 4820
rect 23072 4768 23078 4820
rect 23201 4811 23259 4817
rect 23201 4777 23213 4811
rect 23247 4808 23259 4811
rect 23382 4808 23388 4820
rect 23247 4780 23388 4808
rect 23247 4777 23259 4780
rect 23201 4771 23259 4777
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 17788 4712 18828 4740
rect 17129 4703 17187 4709
rect 9876 4644 10180 4672
rect 9539 4576 9628 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 9876 4604 9904 4644
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 11204 4644 12357 4672
rect 11204 4632 11210 4644
rect 12345 4641 12357 4644
rect 12391 4672 12403 4675
rect 13998 4672 14004 4684
rect 12391 4644 14004 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 17144 4616 17172 4703
rect 20272 4672 20300 4768
rect 22097 4743 22155 4749
rect 22097 4709 22109 4743
rect 22143 4740 22155 4743
rect 22664 4740 22692 4768
rect 22143 4712 22692 4740
rect 22143 4709 22155 4712
rect 22097 4703 22155 4709
rect 22554 4672 22560 4684
rect 20272 4644 20852 4672
rect 9810 4576 9904 4604
rect 9810 4548 9838 4576
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 11054 4604 11060 4616
rect 10367 4576 11060 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 11974 4604 11980 4616
rect 11931 4576 11980 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 12084 4576 13461 4604
rect 750 4496 756 4548
rect 808 4536 814 4548
rect 1489 4539 1547 4545
rect 1489 4536 1501 4539
rect 808 4508 1501 4536
rect 808 4496 814 4508
rect 1489 4505 1501 4508
rect 1535 4505 1547 4539
rect 1489 4499 1547 4505
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 2130 4536 2136 4548
rect 1719 4508 2136 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 2130 4496 2136 4508
rect 2188 4536 2194 4548
rect 2188 4508 7236 4536
rect 2188 4496 2194 4508
rect 5626 4428 5632 4480
rect 5684 4428 5690 4480
rect 6914 4428 6920 4480
rect 6972 4428 6978 4480
rect 7208 4468 7236 4508
rect 7282 4496 7288 4548
rect 7340 4496 7346 4548
rect 7561 4539 7619 4545
rect 7561 4505 7573 4539
rect 7607 4505 7619 4539
rect 7561 4499 7619 4505
rect 7576 4468 7604 4499
rect 9398 4496 9404 4548
rect 9456 4496 9462 4548
rect 9582 4496 9588 4548
rect 9640 4496 9646 4548
rect 9766 4496 9772 4548
rect 9824 4545 9838 4548
rect 9824 4539 9853 4545
rect 9841 4505 9853 4539
rect 10781 4539 10839 4545
rect 10781 4536 10793 4539
rect 9824 4499 9853 4505
rect 9968 4508 10793 4536
rect 9824 4496 9830 4499
rect 9968 4468 9996 4508
rect 10781 4505 10793 4508
rect 10827 4536 10839 4539
rect 12084 4536 12112 4576
rect 13449 4573 13461 4576
rect 13495 4604 13507 4607
rect 13538 4604 13544 4616
rect 13495 4576 13544 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 16850 4564 16856 4616
rect 16908 4564 16914 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 17034 4604 17040 4616
rect 16991 4576 17040 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17126 4564 17132 4616
rect 17184 4564 17190 4616
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 10827 4508 12112 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 12250 4496 12256 4548
rect 12308 4536 12314 4548
rect 13906 4536 13912 4548
rect 12308 4508 13912 4536
rect 12308 4496 12314 4508
rect 13906 4496 13912 4508
rect 13964 4536 13970 4548
rect 17880 4536 17908 4567
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19245 4607 19303 4613
rect 19245 4604 19257 4607
rect 18656 4576 19257 4604
rect 18656 4564 18662 4576
rect 19245 4573 19257 4576
rect 19291 4604 19303 4607
rect 20070 4604 20076 4616
rect 19291 4576 20076 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 20070 4564 20076 4576
rect 20128 4604 20134 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20128 4576 20729 4604
rect 20128 4564 20134 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20824 4604 20852 4644
rect 22204 4644 22560 4672
rect 22204 4613 22232 4644
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 22189 4607 22247 4613
rect 22189 4604 22201 4607
rect 20824 4576 22201 4604
rect 20717 4567 20775 4573
rect 22189 4573 22201 4576
rect 22235 4573 22247 4607
rect 22189 4567 22247 4573
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 22664 4604 22692 4712
rect 22419 4576 22692 4604
rect 22756 4644 23980 4672
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 19512 4539 19570 4545
rect 13964 4508 15608 4536
rect 13964 4496 13970 4508
rect 7208 4440 9996 4468
rect 10134 4428 10140 4480
rect 10192 4428 10198 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11606 4468 11612 4480
rect 11112 4440 11612 4468
rect 11112 4428 11118 4440
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 11698 4428 11704 4480
rect 11756 4428 11762 4480
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 14090 4428 14096 4480
rect 14148 4428 14154 4480
rect 15470 4428 15476 4480
rect 15528 4428 15534 4480
rect 15580 4468 15608 4508
rect 16316 4508 19334 4536
rect 16316 4468 16344 4508
rect 15580 4440 16344 4468
rect 19306 4468 19334 4508
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 19702 4536 19708 4548
rect 19558 4508 19708 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 20990 4545 20996 4548
rect 20984 4499 20996 4545
rect 20990 4496 20996 4499
rect 21048 4496 21054 4548
rect 22557 4539 22615 4545
rect 22557 4505 22569 4539
rect 22603 4536 22615 4539
rect 22756 4536 22784 4644
rect 22940 4576 23428 4604
rect 22603 4508 22784 4536
rect 22603 4505 22615 4508
rect 22557 4499 22615 4505
rect 22830 4496 22836 4548
rect 22888 4496 22894 4548
rect 22940 4468 22968 4576
rect 23106 4545 23112 4548
rect 23049 4539 23112 4545
rect 23049 4505 23061 4539
rect 23095 4505 23112 4539
rect 23049 4499 23112 4505
rect 23106 4496 23112 4499
rect 23164 4496 23170 4548
rect 23290 4496 23296 4548
rect 23348 4496 23354 4548
rect 23400 4536 23428 4576
rect 23474 4564 23480 4616
rect 23532 4564 23538 4616
rect 23952 4613 23980 4644
rect 23937 4607 23995 4613
rect 23937 4573 23949 4607
rect 23983 4573 23995 4607
rect 23937 4567 23995 4573
rect 23400 4508 24900 4536
rect 24872 4480 24900 4508
rect 19306 4440 22968 4468
rect 23658 4428 23664 4480
rect 23716 4428 23722 4480
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 24854 4428 24860 4480
rect 24912 4428 24918 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 6822 4264 6828 4276
rect 6227 4236 6828 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 6914 4224 6920 4276
rect 6972 4224 6978 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8536 4236 9045 4264
rect 8536 4224 8542 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 5068 4131 5126 4137
rect 5068 4097 5080 4131
rect 5114 4128 5126 4131
rect 5644 4128 5672 4156
rect 6932 4137 6960 4224
rect 9048 4196 9076 4227
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 13446 4264 13452 4276
rect 9364 4236 13452 4264
rect 9364 4224 9370 4236
rect 9508 4205 9536 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 15013 4267 15071 4273
rect 15013 4233 15025 4267
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 9401 4199 9459 4205
rect 9401 4196 9413 4199
rect 9048 4168 9413 4196
rect 9401 4165 9413 4168
rect 9447 4165 9459 4199
rect 9401 4159 9459 4165
rect 9493 4199 9551 4205
rect 9493 4165 9505 4199
rect 9539 4165 9551 4199
rect 9493 4159 9551 4165
rect 9631 4199 9689 4205
rect 9631 4165 9643 4199
rect 9677 4196 9689 4199
rect 9766 4196 9772 4208
rect 9677 4168 9772 4196
rect 9677 4165 9689 4168
rect 9631 4159 9689 4165
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 10134 4196 10140 4208
rect 9916 4168 10140 4196
rect 9916 4156 9922 4168
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 11057 4199 11115 4205
rect 11057 4165 11069 4199
rect 11103 4196 11115 4199
rect 11146 4196 11152 4208
rect 11103 4168 11152 4196
rect 11103 4165 11115 4168
rect 11057 4159 11115 4165
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11701 4199 11759 4205
rect 11701 4196 11713 4199
rect 11664 4168 11713 4196
rect 11664 4156 11670 4168
rect 11701 4165 11713 4168
rect 11747 4196 11759 4199
rect 12250 4196 12256 4208
rect 11747 4168 12256 4196
rect 11747 4165 11759 4168
rect 11701 4159 11759 4165
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 12526 4196 12532 4208
rect 12360 4168 12532 4196
rect 5114 4100 5672 4128
rect 6917 4131 6975 4137
rect 5114 4097 5126 4100
rect 5068 4091 5126 4097
rect 6917 4097 6929 4131
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 7926 4137 7932 4140
rect 7920 4091 7932 4137
rect 7926 4088 7932 4091
rect 7984 4088 7990 4140
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 9088 4100 9137 4128
rect 9088 4088 9094 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 10502 4128 10508 4140
rect 9692 4100 10508 4128
rect 9692 4072 9720 4100
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4128 12219 4131
rect 12360 4128 12388 4168
rect 12526 4156 12532 4168
rect 12584 4196 12590 4208
rect 13900 4199 13958 4205
rect 12584 4168 13032 4196
rect 12584 4156 12590 4168
rect 12207 4100 12388 4128
rect 12428 4131 12486 4137
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 12428 4097 12440 4131
rect 12474 4128 12486 4131
rect 12894 4128 12900 4140
rect 12474 4100 12900 4128
rect 12474 4097 12486 4100
rect 12428 4091 12486 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13004 4128 13032 4168
rect 13900 4165 13912 4199
rect 13946 4196 13958 4199
rect 14090 4196 14096 4208
rect 13946 4168 14096 4196
rect 13946 4165 13958 4168
rect 13900 4159 13958 4165
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13004 4100 13645 4128
rect 13633 4097 13645 4100
rect 13679 4128 13691 4131
rect 15028 4128 15056 4227
rect 16482 4224 16488 4276
rect 16540 4224 16546 4276
rect 16669 4267 16727 4273
rect 16669 4233 16681 4267
rect 16715 4233 16727 4267
rect 16669 4227 16727 4233
rect 15372 4199 15430 4205
rect 15372 4165 15384 4199
rect 15418 4196 15430 4199
rect 15470 4196 15476 4208
rect 15418 4168 15476 4196
rect 15418 4165 15430 4168
rect 15372 4159 15430 4165
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 16684 4196 16712 4227
rect 19702 4224 19708 4276
rect 19760 4224 19766 4276
rect 20806 4224 20812 4276
rect 20864 4224 20870 4276
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 20990 4264 20996 4276
rect 20947 4236 20996 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 22554 4224 22560 4276
rect 22612 4264 22618 4276
rect 23290 4264 23296 4276
rect 22612 4236 23296 4264
rect 22612 4224 22618 4236
rect 23290 4224 23296 4236
rect 23348 4224 23354 4276
rect 23474 4224 23480 4276
rect 23532 4264 23538 4276
rect 23569 4267 23627 4273
rect 23569 4264 23581 4267
rect 23532 4236 23581 4264
rect 23532 4224 23538 4236
rect 23569 4233 23581 4236
rect 23615 4233 23627 4267
rect 23569 4227 23627 4233
rect 15896 4168 16712 4196
rect 15896 4156 15902 4168
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17782 4199 17840 4205
rect 17782 4196 17794 4199
rect 17184 4168 17794 4196
rect 17184 4156 17190 4168
rect 17782 4165 17794 4168
rect 17828 4165 17840 4199
rect 17782 4159 17840 4165
rect 18690 4156 18696 4208
rect 18748 4196 18754 4208
rect 19153 4199 19211 4205
rect 19153 4196 19165 4199
rect 18748 4168 19165 4196
rect 18748 4156 18754 4168
rect 19153 4165 19165 4168
rect 19199 4165 19211 4199
rect 19153 4159 19211 4165
rect 15194 4128 15200 4140
rect 13679 4100 14780 4128
rect 15028 4100 15200 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 14752 4072 14780 4100
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17552 4100 18061 4128
rect 17552 4088 17558 4100
rect 18049 4097 18061 4100
rect 18095 4128 18107 4131
rect 18598 4128 18604 4140
rect 18095 4100 18604 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19628 4100 19901 4128
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 9674 4020 9680 4072
rect 9732 4020 9738 4072
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 10060 4032 11008 4060
rect 10060 3992 10088 4032
rect 6104 3964 7696 3992
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 6104 3924 6132 3964
rect 4120 3896 6132 3924
rect 4120 3884 4126 3896
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 6604 3896 6745 3924
rect 6604 3884 6610 3896
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 7668 3924 7696 3964
rect 8956 3964 10088 3992
rect 10137 3995 10195 4001
rect 8956 3924 8984 3964
rect 10137 3961 10149 3995
rect 10183 3961 10195 3995
rect 10137 3955 10195 3961
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3961 10747 3995
rect 10980 3992 11008 4032
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 19628 4069 19656 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 20824 4128 20852 4224
rect 23750 4156 23756 4208
rect 23808 4156 23814 4208
rect 22278 4128 22284 4140
rect 20763 4100 20852 4128
rect 22204 4100 22284 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14792 4032 15117 4060
rect 14792 4020 14798 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4029 19671 4063
rect 19613 4023 19671 4029
rect 21634 4020 21640 4072
rect 21692 4060 21698 4072
rect 22204 4069 22232 4100
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22456 4131 22514 4137
rect 22456 4097 22468 4131
rect 22502 4128 22514 4131
rect 23768 4128 23796 4156
rect 22502 4100 23796 4128
rect 22502 4097 22514 4100
rect 22456 4091 22514 4097
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24774 4131 24832 4137
rect 24774 4128 24786 4131
rect 23900 4100 24786 4128
rect 23900 4088 23906 4100
rect 24774 4097 24786 4100
rect 24820 4097 24832 4131
rect 24774 4091 24832 4097
rect 22189 4063 22247 4069
rect 22189 4060 22201 4063
rect 21692 4032 22201 4060
rect 21692 4020 21698 4032
rect 22189 4029 22201 4032
rect 22235 4029 22247 4063
rect 22189 4023 22247 4029
rect 25038 4020 25044 4072
rect 25096 4020 25102 4072
rect 10980 3964 11744 3992
rect 10689 3955 10747 3961
rect 7668 3896 8984 3924
rect 6733 3887 6791 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 10152 3924 10180 3955
rect 9272 3896 10180 3924
rect 9272 3884 9278 3896
rect 10318 3884 10324 3936
rect 10376 3884 10382 3936
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 10704 3924 10732 3955
rect 10778 3924 10784 3936
rect 10704 3896 10784 3924
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 11296 3896 11621 3924
rect 11296 3884 11302 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11716 3924 11744 3964
rect 13464 3964 13676 3992
rect 13464 3924 13492 3964
rect 11716 3896 13492 3924
rect 11609 3887 11667 3893
rect 13538 3884 13544 3936
rect 13596 3884 13602 3936
rect 13648 3924 13676 3964
rect 14936 3964 15148 3992
rect 14936 3924 14964 3964
rect 13648 3896 14964 3924
rect 15120 3924 15148 3964
rect 16408 3964 16804 3992
rect 16408 3924 16436 3964
rect 15120 3896 16436 3924
rect 16776 3924 16804 3964
rect 19426 3952 19432 4004
rect 19484 3952 19490 4004
rect 19536 3964 22094 3992
rect 19536 3924 19564 3964
rect 16776 3896 19564 3924
rect 22066 3924 22094 3964
rect 23124 3964 24164 3992
rect 23124 3924 23152 3964
rect 22066 3896 23152 3924
rect 23566 3884 23572 3936
rect 23624 3924 23630 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23624 3896 23673 3924
rect 23624 3884 23630 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 24136 3924 24164 3964
rect 25866 3952 25872 4004
rect 25924 3952 25930 4004
rect 25884 3924 25912 3952
rect 24136 3896 25912 3924
rect 23661 3887 23719 3893
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 5810 3720 5816 3732
rect 5767 3692 5816 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6638 3720 6644 3732
rect 6288 3692 6644 3720
rect 5629 3655 5687 3661
rect 5629 3621 5641 3655
rect 5675 3621 5687 3655
rect 5629 3615 5687 3621
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 5644 3448 5672 3615
rect 6288 3593 6316 3692
rect 6638 3680 6644 3692
rect 6696 3720 6702 3732
rect 7650 3720 7656 3732
rect 6696 3692 7656 3720
rect 6696 3680 6702 3692
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 8113 3723 8171 3729
rect 8113 3720 8125 3723
rect 7984 3692 8125 3720
rect 7984 3680 7990 3692
rect 8113 3689 8125 3692
rect 8159 3689 8171 3723
rect 10594 3720 10600 3732
rect 8113 3683 8171 3689
rect 8312 3692 10600 3720
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6546 3525 6552 3528
rect 6540 3516 6552 3525
rect 6507 3488 6552 3516
rect 6540 3479 6552 3488
rect 6546 3476 6552 3479
rect 6604 3476 6610 3528
rect 8312 3525 8340 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11606 3720 11612 3732
rect 11379 3692 11612 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 11606 3680 11612 3692
rect 11664 3720 11670 3732
rect 12158 3720 12164 3732
rect 11664 3692 12164 3720
rect 11664 3680 11670 3692
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12526 3680 12532 3732
rect 12584 3680 12590 3732
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12768 3692 12817 3720
rect 12768 3680 12774 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 12894 3680 12900 3732
rect 12952 3680 12958 3732
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14274 3720 14280 3732
rect 14139 3692 14280 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 15712 3692 15761 3720
rect 15712 3680 15718 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 15749 3683 15807 3689
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 17092 3692 17141 3720
rect 17092 3680 17098 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 19058 3680 19064 3732
rect 19116 3680 19122 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 23566 3720 23572 3732
rect 19484 3692 23572 3720
rect 19484 3680 19490 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 23842 3680 23848 3732
rect 23900 3680 23906 3732
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3516 9919 3519
rect 9950 3516 9956 3528
rect 9907 3488 9956 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 9950 3476 9956 3488
rect 10008 3516 10014 3528
rect 11698 3525 11704 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10008 3488 11437 3516
rect 10008 3476 10014 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11692 3516 11704 3525
rect 11659 3488 11704 3516
rect 11425 3479 11483 3485
rect 11692 3479 11704 3488
rect 5644 3420 7696 3448
rect 7668 3389 7696 3420
rect 9582 3408 9588 3460
rect 9640 3408 9646 3460
rect 10226 3457 10232 3460
rect 10220 3411 10232 3457
rect 10226 3408 10232 3411
rect 10284 3408 10290 3460
rect 11440 3448 11468 3479
rect 11698 3476 11704 3479
rect 11756 3476 11762 3528
rect 12544 3448 12572 3680
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 14185 3655 14243 3661
rect 14185 3652 14197 3655
rect 13596 3624 14197 3652
rect 13596 3612 13602 3624
rect 14185 3621 14197 3624
rect 14231 3652 14243 3655
rect 15565 3655 15623 3661
rect 14231 3624 15148 3652
rect 14231 3621 14243 3624
rect 14185 3615 14243 3621
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14056 3556 14565 3584
rect 14056 3544 14062 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12860 3488 13093 3516
rect 12860 3476 12866 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 15120 3516 15148 3624
rect 15565 3621 15577 3655
rect 15611 3652 15623 3655
rect 15838 3652 15844 3664
rect 15611 3624 15844 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 16025 3655 16083 3661
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16482 3652 16488 3664
rect 16071 3624 16488 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 16945 3655 17003 3661
rect 16945 3621 16957 3655
rect 16991 3621 17003 3655
rect 19076 3652 19104 3680
rect 19521 3655 19579 3661
rect 19521 3652 19533 3655
rect 19076 3624 19533 3652
rect 16945 3615 17003 3621
rect 19521 3621 19533 3624
rect 19567 3621 19579 3655
rect 19521 3615 19579 3621
rect 16960 3584 16988 3615
rect 21266 3612 21272 3664
rect 21324 3652 21330 3664
rect 21453 3655 21511 3661
rect 21453 3652 21465 3655
rect 21324 3624 21465 3652
rect 21324 3612 21330 3624
rect 21453 3621 21465 3624
rect 21499 3621 21511 3655
rect 21453 3615 21511 3621
rect 19705 3587 19763 3593
rect 16960 3556 17816 3584
rect 17310 3516 17316 3528
rect 15120 3488 17316 3516
rect 13081 3479 13139 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17402 3476 17408 3528
rect 17460 3476 17466 3528
rect 17494 3476 17500 3528
rect 17552 3516 17558 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17552 3488 17693 3516
rect 17552 3476 17558 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17788 3516 17816 3556
rect 19705 3553 19717 3587
rect 19751 3553 19763 3587
rect 23198 3584 23204 3596
rect 19705 3547 19763 3553
rect 19904 3556 20208 3584
rect 19720 3516 19748 3547
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 17788 3488 19380 3516
rect 19720 3488 19809 3516
rect 17681 3479 17739 3485
rect 11440 3420 12020 3448
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 9600 3380 9628 3408
rect 11992 3392 12020 3420
rect 12406 3420 12572 3448
rect 15289 3451 15347 3457
rect 7699 3352 9628 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 11238 3380 11244 3392
rect 10100 3352 11244 3380
rect 10100 3340 10106 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12406 3380 12434 3420
rect 15289 3417 15301 3451
rect 15335 3448 15347 3451
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15335 3420 16313 3448
rect 15335 3417 15347 3420
rect 15289 3411 15347 3417
rect 16301 3417 16313 3420
rect 16347 3448 16359 3451
rect 16666 3448 16672 3460
rect 16347 3420 16672 3448
rect 16347 3417 16359 3420
rect 16301 3411 16359 3417
rect 12032 3352 12434 3380
rect 12032 3340 12038 3352
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 15304 3380 15332 3411
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 17926 3451 17984 3457
rect 17926 3448 17938 3451
rect 17604 3420 17938 3448
rect 13688 3352 15332 3380
rect 13688 3340 13694 3352
rect 15838 3340 15844 3392
rect 15896 3340 15902 3392
rect 17604 3389 17632 3420
rect 17926 3417 17938 3420
rect 17972 3417 17984 3451
rect 17926 3411 17984 3417
rect 19242 3408 19248 3460
rect 19300 3408 19306 3460
rect 19352 3448 19380 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 19904 3448 19932 3556
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 20180 3516 20208 3556
rect 22066 3556 23204 3584
rect 22066 3516 22094 3556
rect 23198 3544 23204 3556
rect 23256 3544 23262 3596
rect 20180 3488 22094 3516
rect 22646 3476 22652 3528
rect 22704 3476 22710 3528
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 20318 3451 20376 3457
rect 20318 3448 20330 3451
rect 19352 3420 19932 3448
rect 19996 3420 20330 3448
rect 19996 3389 20024 3420
rect 20318 3417 20330 3420
rect 20364 3417 20376 3451
rect 20318 3411 20376 3417
rect 17589 3383 17647 3389
rect 17589 3349 17601 3383
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3349 20039 3383
rect 19981 3343 20039 3349
rect 22830 3340 22836 3392
rect 22888 3340 22894 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 10226 3176 10232 3188
rect 10183 3148 10232 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 15194 3176 15200 3188
rect 10836 3148 15200 3176
rect 10836 3136 10842 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16209 3179 16267 3185
rect 16209 3145 16221 3179
rect 16255 3145 16267 3179
rect 16209 3139 16267 3145
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 9769 3111 9827 3117
rect 9769 3108 9781 3111
rect 9732 3080 9781 3108
rect 9732 3068 9738 3080
rect 9769 3077 9781 3080
rect 9815 3108 9827 3111
rect 10042 3108 10048 3120
rect 9815 3080 10048 3108
rect 9815 3077 9827 3080
rect 9769 3071 9827 3077
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3040 8723 3043
rect 9953 3043 10011 3049
rect 8711 3012 9352 3040
rect 8711 3009 8723 3012
rect 8665 3003 8723 3009
rect 9324 2981 9352 3012
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10336 3040 10364 3136
rect 16022 3108 16028 3120
rect 9999 3012 10364 3040
rect 11532 3080 16028 3108
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 11532 2972 11560 3080
rect 16022 3068 16028 3080
rect 16080 3108 16086 3120
rect 16224 3108 16252 3139
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17460 3148 17693 3176
rect 17460 3136 17466 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 22462 3136 22468 3188
rect 22520 3136 22526 3188
rect 22830 3136 22836 3188
rect 22888 3136 22894 3188
rect 16080 3080 16252 3108
rect 18141 3111 18199 3117
rect 16080 3068 16086 3080
rect 18141 3077 18153 3111
rect 18187 3108 18199 3111
rect 19242 3108 19248 3120
rect 18187 3080 19248 3108
rect 18187 3077 18199 3080
rect 18141 3071 18199 3077
rect 19242 3068 19248 3080
rect 19300 3108 19306 3120
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 19300 3080 19993 3108
rect 19300 3068 19306 3080
rect 19981 3077 19993 3080
rect 20027 3108 20039 3111
rect 22278 3108 22284 3120
rect 20027 3080 22284 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 22278 3068 22284 3080
rect 22336 3108 22342 3120
rect 22373 3111 22431 3117
rect 22373 3108 22385 3111
rect 22336 3080 22385 3108
rect 22336 3068 22342 3080
rect 22373 3077 22385 3080
rect 22419 3077 22431 3111
rect 22373 3071 22431 3077
rect 11606 3000 11612 3052
rect 11664 3000 11670 3052
rect 12250 3000 12256 3052
rect 12308 3040 12314 3052
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 12308 3012 12357 3040
rect 12308 3000 12314 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 15096 3043 15154 3049
rect 15096 3009 15108 3043
rect 15142 3040 15154 3043
rect 15378 3040 15384 3052
rect 15142 3012 15384 3040
rect 15142 3009 15154 3012
rect 15096 3003 15154 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3009 21051 3043
rect 20993 3003 21051 3009
rect 9309 2935 9367 2941
rect 9646 2944 11560 2972
rect 9493 2907 9551 2913
rect 9493 2873 9505 2907
rect 9539 2904 9551 2907
rect 9646 2904 9674 2944
rect 9539 2876 9674 2904
rect 11624 2904 11652 3000
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 12115 2944 12173 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12161 2941 12173 2944
rect 12207 2972 12219 2975
rect 12207 2944 12434 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 11624 2876 11713 2904
rect 9539 2873 9551 2876
rect 9493 2867 9551 2873
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 11701 2867 11759 2873
rect 8478 2796 8484 2848
rect 8536 2796 8542 2848
rect 11609 2839 11667 2845
rect 11609 2805 11621 2839
rect 11655 2836 11667 2839
rect 11790 2836 11796 2848
rect 11655 2808 11796 2836
rect 11655 2805 11667 2808
rect 11609 2799 11667 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12406 2836 12434 2944
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14792 2944 14841 2972
rect 14792 2932 14798 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 21008 2972 21036 3003
rect 21913 2975 21971 2981
rect 21913 2972 21925 2975
rect 21008 2944 21925 2972
rect 14829 2935 14887 2941
rect 21913 2941 21925 2944
rect 21959 2941 21971 2975
rect 21913 2935 21971 2941
rect 17865 2907 17923 2913
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 18046 2904 18052 2916
rect 17911 2876 18052 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 19702 2864 19708 2916
rect 19760 2864 19766 2916
rect 21634 2864 21640 2916
rect 21692 2864 21698 2916
rect 22097 2907 22155 2913
rect 22097 2873 22109 2907
rect 22143 2904 22155 2907
rect 22480 2904 22508 3136
rect 22848 3108 22876 3136
rect 23578 3111 23636 3117
rect 23578 3108 23590 3111
rect 22848 3080 23590 3108
rect 23578 3077 23590 3080
rect 23624 3077 23636 3111
rect 23578 3071 23636 3077
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2972 23903 2975
rect 25038 2972 25044 2984
rect 23891 2944 25044 2972
rect 23891 2941 23903 2944
rect 23845 2935 23903 2941
rect 22143 2876 22508 2904
rect 22143 2873 22155 2876
rect 22097 2867 22155 2873
rect 13446 2836 13452 2848
rect 12406 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 19518 2796 19524 2848
rect 19576 2796 19582 2848
rect 20806 2796 20812 2848
rect 20864 2796 20870 2848
rect 21652 2836 21680 2864
rect 23860 2836 23888 2935
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 21652 2808 23888 2836
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7800 2604 8125 2632
rect 7800 2592 7806 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 9232 2604 9812 2632
rect 9232 2573 9260 2604
rect 9784 2576 9812 2604
rect 11974 2592 11980 2644
rect 12032 2592 12038 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 13320 2604 13369 2632
rect 13320 2592 13326 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2533 9275 2567
rect 9674 2564 9680 2576
rect 9217 2527 9275 2533
rect 9324 2536 9680 2564
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6733 2499 6791 2505
rect 6733 2496 6745 2499
rect 6696 2468 6745 2496
rect 6696 2456 6702 2468
rect 6733 2465 6745 2468
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2496 8999 2499
rect 9324 2496 9352 2536
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 9766 2524 9772 2576
rect 9824 2524 9830 2576
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 11011 2536 11836 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 8987 2468 9352 2496
rect 9401 2499 9459 2505
rect 8987 2465 8999 2468
rect 8941 2459 8999 2465
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9416 2428 9444 2459
rect 11238 2456 11244 2508
rect 11296 2456 11302 2508
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 9416 2400 9689 2428
rect 9677 2397 9689 2400
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 11808 2428 11836 2536
rect 11992 2505 12020 2592
rect 13372 2564 13400 2595
rect 15378 2592 15384 2644
rect 15436 2592 15442 2644
rect 18046 2592 18052 2644
rect 18104 2592 18110 2644
rect 18233 2635 18291 2641
rect 18233 2601 18245 2635
rect 18279 2632 18291 2635
rect 18874 2632 18880 2644
rect 18279 2604 18880 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 19702 2592 19708 2644
rect 19760 2632 19766 2644
rect 20346 2632 20352 2644
rect 19760 2604 20352 2632
rect 19760 2592 19766 2604
rect 20346 2592 20352 2604
rect 20404 2632 20410 2644
rect 22097 2635 22155 2641
rect 22097 2632 22109 2635
rect 20404 2604 22109 2632
rect 20404 2592 20410 2604
rect 22097 2601 22109 2604
rect 22143 2601 22155 2635
rect 22097 2595 22155 2601
rect 22646 2592 22652 2644
rect 22704 2632 22710 2644
rect 22741 2635 22799 2641
rect 22741 2632 22753 2635
rect 22704 2604 22753 2632
rect 22704 2592 22710 2604
rect 22741 2601 22753 2604
rect 22787 2601 22799 2635
rect 22741 2595 22799 2601
rect 13725 2567 13783 2573
rect 13725 2564 13737 2567
rect 13372 2536 13737 2564
rect 13725 2533 13737 2536
rect 13771 2533 13783 2567
rect 18064 2564 18092 2592
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 18064 2536 19257 2564
rect 13725 2527 13783 2533
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 23014 2564 23020 2576
rect 22603 2536 23020 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 23014 2524 23020 2536
rect 23072 2524 23078 2576
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 13924 2428 13952 2459
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 11808 2400 13584 2428
rect 13924 2400 14105 2428
rect 7000 2363 7058 2369
rect 7000 2329 7012 2363
rect 7046 2360 7058 2363
rect 7190 2360 7196 2372
rect 7046 2332 7196 2360
rect 7046 2329 7058 2332
rect 7000 2323 7058 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 12222 2363 12280 2369
rect 12222 2360 12234 2363
rect 9088 2332 10824 2360
rect 9088 2320 9094 2332
rect 9490 2252 9496 2304
rect 9548 2252 9554 2304
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 10796 2301 10824 2332
rect 11900 2332 12234 2360
rect 11900 2301 11928 2332
rect 12222 2329 12234 2332
rect 12268 2329 12280 2363
rect 12222 2323 12280 2329
rect 13446 2320 13452 2372
rect 13504 2320 13510 2372
rect 13556 2360 13584 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2428 15623 2431
rect 15838 2428 15844 2440
rect 15611 2400 15844 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 17494 2428 17500 2440
rect 16899 2400 17500 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 19886 2388 19892 2440
rect 19944 2428 19950 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 19944 2400 20637 2428
rect 19944 2388 19950 2400
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20671 2400 20729 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 20973 2431 21031 2437
rect 20973 2428 20985 2431
rect 20864 2400 20985 2428
rect 20864 2388 20870 2400
rect 20973 2397 20985 2400
rect 21019 2397 21031 2431
rect 20973 2391 21031 2397
rect 13556 2332 14504 2360
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 14366 2292 14372 2304
rect 14323 2264 14372 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 14476 2292 14504 2332
rect 16482 2320 16488 2372
rect 16540 2360 16546 2372
rect 17098 2363 17156 2369
rect 17098 2360 17110 2363
rect 16540 2332 17110 2360
rect 16540 2320 16546 2332
rect 17098 2329 17110 2332
rect 17144 2329 17156 2363
rect 17098 2323 17156 2329
rect 19610 2320 19616 2372
rect 19668 2360 19674 2372
rect 20358 2363 20416 2369
rect 20358 2360 20370 2363
rect 19668 2332 20370 2360
rect 19668 2320 19674 2332
rect 20358 2329 20370 2332
rect 20404 2329 20416 2363
rect 20358 2323 20416 2329
rect 22278 2320 22284 2372
rect 22336 2320 22342 2372
rect 18690 2292 18696 2304
rect 14476 2264 18696 2292
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 7190 2048 7196 2100
rect 7248 2048 7254 2100
rect 9030 2088 9036 2100
rect 7392 2060 9036 2088
rect 6638 1912 6644 1964
rect 6696 1912 6702 1964
rect 7392 1961 7420 2060
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 9309 2091 9367 2097
rect 9309 2057 9321 2091
rect 9355 2088 9367 2091
rect 9766 2088 9772 2100
rect 9355 2060 9772 2088
rect 9355 2057 9367 2060
rect 9309 2051 9367 2057
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
rect 9861 2091 9919 2097
rect 9861 2057 9873 2091
rect 9907 2088 9919 2091
rect 10042 2088 10048 2100
rect 9907 2060 10048 2088
rect 9907 2057 9919 2060
rect 9861 2051 9919 2057
rect 10042 2048 10048 2060
rect 10100 2048 10106 2100
rect 14553 2091 14611 2097
rect 11532 2060 12434 2088
rect 8196 2023 8254 2029
rect 8196 1989 8208 2023
rect 8242 2020 8254 2023
rect 8478 2020 8484 2032
rect 8242 1992 8484 2020
rect 8242 1989 8254 1992
rect 8196 1983 8254 1989
rect 8478 1980 8484 1992
rect 8536 1980 8542 2032
rect 9401 2023 9459 2029
rect 9401 1989 9413 2023
rect 9447 2020 9459 2023
rect 9674 2020 9680 2032
rect 9447 1992 9680 2020
rect 9447 1989 9459 1992
rect 9401 1983 9459 1989
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 10226 2029 10232 2032
rect 10220 2020 10232 2029
rect 10187 1992 10232 2020
rect 10220 1983 10232 1992
rect 10226 1980 10232 1983
rect 10284 1980 10290 2032
rect 11238 1980 11244 2032
rect 11296 2020 11302 2032
rect 11532 2029 11560 2060
rect 11517 2023 11575 2029
rect 11517 2020 11529 2023
rect 11296 1992 11529 2020
rect 11296 1980 11302 1992
rect 11517 1989 11529 1992
rect 11563 1989 11575 2023
rect 12406 2020 12434 2060
rect 14553 2057 14565 2091
rect 14599 2057 14611 2091
rect 14553 2051 14611 2057
rect 12406 1992 12480 2020
rect 11517 1983 11575 1989
rect 7377 1955 7435 1961
rect 7377 1921 7389 1955
rect 7423 1921 7435 1955
rect 7377 1915 7435 1921
rect 9950 1912 9956 1964
rect 10008 1912 10014 1964
rect 11974 1912 11980 1964
rect 12032 1952 12038 1964
rect 12069 1955 12127 1961
rect 12069 1952 12081 1955
rect 12032 1924 12081 1952
rect 12032 1912 12038 1924
rect 12069 1921 12081 1924
rect 12115 1921 12127 1955
rect 12069 1915 12127 1921
rect 12158 1912 12164 1964
rect 12216 1952 12222 1964
rect 12325 1955 12383 1961
rect 12325 1952 12337 1955
rect 12216 1924 12337 1952
rect 12216 1912 12222 1924
rect 12325 1921 12337 1924
rect 12371 1921 12383 1955
rect 12452 1952 12480 1992
rect 13446 1980 13452 2032
rect 13504 2020 13510 2032
rect 14568 2020 14596 2051
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 17494 2048 17500 2100
rect 17552 2048 17558 2100
rect 18690 2048 18696 2100
rect 18748 2048 18754 2100
rect 19518 2048 19524 2100
rect 19576 2048 19582 2100
rect 19610 2048 19616 2100
rect 19668 2048 19674 2100
rect 21637 2091 21695 2097
rect 21637 2057 21649 2091
rect 21683 2057 21695 2091
rect 21637 2051 21695 2057
rect 14982 2023 15040 2029
rect 14982 2020 14994 2023
rect 13504 1992 14504 2020
rect 14568 1992 14994 2020
rect 13504 1980 13510 1992
rect 13630 1952 13636 1964
rect 12452 1924 13636 1952
rect 12325 1915 12383 1921
rect 13630 1912 13636 1924
rect 13688 1912 13694 1964
rect 14369 1955 14427 1961
rect 14369 1921 14381 1955
rect 14415 1921 14427 1955
rect 14476 1952 14504 1992
rect 14982 1989 14994 1992
rect 15028 1989 15040 2023
rect 17512 2020 17540 2048
rect 14982 1983 15040 1989
rect 15120 1992 17172 2020
rect 15120 1952 15148 1992
rect 14476 1924 15148 1952
rect 16301 1955 16359 1961
rect 14369 1915 14427 1921
rect 16301 1921 16313 1955
rect 16347 1952 16359 1955
rect 16347 1924 16574 1952
rect 16347 1921 16359 1924
rect 16301 1915 16359 1921
rect 6656 1884 6684 1912
rect 7926 1884 7932 1896
rect 6656 1856 7932 1884
rect 7926 1844 7932 1856
rect 7984 1844 7990 1896
rect 14093 1887 14151 1893
rect 14093 1853 14105 1887
rect 14139 1884 14151 1887
rect 14384 1884 14412 1915
rect 14139 1856 14412 1884
rect 14139 1853 14151 1856
rect 14093 1847 14151 1853
rect 14458 1844 14464 1896
rect 14516 1884 14522 1896
rect 14737 1887 14795 1893
rect 14737 1884 14749 1887
rect 14516 1856 14749 1884
rect 14516 1844 14522 1856
rect 14737 1853 14749 1856
rect 14783 1853 14795 1887
rect 16546 1884 16574 1924
rect 17144 1893 17172 1992
rect 17328 1992 19380 2020
rect 17328 1961 17356 1992
rect 17313 1955 17371 1961
rect 17313 1921 17325 1955
rect 17359 1921 17371 1955
rect 17313 1915 17371 1921
rect 17402 1912 17408 1964
rect 17460 1952 17466 1964
rect 17569 1955 17627 1961
rect 17569 1952 17581 1955
rect 17460 1924 17581 1952
rect 17460 1912 17466 1924
rect 17569 1921 17581 1924
rect 17615 1921 17627 1955
rect 17569 1915 17627 1921
rect 18785 1955 18843 1961
rect 18785 1921 18797 1955
rect 18831 1952 18843 1955
rect 19242 1952 19248 1964
rect 18831 1924 19248 1952
rect 18831 1921 18843 1924
rect 18785 1915 18843 1921
rect 16669 1887 16727 1893
rect 16669 1884 16681 1887
rect 16546 1856 16681 1884
rect 14737 1847 14795 1853
rect 16669 1853 16681 1856
rect 16715 1853 16727 1887
rect 16669 1847 16727 1853
rect 17129 1887 17187 1893
rect 17129 1853 17141 1887
rect 17175 1884 17187 1887
rect 17175 1856 17356 1884
rect 17175 1853 17187 1856
rect 17129 1847 17187 1853
rect 9769 1819 9827 1825
rect 9769 1785 9781 1819
rect 9815 1816 9827 1819
rect 9858 1816 9864 1828
rect 9815 1788 9864 1816
rect 9815 1785 9827 1788
rect 9769 1779 9827 1785
rect 9858 1776 9864 1788
rect 9916 1776 9922 1828
rect 11333 1819 11391 1825
rect 11333 1785 11345 1819
rect 11379 1816 11391 1819
rect 11882 1816 11888 1828
rect 11379 1788 11888 1816
rect 11379 1785 11391 1788
rect 11333 1779 11391 1785
rect 11882 1776 11888 1788
rect 11940 1776 11946 1828
rect 13909 1819 13967 1825
rect 13909 1816 13921 1819
rect 13740 1788 13921 1816
rect 13740 1760 13768 1788
rect 13909 1785 13921 1788
rect 13955 1785 13967 1819
rect 13909 1779 13967 1785
rect 16390 1776 16396 1828
rect 16448 1816 16454 1828
rect 16761 1819 16819 1825
rect 16761 1816 16773 1819
rect 16448 1788 16773 1816
rect 16448 1776 16454 1788
rect 16761 1785 16773 1788
rect 16807 1785 16819 1819
rect 16761 1779 16819 1785
rect 11974 1708 11980 1760
rect 12032 1708 12038 1760
rect 13449 1751 13507 1757
rect 13449 1717 13461 1751
rect 13495 1748 13507 1751
rect 13722 1748 13728 1760
rect 13495 1720 13728 1748
rect 13495 1717 13507 1720
rect 13449 1711 13507 1717
rect 13722 1708 13728 1720
rect 13780 1708 13786 1760
rect 16117 1751 16175 1757
rect 16117 1717 16129 1751
rect 16163 1748 16175 1751
rect 17034 1748 17040 1760
rect 16163 1720 17040 1748
rect 16163 1717 16175 1720
rect 16117 1711 16175 1717
rect 17034 1708 17040 1720
rect 17092 1708 17098 1760
rect 17328 1748 17356 1856
rect 18800 1816 18828 1915
rect 19242 1912 19248 1924
rect 19300 1912 19306 1964
rect 19352 1884 19380 1992
rect 19429 1955 19487 1961
rect 19429 1921 19441 1955
rect 19475 1952 19487 1955
rect 19536 1952 19564 2048
rect 21652 2020 21680 2051
rect 23014 2048 23020 2100
rect 23072 2088 23078 2100
rect 23201 2091 23259 2097
rect 23201 2088 23213 2091
rect 23072 2060 23213 2088
rect 23072 2048 23078 2060
rect 23201 2057 23213 2060
rect 23247 2057 23259 2091
rect 23201 2051 23259 2057
rect 22066 2023 22124 2029
rect 22066 2020 22078 2023
rect 21652 1992 22078 2020
rect 22066 1989 22078 1992
rect 22112 1989 22124 2023
rect 22066 1983 22124 1989
rect 19475 1924 19564 1952
rect 19475 1921 19487 1924
rect 19429 1915 19487 1921
rect 19610 1912 19616 1964
rect 19668 1952 19674 1964
rect 20145 1955 20203 1961
rect 20145 1952 20157 1955
rect 19668 1924 20157 1952
rect 19668 1912 19674 1924
rect 20145 1921 20157 1924
rect 20191 1921 20203 1955
rect 20145 1915 20203 1921
rect 21450 1912 21456 1964
rect 21508 1912 21514 1964
rect 21634 1912 21640 1964
rect 21692 1952 21698 1964
rect 21821 1955 21879 1961
rect 21821 1952 21833 1955
rect 21692 1924 21833 1952
rect 21692 1912 21698 1924
rect 21821 1921 21833 1924
rect 21867 1921 21879 1955
rect 21821 1915 21879 1921
rect 19886 1884 19892 1896
rect 19352 1856 19892 1884
rect 19886 1844 19892 1856
rect 19944 1844 19950 1896
rect 18248 1788 18828 1816
rect 18248 1748 18276 1788
rect 18874 1776 18880 1828
rect 18932 1816 18938 1828
rect 19061 1819 19119 1825
rect 19061 1816 19073 1819
rect 18932 1788 19073 1816
rect 18932 1776 18938 1788
rect 19061 1785 19073 1788
rect 19107 1785 19119 1819
rect 19061 1779 19119 1785
rect 17328 1720 18276 1748
rect 19242 1708 19248 1760
rect 19300 1708 19306 1760
rect 21269 1751 21327 1757
rect 21269 1717 21281 1751
rect 21315 1748 21327 1751
rect 22186 1748 22192 1760
rect 21315 1720 22192 1748
rect 21315 1717 21327 1720
rect 21269 1711 21327 1717
rect 22186 1708 22192 1720
rect 22244 1708 22250 1760
rect 1104 1658 28888 1680
rect 1104 1606 4423 1658
rect 4475 1606 4487 1658
rect 4539 1606 4551 1658
rect 4603 1606 4615 1658
rect 4667 1606 4679 1658
rect 4731 1606 11369 1658
rect 11421 1606 11433 1658
rect 11485 1606 11497 1658
rect 11549 1606 11561 1658
rect 11613 1606 11625 1658
rect 11677 1606 18315 1658
rect 18367 1606 18379 1658
rect 18431 1606 18443 1658
rect 18495 1606 18507 1658
rect 18559 1606 18571 1658
rect 18623 1606 25261 1658
rect 25313 1606 25325 1658
rect 25377 1606 25389 1658
rect 25441 1606 25453 1658
rect 25505 1606 25517 1658
rect 25569 1606 28888 1658
rect 1104 1584 28888 1606
rect 9858 1504 9864 1556
rect 9916 1544 9922 1556
rect 10321 1547 10379 1553
rect 10321 1544 10333 1547
rect 9916 1516 10333 1544
rect 9916 1504 9922 1516
rect 10321 1513 10333 1516
rect 10367 1513 10379 1547
rect 10321 1507 10379 1513
rect 12158 1504 12164 1556
rect 12216 1504 12222 1556
rect 15473 1547 15531 1553
rect 15473 1513 15485 1547
rect 15519 1544 15531 1547
rect 16390 1544 16396 1556
rect 15519 1516 16396 1544
rect 15519 1513 15531 1516
rect 15473 1507 15531 1513
rect 16390 1504 16396 1516
rect 16448 1504 16454 1556
rect 17402 1504 17408 1556
rect 17460 1504 17466 1556
rect 19150 1504 19156 1556
rect 19208 1504 19214 1556
rect 19610 1504 19616 1556
rect 19668 1504 19674 1556
rect 21450 1504 21456 1556
rect 21508 1544 21514 1556
rect 21821 1547 21879 1553
rect 21821 1544 21833 1547
rect 21508 1516 21833 1544
rect 21508 1504 21514 1516
rect 21821 1513 21833 1516
rect 21867 1513 21879 1547
rect 21821 1507 21879 1513
rect 17034 1436 17040 1488
rect 17092 1476 17098 1488
rect 19168 1476 19196 1504
rect 17092 1448 19196 1476
rect 22005 1479 22063 1485
rect 17092 1436 17098 1448
rect 22005 1445 22017 1479
rect 22051 1476 22063 1479
rect 22186 1476 22192 1488
rect 22051 1448 22192 1476
rect 22051 1445 22063 1448
rect 22005 1439 22063 1445
rect 22186 1436 22192 1448
rect 22244 1436 22250 1488
rect 7926 1368 7932 1420
rect 7984 1408 7990 1420
rect 8941 1411 8999 1417
rect 8941 1408 8953 1411
rect 7984 1380 8953 1408
rect 7984 1368 7990 1380
rect 8941 1377 8953 1380
rect 8987 1377 8999 1411
rect 8941 1371 8999 1377
rect 22278 1368 22284 1420
rect 22336 1368 22342 1420
rect 9208 1343 9266 1349
rect 9208 1309 9220 1343
rect 9254 1340 9266 1343
rect 9490 1340 9496 1352
rect 9254 1312 9496 1340
rect 9254 1309 9266 1312
rect 9208 1303 9266 1309
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 11974 1300 11980 1352
rect 12032 1300 12038 1352
rect 14366 1349 14372 1352
rect 14093 1343 14151 1349
rect 14093 1309 14105 1343
rect 14139 1309 14151 1343
rect 14360 1340 14372 1349
rect 14327 1312 14372 1340
rect 14093 1303 14151 1309
rect 14360 1303 14372 1312
rect 14108 1272 14136 1303
rect 14366 1300 14372 1303
rect 14424 1300 14430 1352
rect 14734 1300 14740 1352
rect 14792 1300 14798 1352
rect 16666 1300 16672 1352
rect 16724 1300 16730 1352
rect 17221 1343 17279 1349
rect 17221 1340 17233 1343
rect 17144 1312 17233 1340
rect 14752 1272 14780 1300
rect 14108 1244 14780 1272
rect 17144 1213 17172 1312
rect 17221 1309 17233 1312
rect 17267 1309 17279 1343
rect 17221 1303 17279 1309
rect 19242 1300 19248 1352
rect 19300 1340 19306 1352
rect 19429 1343 19487 1349
rect 19429 1340 19441 1343
rect 19300 1312 19441 1340
rect 19300 1300 19306 1312
rect 19429 1309 19441 1312
rect 19475 1309 19487 1343
rect 19429 1303 19487 1309
rect 17129 1207 17187 1213
rect 17129 1173 17141 1207
rect 17175 1173 17187 1207
rect 17129 1167 17187 1173
rect 1104 1114 29048 1136
rect 1104 1062 7896 1114
rect 7948 1062 7960 1114
rect 8012 1062 8024 1114
rect 8076 1062 8088 1114
rect 8140 1062 8152 1114
rect 8204 1062 14842 1114
rect 14894 1062 14906 1114
rect 14958 1062 14970 1114
rect 15022 1062 15034 1114
rect 15086 1062 15098 1114
rect 15150 1062 21788 1114
rect 21840 1062 21852 1114
rect 21904 1062 21916 1114
rect 21968 1062 21980 1114
rect 22032 1062 22044 1114
rect 22096 1062 28734 1114
rect 28786 1062 28798 1114
rect 28850 1062 28862 1114
rect 28914 1062 28926 1114
rect 28978 1062 28990 1114
rect 29042 1062 29048 1114
rect 1104 1040 29048 1062
<< via1 >>
rect 7896 32614 7948 32666
rect 7960 32614 8012 32666
rect 8024 32614 8076 32666
rect 8088 32614 8140 32666
rect 8152 32614 8204 32666
rect 14842 32614 14894 32666
rect 14906 32614 14958 32666
rect 14970 32614 15022 32666
rect 15034 32614 15086 32666
rect 15098 32614 15150 32666
rect 21788 32614 21840 32666
rect 21852 32614 21904 32666
rect 21916 32614 21968 32666
rect 21980 32614 22032 32666
rect 22044 32614 22096 32666
rect 28734 32614 28786 32666
rect 28798 32614 28850 32666
rect 28862 32614 28914 32666
rect 28926 32614 28978 32666
rect 28990 32614 29042 32666
rect 3976 32308 4028 32360
rect 4252 32351 4304 32360
rect 4252 32317 4261 32351
rect 4261 32317 4295 32351
rect 4295 32317 4304 32351
rect 4252 32308 4304 32317
rect 4344 32215 4396 32224
rect 4344 32181 4353 32215
rect 4353 32181 4387 32215
rect 4387 32181 4396 32215
rect 6460 32308 6512 32360
rect 7840 32308 7892 32360
rect 9588 32308 9640 32360
rect 4344 32172 4396 32181
rect 11060 32215 11112 32224
rect 11060 32181 11069 32215
rect 11069 32181 11103 32215
rect 11103 32181 11112 32215
rect 11060 32172 11112 32181
rect 4423 32070 4475 32122
rect 4487 32070 4539 32122
rect 4551 32070 4603 32122
rect 4615 32070 4667 32122
rect 4679 32070 4731 32122
rect 11369 32070 11421 32122
rect 11433 32070 11485 32122
rect 11497 32070 11549 32122
rect 11561 32070 11613 32122
rect 11625 32070 11677 32122
rect 18315 32070 18367 32122
rect 18379 32070 18431 32122
rect 18443 32070 18495 32122
rect 18507 32070 18559 32122
rect 18571 32070 18623 32122
rect 25261 32070 25313 32122
rect 25325 32070 25377 32122
rect 25389 32070 25441 32122
rect 25453 32070 25505 32122
rect 25517 32070 25569 32122
rect 11060 31968 11112 32020
rect 4252 31943 4304 31952
rect 4252 31909 4261 31943
rect 4261 31909 4295 31943
rect 4295 31909 4304 31943
rect 4252 31900 4304 31909
rect 3976 31764 4028 31816
rect 4988 31764 5040 31816
rect 6460 31875 6512 31884
rect 6460 31841 6469 31875
rect 6469 31841 6503 31875
rect 6503 31841 6512 31875
rect 6460 31832 6512 31841
rect 7840 31875 7892 31884
rect 7288 31807 7340 31816
rect 7288 31773 7297 31807
rect 7297 31773 7331 31807
rect 7331 31773 7340 31807
rect 7840 31841 7849 31875
rect 7849 31841 7883 31875
rect 7883 31841 7892 31875
rect 7840 31832 7892 31841
rect 9588 31832 9640 31884
rect 7288 31764 7340 31773
rect 8668 31764 8720 31816
rect 9312 31807 9364 31816
rect 9312 31773 9321 31807
rect 9321 31773 9355 31807
rect 9355 31773 9364 31807
rect 9312 31764 9364 31773
rect 9680 31807 9732 31816
rect 9680 31773 9689 31807
rect 9689 31773 9723 31807
rect 9723 31773 9732 31807
rect 9680 31764 9732 31773
rect 4344 31628 4396 31680
rect 9588 31628 9640 31680
rect 9680 31671 9732 31680
rect 9680 31637 9689 31671
rect 9689 31637 9723 31671
rect 9723 31637 9732 31671
rect 9680 31628 9732 31637
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 2412 31467 2464 31476
rect 2412 31433 2421 31467
rect 2421 31433 2455 31467
rect 2455 31433 2464 31467
rect 2412 31424 2464 31433
rect 2504 31288 2556 31340
rect 4344 31424 4396 31476
rect 3976 31288 4028 31340
rect 4252 31331 4304 31340
rect 4252 31297 4261 31331
rect 4261 31297 4295 31331
rect 4295 31297 4304 31331
rect 4252 31288 4304 31297
rect 4988 31288 5040 31340
rect 1860 31084 1912 31136
rect 2412 31084 2464 31136
rect 2780 31084 2832 31136
rect 3056 31152 3108 31204
rect 4804 31263 4856 31272
rect 4804 31229 4813 31263
rect 4813 31229 4847 31263
rect 4847 31229 4856 31263
rect 4804 31220 4856 31229
rect 7288 31288 7340 31340
rect 9588 31288 9640 31340
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 10324 31331 10376 31340
rect 10324 31297 10333 31331
rect 10333 31297 10367 31331
rect 10367 31297 10376 31331
rect 10324 31288 10376 31297
rect 8484 31263 8536 31272
rect 8484 31229 8493 31263
rect 8493 31229 8527 31263
rect 8527 31229 8536 31263
rect 8484 31220 8536 31229
rect 9312 31263 9364 31272
rect 9312 31229 9321 31263
rect 9321 31229 9355 31263
rect 9355 31229 9364 31263
rect 9312 31220 9364 31229
rect 8944 31084 8996 31136
rect 9404 31084 9456 31136
rect 9680 31127 9732 31136
rect 9680 31093 9689 31127
rect 9689 31093 9723 31127
rect 9723 31093 9732 31127
rect 9680 31084 9732 31093
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 10876 31127 10928 31136
rect 10876 31093 10885 31127
rect 10885 31093 10919 31127
rect 10919 31093 10928 31127
rect 10876 31084 10928 31093
rect 11244 31084 11296 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 1032 30880 1084 30932
rect 3976 30880 4028 30932
rect 4252 30880 4304 30932
rect 4988 30923 5040 30932
rect 4988 30889 4997 30923
rect 4997 30889 5031 30923
rect 5031 30889 5040 30923
rect 4988 30880 5040 30889
rect 8484 30880 8536 30932
rect 1952 30744 2004 30796
rect 2504 30744 2556 30796
rect 4804 30812 4856 30864
rect 1860 30719 1912 30728
rect 1860 30685 1869 30719
rect 1869 30685 1903 30719
rect 1903 30685 1912 30719
rect 1860 30676 1912 30685
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 2872 30608 2924 30660
rect 1860 30540 1912 30592
rect 4344 30676 4396 30728
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 5724 30676 5776 30728
rect 8668 30719 8720 30728
rect 8668 30685 8677 30719
rect 8677 30685 8711 30719
rect 8711 30685 8720 30719
rect 8668 30676 8720 30685
rect 8944 30719 8996 30728
rect 8944 30685 8953 30719
rect 8953 30685 8987 30719
rect 8987 30685 8996 30719
rect 8944 30676 8996 30685
rect 9312 30744 9364 30796
rect 9956 30812 10008 30864
rect 10416 30812 10468 30864
rect 12072 30812 12124 30864
rect 9588 30787 9640 30796
rect 9588 30753 9597 30787
rect 9597 30753 9631 30787
rect 9631 30753 9640 30787
rect 9588 30744 9640 30753
rect 9404 30676 9456 30728
rect 9864 30676 9916 30728
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 11244 30744 11296 30796
rect 10600 30676 10652 30685
rect 3056 30540 3108 30592
rect 3424 30540 3476 30592
rect 9772 30608 9824 30660
rect 10876 30608 10928 30660
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 12164 30540 12216 30592
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 3056 30336 3108 30388
rect 4804 30336 4856 30388
rect 9404 30336 9456 30388
rect 10048 30336 10100 30388
rect 10692 30336 10744 30388
rect 4068 30311 4120 30320
rect 4068 30277 4077 30311
rect 4077 30277 4111 30311
rect 4111 30277 4120 30311
rect 4068 30268 4120 30277
rect 6920 30200 6972 30252
rect 7196 30200 7248 30252
rect 9956 30243 10008 30252
rect 9956 30209 9965 30243
rect 9965 30209 9999 30243
rect 9999 30209 10008 30243
rect 9956 30200 10008 30209
rect 10600 30200 10652 30252
rect 15844 30243 15896 30252
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 1952 30175 2004 30184
rect 1952 30141 1961 30175
rect 1961 30141 1995 30175
rect 1995 30141 2004 30175
rect 1952 30132 2004 30141
rect 2964 30132 3016 30184
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 3424 30132 3476 30184
rect 3884 30132 3936 30184
rect 9864 30132 9916 30184
rect 10232 30132 10284 30184
rect 10968 30175 11020 30184
rect 10968 30141 10977 30175
rect 10977 30141 11011 30175
rect 11011 30141 11020 30175
rect 10968 30132 11020 30141
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 12164 30132 12216 30184
rect 2688 29996 2740 30048
rect 6644 30039 6696 30048
rect 6644 30005 6653 30039
rect 6653 30005 6687 30039
rect 6687 30005 6696 30039
rect 6644 29996 6696 30005
rect 15660 30039 15712 30048
rect 15660 30005 15669 30039
rect 15669 30005 15703 30039
rect 15703 30005 15712 30039
rect 15660 29996 15712 30005
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 3240 29792 3292 29844
rect 4804 29792 4856 29844
rect 1860 29699 1912 29708
rect 1860 29665 1869 29699
rect 1869 29665 1903 29699
rect 1903 29665 1912 29699
rect 1860 29656 1912 29665
rect 2136 29656 2188 29708
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 2688 29631 2740 29640
rect 2688 29597 2697 29631
rect 2697 29597 2731 29631
rect 2731 29597 2740 29631
rect 2688 29588 2740 29597
rect 4252 29588 4304 29640
rect 5080 29520 5132 29572
rect 6368 29520 6420 29572
rect 7656 29563 7708 29572
rect 7656 29529 7690 29563
rect 7690 29529 7708 29563
rect 7656 29520 7708 29529
rect 8300 29520 8352 29572
rect 1860 29452 1912 29504
rect 3056 29452 3108 29504
rect 3516 29452 3568 29504
rect 6000 29452 6052 29504
rect 7196 29452 7248 29504
rect 7564 29452 7616 29504
rect 9772 29631 9824 29640
rect 9772 29597 9781 29631
rect 9781 29597 9815 29631
rect 9815 29597 9824 29631
rect 9772 29588 9824 29597
rect 10324 29792 10376 29844
rect 12072 29792 12124 29844
rect 12164 29792 12216 29844
rect 15844 29792 15896 29844
rect 10600 29767 10652 29776
rect 10600 29733 10609 29767
rect 10609 29733 10643 29767
rect 10643 29733 10652 29767
rect 10600 29724 10652 29733
rect 11152 29724 11204 29776
rect 10968 29699 11020 29708
rect 10968 29665 10977 29699
rect 10977 29665 11011 29699
rect 11011 29665 11020 29699
rect 10968 29656 11020 29665
rect 14648 29724 14700 29776
rect 15752 29724 15804 29776
rect 9864 29520 9916 29572
rect 14464 29588 14516 29640
rect 14372 29520 14424 29572
rect 14740 29520 14792 29572
rect 10692 29452 10744 29504
rect 14096 29495 14148 29504
rect 14096 29461 14105 29495
rect 14105 29461 14139 29495
rect 14139 29461 14148 29495
rect 14096 29452 14148 29461
rect 15476 29452 15528 29504
rect 18788 29588 18840 29640
rect 16488 29520 16540 29572
rect 17960 29563 18012 29572
rect 17960 29529 17978 29563
rect 17978 29529 18012 29563
rect 17960 29520 18012 29529
rect 20812 29452 20864 29504
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 1860 29291 1912 29300
rect 1860 29257 1869 29291
rect 1869 29257 1903 29291
rect 1903 29257 1912 29291
rect 1860 29248 1912 29257
rect 3056 29248 3108 29300
rect 5080 29291 5132 29300
rect 5080 29257 5089 29291
rect 5089 29257 5123 29291
rect 5123 29257 5132 29291
rect 5080 29248 5132 29257
rect 3516 29180 3568 29232
rect 4068 29180 4120 29232
rect 2136 29112 2188 29164
rect 2964 29112 3016 29164
rect 3240 29112 3292 29164
rect 3884 29112 3936 29164
rect 5172 29155 5224 29164
rect 5172 29121 5181 29155
rect 5181 29121 5215 29155
rect 5215 29121 5224 29155
rect 5172 29112 5224 29121
rect 6920 29248 6972 29300
rect 11152 29291 11204 29300
rect 11152 29257 11161 29291
rect 11161 29257 11195 29291
rect 11195 29257 11204 29291
rect 11152 29248 11204 29257
rect 12072 29248 12124 29300
rect 14464 29248 14516 29300
rect 15660 29248 15712 29300
rect 20812 29291 20864 29300
rect 20812 29257 20821 29291
rect 20821 29257 20855 29291
rect 20855 29257 20864 29291
rect 20812 29248 20864 29257
rect 5448 29180 5500 29232
rect 9680 29112 9732 29164
rect 10324 29112 10376 29164
rect 12440 29112 12492 29164
rect 13544 29155 13596 29164
rect 13544 29121 13578 29155
rect 13578 29121 13596 29155
rect 13544 29112 13596 29121
rect 16488 29180 16540 29232
rect 15476 29112 15528 29164
rect 2780 29044 2832 29096
rect 4344 29044 4396 29096
rect 4804 29044 4856 29096
rect 1860 29019 1912 29028
rect 1860 28985 1869 29019
rect 1869 28985 1903 29019
rect 1903 28985 1912 29019
rect 1860 28976 1912 28985
rect 3056 28976 3108 29028
rect 4988 29044 5040 29096
rect 6000 29044 6052 29096
rect 7196 29087 7248 29096
rect 7196 29053 7205 29087
rect 7205 29053 7239 29087
rect 7239 29053 7248 29087
rect 7196 29044 7248 29053
rect 8392 29087 8444 29096
rect 8392 29053 8401 29087
rect 8401 29053 8435 29087
rect 8435 29053 8444 29087
rect 8392 29044 8444 29053
rect 5724 28976 5776 29028
rect 6184 28908 6236 28960
rect 7564 28908 7616 28960
rect 7748 28951 7800 28960
rect 7748 28917 7757 28951
rect 7757 28917 7791 28951
rect 7791 28917 7800 28951
rect 7748 28908 7800 28917
rect 16304 29019 16356 29028
rect 16304 28985 16313 29019
rect 16313 28985 16347 29019
rect 16347 28985 16356 29019
rect 16304 28976 16356 28985
rect 18052 29155 18104 29164
rect 18052 29121 18086 29155
rect 18086 29121 18104 29155
rect 18052 29112 18104 29121
rect 19708 29155 19760 29164
rect 19708 29121 19742 29155
rect 19742 29121 19760 29155
rect 19708 29112 19760 29121
rect 17408 29019 17460 29028
rect 17408 28985 17417 29019
rect 17417 28985 17451 29019
rect 17451 28985 17460 29019
rect 17408 28976 17460 28985
rect 8484 28908 8536 28960
rect 8852 28908 8904 28960
rect 14556 28908 14608 28960
rect 15292 28908 15344 28960
rect 16488 28908 16540 28960
rect 17132 28951 17184 28960
rect 17132 28917 17141 28951
rect 17141 28917 17175 28951
rect 17175 28917 17184 28951
rect 17132 28908 17184 28917
rect 17224 28951 17276 28960
rect 17224 28917 17233 28951
rect 17233 28917 17267 28951
rect 17267 28917 17276 28951
rect 17224 28908 17276 28917
rect 19064 28976 19116 29028
rect 18880 28908 18932 28960
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 1584 28747 1636 28756
rect 1584 28713 1593 28747
rect 1593 28713 1627 28747
rect 1627 28713 1636 28747
rect 1584 28704 1636 28713
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 2044 28543 2096 28552
rect 2044 28509 2053 28543
rect 2053 28509 2087 28543
rect 2087 28509 2096 28543
rect 2044 28500 2096 28509
rect 2780 28704 2832 28756
rect 5172 28704 5224 28756
rect 6368 28747 6420 28756
rect 6368 28713 6377 28747
rect 6377 28713 6411 28747
rect 6411 28713 6420 28747
rect 6368 28704 6420 28713
rect 7656 28704 7708 28756
rect 9680 28704 9732 28756
rect 13544 28704 13596 28756
rect 5448 28636 5500 28688
rect 2136 28407 2188 28416
rect 2136 28373 2145 28407
rect 2145 28373 2179 28407
rect 2179 28373 2188 28407
rect 2136 28364 2188 28373
rect 5540 28500 5592 28552
rect 6184 28500 6236 28552
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 6644 28500 6696 28552
rect 6920 28500 6972 28552
rect 7472 28543 7524 28552
rect 7472 28509 7481 28543
rect 7481 28509 7515 28543
rect 7515 28509 7524 28543
rect 7472 28500 7524 28509
rect 8484 28500 8536 28552
rect 8300 28432 8352 28484
rect 2964 28407 3016 28416
rect 2964 28373 2973 28407
rect 2973 28373 3007 28407
rect 3007 28373 3016 28407
rect 2964 28364 3016 28373
rect 3240 28364 3292 28416
rect 3516 28407 3568 28416
rect 3516 28373 3525 28407
rect 3525 28373 3559 28407
rect 3559 28373 3568 28407
rect 3516 28364 3568 28373
rect 3792 28364 3844 28416
rect 6276 28407 6328 28416
rect 6276 28373 6285 28407
rect 6285 28373 6319 28407
rect 6319 28373 6328 28407
rect 6276 28364 6328 28373
rect 6736 28407 6788 28416
rect 6736 28373 6745 28407
rect 6745 28373 6779 28407
rect 6779 28373 6788 28407
rect 6736 28364 6788 28373
rect 7288 28364 7340 28416
rect 8852 28500 8904 28552
rect 9036 28432 9088 28484
rect 9864 28568 9916 28620
rect 14372 28704 14424 28756
rect 14556 28679 14608 28688
rect 14556 28645 14565 28679
rect 14565 28645 14599 28679
rect 14599 28645 14608 28679
rect 14556 28636 14608 28645
rect 14740 28704 14792 28756
rect 17132 28704 17184 28756
rect 18052 28704 18104 28756
rect 9772 28543 9824 28552
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 10324 28543 10376 28552
rect 10324 28509 10333 28543
rect 10333 28509 10367 28543
rect 10367 28509 10376 28543
rect 10324 28500 10376 28509
rect 10600 28543 10652 28552
rect 10600 28509 10609 28543
rect 10609 28509 10643 28543
rect 10643 28509 10652 28543
rect 10600 28500 10652 28509
rect 14096 28500 14148 28552
rect 17960 28636 18012 28688
rect 15292 28500 15344 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 17224 28500 17276 28552
rect 18144 28500 18196 28552
rect 18880 28500 18932 28552
rect 21456 28543 21508 28552
rect 21456 28509 21465 28543
rect 21465 28509 21499 28543
rect 21499 28509 21508 28543
rect 21456 28500 21508 28509
rect 9312 28364 9364 28416
rect 11704 28407 11756 28416
rect 11704 28373 11713 28407
rect 11713 28373 11747 28407
rect 11747 28373 11756 28407
rect 11704 28364 11756 28373
rect 15200 28407 15252 28416
rect 15200 28373 15209 28407
rect 15209 28373 15243 28407
rect 15243 28373 15252 28407
rect 15200 28364 15252 28373
rect 18052 28407 18104 28416
rect 18052 28373 18061 28407
rect 18061 28373 18095 28407
rect 18095 28373 18104 28407
rect 18052 28364 18104 28373
rect 19156 28432 19208 28484
rect 25872 28432 25924 28484
rect 20628 28407 20680 28416
rect 20628 28373 20637 28407
rect 20637 28373 20671 28407
rect 20671 28373 20680 28407
rect 20628 28364 20680 28373
rect 21640 28407 21692 28416
rect 21640 28373 21649 28407
rect 21649 28373 21683 28407
rect 21683 28373 21692 28407
rect 21640 28364 21692 28373
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 1768 28203 1820 28212
rect 1768 28169 1801 28203
rect 1801 28169 1820 28203
rect 1768 28160 1820 28169
rect 2136 28160 2188 28212
rect 2596 28092 2648 28144
rect 2044 28067 2096 28076
rect 2044 28033 2053 28067
rect 2053 28033 2087 28067
rect 2087 28033 2096 28067
rect 2044 28024 2096 28033
rect 2504 28024 2556 28076
rect 3516 28160 3568 28212
rect 5632 28160 5684 28212
rect 6276 28160 6328 28212
rect 6736 28160 6788 28212
rect 7748 28160 7800 28212
rect 9036 28160 9088 28212
rect 6920 28092 6972 28144
rect 3516 28067 3568 28076
rect 3516 28033 3524 28067
rect 3524 28033 3568 28067
rect 3516 28024 3568 28033
rect 4252 28024 4304 28076
rect 4804 28024 4856 28076
rect 3148 27956 3200 28008
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 5264 27888 5316 27940
rect 8392 28092 8444 28144
rect 9312 28160 9364 28212
rect 10600 28160 10652 28212
rect 15200 28160 15252 28212
rect 18052 28160 18104 28212
rect 19156 28203 19208 28212
rect 19156 28169 19165 28203
rect 19165 28169 19199 28203
rect 19199 28169 19208 28203
rect 19156 28160 19208 28169
rect 19708 28203 19760 28212
rect 19708 28169 19717 28203
rect 19717 28169 19751 28203
rect 19751 28169 19760 28203
rect 19708 28160 19760 28169
rect 21640 28160 21692 28212
rect 9772 28092 9824 28144
rect 20720 28092 20772 28144
rect 9864 28067 9916 28076
rect 9864 28033 9873 28067
rect 9873 28033 9907 28067
rect 9907 28033 9916 28067
rect 9864 28024 9916 28033
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 12808 28067 12860 28076
rect 12808 28033 12817 28067
rect 12817 28033 12851 28067
rect 12851 28033 12860 28067
rect 12808 28024 12860 28033
rect 2780 27820 2832 27872
rect 3056 27820 3108 27872
rect 3332 27820 3384 27872
rect 5080 27820 5132 27872
rect 5540 27863 5592 27872
rect 5540 27829 5549 27863
rect 5549 27829 5583 27863
rect 5583 27829 5592 27863
rect 5540 27820 5592 27829
rect 5908 27863 5960 27872
rect 5908 27829 5917 27863
rect 5917 27829 5951 27863
rect 5951 27829 5960 27863
rect 5908 27820 5960 27829
rect 6552 27820 6604 27872
rect 6736 27820 6788 27872
rect 7196 27863 7248 27872
rect 7196 27829 7205 27863
rect 7205 27829 7239 27863
rect 7239 27829 7248 27863
rect 7196 27820 7248 27829
rect 8484 27820 8536 27872
rect 9312 27820 9364 27872
rect 12624 27863 12676 27872
rect 12624 27829 12633 27863
rect 12633 27829 12667 27863
rect 12667 27829 12676 27863
rect 12624 27820 12676 27829
rect 13912 27863 13964 27872
rect 13912 27829 13921 27863
rect 13921 27829 13955 27863
rect 13955 27829 13964 27863
rect 13912 27820 13964 27829
rect 15660 28024 15712 28076
rect 18972 28067 19024 28076
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 19892 28067 19944 28076
rect 19892 28033 19901 28067
rect 19901 28033 19935 28067
rect 19935 28033 19944 28067
rect 19892 28024 19944 28033
rect 14648 27999 14700 28008
rect 14648 27965 14657 27999
rect 14657 27965 14691 27999
rect 14691 27965 14700 27999
rect 14648 27956 14700 27965
rect 18880 27999 18932 28008
rect 18880 27965 18889 27999
rect 18889 27965 18923 27999
rect 18923 27965 18932 27999
rect 18880 27956 18932 27965
rect 21640 27956 21692 28008
rect 15568 27820 15620 27872
rect 17500 27863 17552 27872
rect 17500 27829 17509 27863
rect 17509 27829 17543 27863
rect 17543 27829 17552 27863
rect 17500 27820 17552 27829
rect 21180 27820 21232 27872
rect 22192 27820 22244 27872
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 4252 27616 4304 27668
rect 2872 27591 2924 27600
rect 2872 27557 2881 27591
rect 2881 27557 2915 27591
rect 2915 27557 2924 27591
rect 2872 27548 2924 27557
rect 4804 27548 4856 27600
rect 7564 27616 7616 27668
rect 9864 27616 9916 27668
rect 10416 27616 10468 27668
rect 1676 27480 1728 27532
rect 3332 27523 3384 27532
rect 3332 27489 3341 27523
rect 3341 27489 3375 27523
rect 3375 27489 3384 27523
rect 3332 27480 3384 27489
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 2228 27412 2280 27421
rect 2504 27412 2556 27464
rect 3148 27412 3200 27464
rect 4988 27480 5040 27532
rect 5356 27480 5408 27532
rect 4804 27412 4856 27464
rect 5172 27412 5224 27464
rect 5448 27412 5500 27464
rect 8944 27548 8996 27600
rect 6920 27455 6972 27464
rect 6920 27421 6929 27455
rect 6929 27421 6963 27455
rect 6963 27421 6972 27455
rect 10324 27480 10376 27532
rect 15200 27548 15252 27600
rect 15292 27548 15344 27600
rect 18144 27659 18196 27668
rect 18144 27625 18153 27659
rect 18153 27625 18187 27659
rect 18187 27625 18196 27659
rect 18144 27616 18196 27625
rect 18972 27616 19024 27668
rect 19892 27616 19944 27668
rect 20720 27659 20772 27668
rect 20720 27625 20729 27659
rect 20729 27625 20763 27659
rect 20763 27625 20772 27659
rect 20720 27616 20772 27625
rect 21456 27659 21508 27668
rect 21456 27625 21465 27659
rect 21465 27625 21499 27659
rect 21499 27625 21508 27659
rect 21456 27616 21508 27625
rect 22192 27616 22244 27668
rect 17408 27548 17460 27600
rect 20628 27548 20680 27600
rect 6920 27412 6972 27421
rect 9312 27455 9364 27464
rect 9312 27421 9321 27455
rect 9321 27421 9355 27455
rect 9355 27421 9364 27455
rect 9312 27412 9364 27421
rect 10692 27455 10744 27464
rect 10692 27421 10701 27455
rect 10701 27421 10735 27455
rect 10735 27421 10744 27455
rect 10692 27412 10744 27421
rect 12440 27412 12492 27464
rect 12624 27455 12676 27464
rect 12624 27421 12658 27455
rect 12658 27421 12676 27455
rect 12624 27412 12676 27421
rect 2044 27276 2096 27328
rect 2136 27319 2188 27328
rect 2136 27285 2145 27319
rect 2145 27285 2179 27319
rect 2179 27285 2188 27319
rect 2136 27276 2188 27285
rect 4160 27319 4212 27328
rect 4160 27285 4169 27319
rect 4169 27285 4203 27319
rect 4203 27285 4212 27319
rect 4160 27276 4212 27285
rect 4252 27319 4304 27328
rect 4252 27285 4261 27319
rect 4261 27285 4295 27319
rect 4295 27285 4304 27319
rect 4252 27276 4304 27285
rect 5908 27344 5960 27396
rect 6736 27344 6788 27396
rect 7196 27387 7248 27396
rect 7196 27353 7230 27387
rect 7230 27353 7248 27387
rect 7196 27344 7248 27353
rect 13636 27344 13688 27396
rect 4896 27276 4948 27328
rect 5540 27276 5592 27328
rect 8484 27276 8536 27328
rect 9128 27276 9180 27328
rect 11704 27276 11756 27328
rect 13176 27276 13228 27328
rect 14556 27412 14608 27464
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 14924 27455 14976 27464
rect 14924 27421 14933 27455
rect 14933 27421 14967 27455
rect 14967 27421 14976 27455
rect 14924 27412 14976 27421
rect 15016 27455 15068 27464
rect 15016 27421 15025 27455
rect 15025 27421 15059 27455
rect 15059 27421 15068 27455
rect 15016 27412 15068 27421
rect 15200 27412 15252 27464
rect 15292 27412 15344 27464
rect 15568 27455 15620 27464
rect 15568 27421 15575 27455
rect 15575 27421 15620 27455
rect 15568 27412 15620 27421
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 16120 27455 16172 27464
rect 16120 27421 16129 27455
rect 16129 27421 16163 27455
rect 16163 27421 16172 27455
rect 16120 27412 16172 27421
rect 21548 27480 21600 27532
rect 19616 27455 19668 27464
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 16580 27344 16632 27396
rect 16856 27344 16908 27396
rect 17684 27387 17736 27396
rect 17684 27353 17693 27387
rect 17693 27353 17727 27387
rect 17727 27353 17736 27387
rect 17684 27344 17736 27353
rect 15292 27319 15344 27328
rect 15292 27285 15301 27319
rect 15301 27285 15335 27319
rect 15335 27285 15344 27319
rect 15292 27276 15344 27285
rect 15568 27276 15620 27328
rect 16028 27319 16080 27328
rect 16028 27285 16037 27319
rect 16037 27285 16071 27319
rect 16071 27285 16080 27319
rect 16028 27276 16080 27285
rect 16120 27276 16172 27328
rect 16488 27276 16540 27328
rect 19432 27344 19484 27396
rect 19800 27387 19852 27396
rect 19800 27353 19809 27387
rect 19809 27353 19843 27387
rect 19843 27353 19852 27387
rect 19800 27344 19852 27353
rect 20444 27387 20496 27396
rect 20444 27353 20453 27387
rect 20453 27353 20487 27387
rect 20487 27353 20496 27387
rect 20444 27344 20496 27353
rect 20536 27344 20588 27396
rect 21180 27344 21232 27396
rect 24400 27412 24452 27464
rect 20812 27276 20864 27328
rect 22928 27276 22980 27328
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 1676 27072 1728 27124
rect 2136 27072 2188 27124
rect 5172 27115 5224 27124
rect 5172 27081 5181 27115
rect 5181 27081 5215 27115
rect 5215 27081 5224 27115
rect 5172 27072 5224 27081
rect 2504 27004 2556 27056
rect 2044 26936 2096 26988
rect 2228 26911 2280 26920
rect 2228 26877 2237 26911
rect 2237 26877 2271 26911
rect 2271 26877 2280 26911
rect 2228 26868 2280 26877
rect 3056 26979 3108 26988
rect 3056 26945 3065 26979
rect 3065 26945 3099 26979
rect 3099 26945 3108 26979
rect 3056 26936 3108 26945
rect 3332 26979 3384 26988
rect 3332 26945 3341 26979
rect 3341 26945 3375 26979
rect 3375 26945 3384 26979
rect 3332 26936 3384 26945
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 4160 27047 4212 27056
rect 4160 27013 4169 27047
rect 4169 27013 4203 27047
rect 4203 27013 4212 27047
rect 6828 27072 6880 27124
rect 7104 27072 7156 27124
rect 10692 27115 10744 27124
rect 10692 27081 10701 27115
rect 10701 27081 10735 27115
rect 10735 27081 10744 27115
rect 10692 27072 10744 27081
rect 4160 27004 4212 27013
rect 2872 26800 2924 26852
rect 2964 26800 3016 26852
rect 3608 26800 3660 26852
rect 5264 26868 5316 26920
rect 5540 27047 5592 27056
rect 5540 27013 5549 27047
rect 5549 27013 5583 27047
rect 5583 27013 5592 27047
rect 5540 27004 5592 27013
rect 6092 27004 6144 27056
rect 8944 27004 8996 27056
rect 6276 26868 6328 26920
rect 7380 26936 7432 26988
rect 8484 26936 8536 26988
rect 6000 26800 6052 26852
rect 6092 26800 6144 26852
rect 8300 26868 8352 26920
rect 9128 26868 9180 26920
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 12440 27004 12492 27056
rect 13912 27072 13964 27124
rect 14740 27072 14792 27124
rect 15292 27072 15344 27124
rect 15384 27115 15436 27124
rect 15384 27081 15393 27115
rect 15393 27081 15427 27115
rect 15427 27081 15436 27115
rect 15384 27072 15436 27081
rect 11980 26979 12032 26988
rect 11980 26945 12014 26979
rect 12014 26945 12032 26979
rect 9404 26868 9456 26920
rect 11980 26936 12032 26945
rect 3700 26732 3752 26784
rect 5080 26732 5132 26784
rect 6368 26732 6420 26784
rect 7012 26775 7064 26784
rect 7012 26741 7021 26775
rect 7021 26741 7055 26775
rect 7055 26741 7064 26775
rect 7012 26732 7064 26741
rect 7656 26732 7708 26784
rect 9220 26732 9272 26784
rect 9496 26732 9548 26784
rect 12900 26868 12952 26920
rect 11060 26732 11112 26784
rect 13084 26775 13136 26784
rect 13084 26741 13093 26775
rect 13093 26741 13127 26775
rect 13127 26741 13136 26775
rect 15660 26936 15712 26988
rect 16488 26936 16540 26988
rect 17500 27072 17552 27124
rect 21548 27072 21600 27124
rect 17408 27004 17460 27056
rect 19616 27004 19668 27056
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 19156 26979 19208 26988
rect 19156 26945 19165 26979
rect 19165 26945 19199 26979
rect 19199 26945 19208 26979
rect 19156 26936 19208 26945
rect 19708 26979 19760 26988
rect 19708 26945 19742 26979
rect 19742 26945 19760 26979
rect 19708 26936 19760 26945
rect 18052 26868 18104 26920
rect 18880 26868 18932 26920
rect 23940 26936 23992 26988
rect 24400 26936 24452 26988
rect 23296 26868 23348 26920
rect 22928 26843 22980 26852
rect 22928 26809 22937 26843
rect 22937 26809 22971 26843
rect 22971 26809 22980 26843
rect 22928 26800 22980 26809
rect 13084 26732 13136 26741
rect 14832 26732 14884 26784
rect 16120 26732 16172 26784
rect 17040 26732 17092 26784
rect 18972 26775 19024 26784
rect 18972 26741 18981 26775
rect 18981 26741 19015 26775
rect 19015 26741 19024 26775
rect 18972 26732 19024 26741
rect 20076 26732 20128 26784
rect 20444 26732 20496 26784
rect 23020 26775 23072 26784
rect 23020 26741 23029 26775
rect 23029 26741 23063 26775
rect 23063 26741 23072 26775
rect 23020 26732 23072 26741
rect 23112 26775 23164 26784
rect 23112 26741 23121 26775
rect 23121 26741 23155 26775
rect 23155 26741 23164 26775
rect 23112 26732 23164 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 2872 26528 2924 26580
rect 3332 26528 3384 26580
rect 4988 26528 5040 26580
rect 5540 26528 5592 26580
rect 6000 26528 6052 26580
rect 6092 26528 6144 26580
rect 6736 26528 6788 26580
rect 7012 26528 7064 26580
rect 9956 26571 10008 26580
rect 9956 26537 9965 26571
rect 9965 26537 9999 26571
rect 9999 26537 10008 26571
rect 9956 26528 10008 26537
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 12808 26528 12860 26580
rect 13084 26528 13136 26580
rect 16580 26571 16632 26580
rect 16580 26537 16589 26571
rect 16589 26537 16623 26571
rect 16623 26537 16632 26571
rect 16580 26528 16632 26537
rect 17316 26528 17368 26580
rect 4344 26460 4396 26512
rect 2688 26392 2740 26444
rect 2964 26324 3016 26376
rect 3516 26324 3568 26376
rect 4528 26367 4580 26376
rect 4528 26333 4537 26367
rect 4537 26333 4571 26367
rect 4571 26333 4580 26367
rect 4528 26324 4580 26333
rect 4804 26324 4856 26376
rect 3424 26299 3476 26308
rect 3424 26265 3433 26299
rect 3433 26265 3467 26299
rect 3467 26265 3476 26299
rect 3424 26256 3476 26265
rect 5080 26392 5132 26444
rect 6276 26392 6328 26444
rect 5908 26367 5960 26376
rect 5908 26333 5917 26367
rect 5917 26333 5951 26367
rect 5951 26333 5960 26367
rect 5908 26324 5960 26333
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 6368 26367 6420 26376
rect 6368 26333 6377 26367
rect 6377 26333 6411 26367
rect 6411 26333 6420 26367
rect 6368 26324 6420 26333
rect 6552 26324 6604 26376
rect 13176 26503 13228 26512
rect 13176 26469 13185 26503
rect 13185 26469 13219 26503
rect 13219 26469 13228 26503
rect 13176 26460 13228 26469
rect 13636 26460 13688 26512
rect 16764 26460 16816 26512
rect 19708 26571 19760 26580
rect 19708 26537 19717 26571
rect 19717 26537 19751 26571
rect 19751 26537 19760 26571
rect 19708 26528 19760 26537
rect 23020 26528 23072 26580
rect 23940 26528 23992 26580
rect 11060 26392 11112 26444
rect 14464 26392 14516 26444
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12164 26324 12216 26333
rect 15752 26367 15804 26376
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 17132 26324 17184 26376
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 18972 26392 19024 26444
rect 2136 26231 2188 26240
rect 2136 26197 2145 26231
rect 2145 26197 2179 26231
rect 2179 26197 2188 26231
rect 2136 26188 2188 26197
rect 4344 26188 4396 26240
rect 9220 26256 9272 26308
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 9496 26299 9548 26308
rect 9496 26265 9505 26299
rect 9505 26265 9539 26299
rect 9539 26265 9548 26299
rect 9496 26256 9548 26265
rect 13084 26256 13136 26308
rect 18052 26324 18104 26376
rect 21364 26324 21416 26376
rect 6552 26188 6604 26240
rect 9128 26188 9180 26240
rect 10600 26188 10652 26240
rect 13268 26231 13320 26240
rect 13268 26197 13277 26231
rect 13277 26197 13311 26231
rect 13311 26197 13320 26231
rect 13268 26188 13320 26197
rect 15660 26188 15712 26240
rect 19432 26256 19484 26308
rect 21456 26256 21508 26308
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 2136 25984 2188 26036
rect 2872 25916 2924 25968
rect 3056 25916 3108 25968
rect 2228 25848 2280 25900
rect 2320 25891 2372 25900
rect 2320 25857 2329 25891
rect 2329 25857 2363 25891
rect 2363 25857 2372 25891
rect 2320 25848 2372 25857
rect 3148 25848 3200 25900
rect 4252 25984 4304 26036
rect 4344 26027 4396 26036
rect 4344 25993 4353 26027
rect 4353 25993 4387 26027
rect 4387 25993 4396 26027
rect 4344 25984 4396 25993
rect 5356 25984 5408 26036
rect 6460 25984 6512 26036
rect 7472 25984 7524 26036
rect 2412 25712 2464 25764
rect 2872 25823 2924 25832
rect 2872 25789 2881 25823
rect 2881 25789 2915 25823
rect 2915 25789 2924 25823
rect 2872 25780 2924 25789
rect 3056 25780 3108 25832
rect 4528 25916 4580 25968
rect 4896 25916 4948 25968
rect 3700 25848 3752 25900
rect 3976 25848 4028 25900
rect 4712 25848 4764 25900
rect 6736 25916 6788 25968
rect 3056 25644 3108 25696
rect 4344 25712 4396 25764
rect 4896 25780 4948 25832
rect 7380 25891 7432 25900
rect 7380 25857 7389 25891
rect 7389 25857 7423 25891
rect 7423 25857 7432 25891
rect 7380 25848 7432 25857
rect 7748 25848 7800 25900
rect 8024 25848 8076 25900
rect 4528 25712 4580 25764
rect 6092 25712 6144 25764
rect 8208 25891 8260 25900
rect 8208 25857 8217 25891
rect 8217 25857 8251 25891
rect 8251 25857 8260 25891
rect 8208 25848 8260 25857
rect 10324 25984 10376 26036
rect 11244 25984 11296 26036
rect 13268 25984 13320 26036
rect 15752 26027 15804 26036
rect 15752 25993 15761 26027
rect 15761 25993 15795 26027
rect 15795 25993 15804 26027
rect 15752 25984 15804 25993
rect 15936 25984 15988 26036
rect 8484 25780 8536 25832
rect 9772 25780 9824 25832
rect 10416 25848 10468 25900
rect 12900 25848 12952 25900
rect 17224 25984 17276 26036
rect 10600 25780 10652 25832
rect 17684 25916 17736 25968
rect 18052 25959 18104 25968
rect 18052 25925 18061 25959
rect 18061 25925 18095 25959
rect 18095 25925 18104 25959
rect 18052 25916 18104 25925
rect 21456 26027 21508 26036
rect 21456 25993 21465 26027
rect 21465 25993 21499 26027
rect 21499 25993 21508 26027
rect 21456 25984 21508 25993
rect 15568 25780 15620 25832
rect 15752 25712 15804 25764
rect 16304 25712 16356 25764
rect 3516 25687 3568 25696
rect 3516 25653 3525 25687
rect 3525 25653 3559 25687
rect 3559 25653 3568 25687
rect 3516 25644 3568 25653
rect 3608 25644 3660 25696
rect 5264 25687 5316 25696
rect 5264 25653 5273 25687
rect 5273 25653 5307 25687
rect 5307 25653 5316 25687
rect 5264 25644 5316 25653
rect 6644 25644 6696 25696
rect 7564 25644 7616 25696
rect 7656 25644 7708 25696
rect 9036 25644 9088 25696
rect 10416 25687 10468 25696
rect 10416 25653 10425 25687
rect 10425 25653 10459 25687
rect 10459 25653 10468 25687
rect 10416 25644 10468 25653
rect 10968 25644 11020 25696
rect 12808 25644 12860 25696
rect 15476 25644 15528 25696
rect 16212 25644 16264 25696
rect 17316 25755 17368 25764
rect 17316 25721 17325 25755
rect 17325 25721 17359 25755
rect 17359 25721 17368 25755
rect 17316 25712 17368 25721
rect 18880 25848 18932 25900
rect 20812 25848 20864 25900
rect 18788 25823 18840 25832
rect 18788 25789 18797 25823
rect 18797 25789 18831 25823
rect 18831 25789 18840 25823
rect 18788 25780 18840 25789
rect 22560 25848 22612 25900
rect 21640 25712 21692 25764
rect 25780 25712 25832 25764
rect 19800 25644 19852 25696
rect 20260 25644 20312 25696
rect 25872 25644 25924 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 2320 25440 2372 25492
rect 3608 25440 3660 25492
rect 4344 25440 4396 25492
rect 5264 25440 5316 25492
rect 5356 25440 5408 25492
rect 2780 25304 2832 25356
rect 3332 25279 3384 25288
rect 3332 25245 3341 25279
rect 3341 25245 3375 25279
rect 3375 25245 3384 25279
rect 3332 25236 3384 25245
rect 6644 25372 6696 25424
rect 4804 25304 4856 25356
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 4252 25279 4304 25288
rect 4252 25245 4261 25279
rect 4261 25245 4295 25279
rect 4295 25245 4304 25279
rect 4252 25236 4304 25245
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 5724 25304 5776 25356
rect 5540 25236 5592 25288
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 8208 25440 8260 25492
rect 10416 25440 10468 25492
rect 10968 25483 11020 25492
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 16764 25440 16816 25492
rect 7288 25372 7340 25424
rect 7748 25372 7800 25424
rect 8392 25372 8444 25424
rect 3700 25100 3752 25152
rect 5356 25100 5408 25152
rect 5816 25100 5868 25152
rect 7380 25236 7432 25288
rect 7472 25236 7524 25288
rect 7564 25236 7616 25288
rect 6828 25168 6880 25220
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 9036 25304 9088 25356
rect 10600 25372 10652 25424
rect 8484 25236 8536 25288
rect 8576 25279 8628 25288
rect 8576 25245 8585 25279
rect 8585 25245 8619 25279
rect 8619 25245 8628 25279
rect 8576 25236 8628 25245
rect 8392 25168 8444 25220
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9588 25279 9640 25288
rect 9588 25245 9597 25279
rect 9597 25245 9631 25279
rect 9631 25245 9640 25279
rect 9588 25236 9640 25245
rect 9864 25236 9916 25288
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 7012 25143 7064 25152
rect 7012 25109 7021 25143
rect 7021 25109 7055 25143
rect 7055 25109 7064 25143
rect 7012 25100 7064 25109
rect 7288 25100 7340 25152
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 7748 25100 7800 25152
rect 8024 25100 8076 25152
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 11244 25236 11296 25288
rect 14740 25372 14792 25424
rect 18880 25440 18932 25492
rect 21640 25440 21692 25492
rect 20260 25372 20312 25424
rect 11796 25236 11848 25288
rect 11888 25279 11940 25288
rect 11888 25245 11897 25279
rect 11897 25245 11931 25279
rect 11931 25245 11940 25279
rect 11888 25236 11940 25245
rect 12440 25304 12492 25356
rect 12348 25236 12400 25288
rect 12808 25279 12860 25288
rect 12808 25245 12842 25279
rect 12842 25245 12860 25279
rect 12808 25236 12860 25245
rect 15476 25236 15528 25288
rect 15660 25279 15712 25288
rect 15660 25245 15694 25279
rect 15694 25245 15712 25279
rect 15660 25236 15712 25245
rect 13636 25100 13688 25152
rect 15936 25168 15988 25220
rect 16212 25168 16264 25220
rect 18788 25304 18840 25356
rect 19248 25304 19300 25356
rect 21364 25236 21416 25288
rect 13912 25143 13964 25152
rect 13912 25109 13921 25143
rect 13921 25109 13955 25143
rect 13955 25109 13964 25143
rect 13912 25100 13964 25109
rect 14648 25143 14700 25152
rect 14648 25109 14657 25143
rect 14657 25109 14691 25143
rect 14691 25109 14700 25143
rect 14648 25100 14700 25109
rect 16948 25100 17000 25152
rect 17408 25168 17460 25220
rect 17776 25168 17828 25220
rect 17868 25168 17920 25220
rect 17960 25100 18012 25152
rect 18880 25100 18932 25152
rect 21272 25168 21324 25220
rect 22468 25211 22520 25220
rect 22468 25177 22502 25211
rect 22502 25177 22520 25211
rect 22468 25168 22520 25177
rect 25780 25483 25832 25492
rect 25780 25449 25789 25483
rect 25789 25449 25823 25483
rect 25823 25449 25832 25483
rect 25780 25440 25832 25449
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 22376 25100 22428 25152
rect 24124 25211 24176 25220
rect 24124 25177 24133 25211
rect 24133 25177 24167 25211
rect 24167 25177 24176 25211
rect 24124 25168 24176 25177
rect 24308 25168 24360 25220
rect 23664 25143 23716 25152
rect 23664 25109 23673 25143
rect 23673 25109 23707 25143
rect 23707 25109 23716 25143
rect 23664 25100 23716 25109
rect 23756 25100 23808 25152
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 4160 24896 4212 24948
rect 6552 24896 6604 24948
rect 6644 24896 6696 24948
rect 7380 24896 7432 24948
rect 2228 24871 2280 24880
rect 2228 24837 2237 24871
rect 2237 24837 2271 24871
rect 2271 24837 2280 24871
rect 2228 24828 2280 24837
rect 2504 24760 2556 24812
rect 2320 24624 2372 24676
rect 2872 24624 2924 24676
rect 5264 24828 5316 24880
rect 6460 24828 6512 24880
rect 4988 24735 5040 24744
rect 4988 24701 4997 24735
rect 4997 24701 5031 24735
rect 5031 24701 5040 24735
rect 4988 24692 5040 24701
rect 1492 24556 1544 24608
rect 2780 24556 2832 24608
rect 3424 24556 3476 24608
rect 4068 24556 4120 24608
rect 4712 24556 4764 24608
rect 4896 24556 4948 24608
rect 5448 24599 5500 24608
rect 5448 24565 5457 24599
rect 5457 24565 5491 24599
rect 5491 24565 5500 24599
rect 5448 24556 5500 24565
rect 5540 24556 5592 24608
rect 5816 24760 5868 24812
rect 6276 24760 6328 24812
rect 7288 24828 7340 24880
rect 6828 24803 6880 24812
rect 6828 24769 6837 24803
rect 6837 24769 6871 24803
rect 6871 24769 6880 24803
rect 6828 24760 6880 24769
rect 7012 24760 7064 24812
rect 7196 24760 7248 24812
rect 7472 24760 7524 24812
rect 9864 24896 9916 24948
rect 8576 24828 8628 24880
rect 8852 24828 8904 24880
rect 9312 24871 9364 24880
rect 9312 24837 9321 24871
rect 9321 24837 9355 24871
rect 9355 24837 9364 24871
rect 9312 24828 9364 24837
rect 10324 24828 10376 24880
rect 9036 24760 9088 24812
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 8852 24692 8904 24744
rect 9496 24760 9548 24812
rect 7564 24624 7616 24676
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 10416 24803 10468 24812
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 10508 24760 10560 24812
rect 11888 24896 11940 24948
rect 17776 24939 17828 24948
rect 17776 24905 17785 24939
rect 17785 24905 17819 24939
rect 17819 24905 17828 24939
rect 17776 24896 17828 24905
rect 17960 24896 18012 24948
rect 21272 24939 21324 24948
rect 21272 24905 21281 24939
rect 21281 24905 21315 24939
rect 21315 24905 21324 24939
rect 21272 24896 21324 24905
rect 22468 24939 22520 24948
rect 22468 24905 22477 24939
rect 22477 24905 22511 24939
rect 22511 24905 22520 24939
rect 22468 24896 22520 24905
rect 23664 24896 23716 24948
rect 24308 24896 24360 24948
rect 10784 24871 10836 24880
rect 10784 24837 10809 24871
rect 10809 24837 10836 24871
rect 10784 24828 10836 24837
rect 14648 24828 14700 24880
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 12348 24760 12400 24812
rect 12440 24760 12492 24812
rect 12992 24760 13044 24812
rect 16580 24760 16632 24812
rect 16948 24871 17000 24880
rect 16948 24837 16957 24871
rect 16957 24837 16991 24871
rect 16991 24837 17000 24871
rect 16948 24828 17000 24837
rect 16856 24803 16908 24812
rect 15936 24735 15988 24744
rect 15936 24701 15945 24735
rect 15945 24701 15979 24735
rect 15979 24701 15988 24735
rect 15936 24692 15988 24701
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 7656 24556 7708 24608
rect 9772 24556 9824 24608
rect 9956 24556 10008 24608
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 16120 24556 16172 24608
rect 17132 24760 17184 24812
rect 17500 24803 17552 24812
rect 17500 24769 17509 24803
rect 17509 24769 17543 24803
rect 17543 24769 17552 24803
rect 17500 24760 17552 24769
rect 17868 24760 17920 24812
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20812 24828 20864 24880
rect 19248 24735 19300 24744
rect 19248 24701 19257 24735
rect 19257 24701 19291 24735
rect 19291 24701 19300 24735
rect 19248 24692 19300 24701
rect 22376 24692 22428 24744
rect 24124 24692 24176 24744
rect 25136 24692 25188 24744
rect 17132 24556 17184 24608
rect 17224 24599 17276 24608
rect 17224 24565 17233 24599
rect 17233 24565 17267 24599
rect 17267 24565 17276 24599
rect 17224 24556 17276 24565
rect 19524 24556 19576 24608
rect 24952 24667 25004 24676
rect 24952 24633 24961 24667
rect 24961 24633 24995 24667
rect 24995 24633 25004 24667
rect 24952 24624 25004 24633
rect 24768 24599 24820 24608
rect 24768 24565 24777 24599
rect 24777 24565 24811 24599
rect 24811 24565 24820 24599
rect 24768 24556 24820 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 2596 24395 2648 24404
rect 2596 24361 2605 24395
rect 2605 24361 2639 24395
rect 2639 24361 2648 24395
rect 2596 24352 2648 24361
rect 3332 24352 3384 24404
rect 4988 24352 5040 24404
rect 2320 24284 2372 24336
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 1952 24148 2004 24200
rect 2780 24216 2832 24268
rect 3240 24216 3292 24268
rect 2320 24191 2372 24200
rect 2320 24157 2329 24191
rect 2329 24157 2363 24191
rect 2363 24157 2372 24191
rect 2320 24148 2372 24157
rect 3700 24216 3752 24268
rect 3884 24216 3936 24268
rect 4896 24216 4948 24268
rect 2780 24080 2832 24132
rect 2964 24080 3016 24132
rect 3148 24080 3200 24132
rect 4344 24080 4396 24132
rect 4252 24055 4304 24064
rect 4252 24021 4261 24055
rect 4261 24021 4295 24055
rect 4295 24021 4304 24055
rect 4252 24012 4304 24021
rect 9588 24352 9640 24404
rect 15476 24352 15528 24404
rect 15752 24352 15804 24404
rect 5448 24284 5500 24336
rect 6000 24284 6052 24336
rect 5356 24148 5408 24200
rect 6828 24216 6880 24268
rect 10784 24284 10836 24336
rect 13912 24284 13964 24336
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 6368 24148 6420 24200
rect 9312 24216 9364 24268
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 7380 24148 7432 24200
rect 7472 24191 7524 24200
rect 7472 24157 7481 24191
rect 7481 24157 7515 24191
rect 7515 24157 7524 24191
rect 7472 24148 7524 24157
rect 6000 24080 6052 24132
rect 8760 24148 8812 24200
rect 9956 24148 10008 24200
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10324 24148 10376 24157
rect 11704 24216 11756 24268
rect 11796 24259 11848 24268
rect 11796 24225 11805 24259
rect 11805 24225 11839 24259
rect 11839 24225 11848 24259
rect 11796 24216 11848 24225
rect 6276 24012 6328 24064
rect 6736 24012 6788 24064
rect 7196 24012 7248 24064
rect 9036 24080 9088 24132
rect 9864 24123 9916 24132
rect 9864 24089 9873 24123
rect 9873 24089 9907 24123
rect 9907 24089 9916 24123
rect 10876 24148 10928 24200
rect 11888 24191 11940 24200
rect 9864 24080 9916 24089
rect 8576 24012 8628 24064
rect 10416 24012 10468 24064
rect 11244 24080 11296 24132
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12348 24148 12400 24200
rect 15568 24216 15620 24268
rect 13084 24080 13136 24132
rect 14464 24080 14516 24132
rect 14648 24080 14700 24132
rect 13728 24055 13780 24064
rect 13728 24021 13737 24055
rect 13737 24021 13771 24055
rect 13771 24021 13780 24055
rect 13728 24012 13780 24021
rect 15292 24012 15344 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 18972 24352 19024 24404
rect 21088 24284 21140 24336
rect 19248 24216 19300 24268
rect 17408 24148 17460 24200
rect 20812 24148 20864 24200
rect 17592 24123 17644 24132
rect 17592 24089 17626 24123
rect 17626 24089 17644 24123
rect 17592 24080 17644 24089
rect 18788 24080 18840 24132
rect 22744 24123 22796 24132
rect 22744 24089 22753 24123
rect 22753 24089 22787 24123
rect 22787 24089 22796 24123
rect 22744 24080 22796 24089
rect 22836 24123 22888 24132
rect 22836 24089 22845 24123
rect 22845 24089 22879 24123
rect 22879 24089 22888 24123
rect 22836 24080 22888 24089
rect 22284 24012 22336 24064
rect 23204 24148 23256 24200
rect 24400 24191 24452 24200
rect 24400 24157 24409 24191
rect 24409 24157 24443 24191
rect 24443 24157 24452 24191
rect 24400 24148 24452 24157
rect 23296 24080 23348 24132
rect 23020 24012 23072 24064
rect 24952 24012 25004 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 2228 23808 2280 23860
rect 2780 23808 2832 23860
rect 4252 23808 4304 23860
rect 5816 23808 5868 23860
rect 6000 23808 6052 23860
rect 6736 23851 6788 23860
rect 6736 23817 6745 23851
rect 6745 23817 6779 23851
rect 6779 23817 6788 23851
rect 6736 23808 6788 23817
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 2688 23740 2740 23792
rect 2320 23715 2372 23724
rect 2320 23681 2329 23715
rect 2329 23681 2363 23715
rect 2363 23681 2372 23715
rect 2320 23672 2372 23681
rect 2504 23536 2556 23588
rect 2228 23468 2280 23520
rect 3148 23672 3200 23724
rect 3148 23536 3200 23588
rect 3884 23672 3936 23724
rect 4068 23740 4120 23792
rect 4252 23672 4304 23724
rect 5632 23740 5684 23792
rect 5724 23740 5776 23792
rect 6644 23740 6696 23792
rect 7288 23783 7340 23792
rect 7288 23749 7297 23783
rect 7297 23749 7331 23783
rect 7331 23749 7340 23783
rect 7288 23740 7340 23749
rect 5356 23672 5408 23724
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 7012 23672 7064 23724
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 10876 23808 10928 23860
rect 12992 23808 13044 23860
rect 13728 23808 13780 23860
rect 16120 23851 16172 23860
rect 16120 23817 16129 23851
rect 16129 23817 16163 23851
rect 16163 23817 16172 23851
rect 16120 23808 16172 23817
rect 17592 23808 17644 23860
rect 9312 23740 9364 23792
rect 10140 23740 10192 23792
rect 10968 23740 11020 23792
rect 4068 23647 4120 23656
rect 4068 23613 4077 23647
rect 4077 23613 4111 23647
rect 4111 23613 4120 23647
rect 4068 23604 4120 23613
rect 4436 23604 4488 23656
rect 4988 23604 5040 23656
rect 5172 23647 5224 23656
rect 5172 23613 5181 23647
rect 5181 23613 5215 23647
rect 5215 23613 5224 23647
rect 5172 23604 5224 23613
rect 5448 23604 5500 23656
rect 5540 23647 5592 23656
rect 5540 23613 5549 23647
rect 5549 23613 5583 23647
rect 5583 23613 5592 23647
rect 5540 23604 5592 23613
rect 5632 23647 5684 23656
rect 5632 23613 5641 23647
rect 5641 23613 5675 23647
rect 5675 23613 5684 23647
rect 5632 23604 5684 23613
rect 5724 23647 5776 23656
rect 5724 23613 5733 23647
rect 5733 23613 5767 23647
rect 5767 23613 5776 23647
rect 5724 23604 5776 23613
rect 6184 23604 6236 23656
rect 6736 23604 6788 23656
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 8392 23672 8444 23724
rect 10048 23672 10100 23724
rect 10324 23604 10376 23656
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 15292 23740 15344 23792
rect 15568 23740 15620 23792
rect 19708 23740 19760 23792
rect 23204 23851 23256 23860
rect 23204 23817 23213 23851
rect 23213 23817 23247 23851
rect 23247 23817 23256 23851
rect 23204 23808 23256 23817
rect 24768 23808 24820 23860
rect 22928 23740 22980 23792
rect 7472 23536 7524 23588
rect 8208 23536 8260 23588
rect 16120 23604 16172 23656
rect 16672 23604 16724 23656
rect 17132 23604 17184 23656
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 21364 23672 21416 23724
rect 22652 23672 22704 23724
rect 23480 23715 23532 23724
rect 23480 23681 23484 23715
rect 23484 23681 23518 23715
rect 23518 23681 23532 23715
rect 23480 23672 23532 23681
rect 23756 23715 23808 23724
rect 23756 23681 23801 23715
rect 23801 23681 23808 23715
rect 23756 23672 23808 23681
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 24400 23604 24452 23656
rect 16856 23536 16908 23588
rect 19340 23536 19392 23588
rect 3976 23468 4028 23520
rect 4804 23468 4856 23520
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 7288 23468 7340 23520
rect 7748 23468 7800 23520
rect 7840 23468 7892 23520
rect 8668 23468 8720 23520
rect 8944 23468 8996 23520
rect 9404 23468 9456 23520
rect 10876 23511 10928 23520
rect 10876 23477 10885 23511
rect 10885 23477 10919 23511
rect 10919 23477 10928 23511
rect 10876 23468 10928 23477
rect 12072 23468 12124 23520
rect 14464 23511 14516 23520
rect 14464 23477 14473 23511
rect 14473 23477 14507 23511
rect 14507 23477 14516 23511
rect 14464 23468 14516 23477
rect 16028 23511 16080 23520
rect 16028 23477 16037 23511
rect 16037 23477 16071 23511
rect 16071 23477 16080 23511
rect 16028 23468 16080 23477
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 18880 23511 18932 23520
rect 18880 23477 18889 23511
rect 18889 23477 18923 23511
rect 18923 23477 18932 23511
rect 18880 23468 18932 23477
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 19984 23511 20036 23520
rect 19984 23477 19993 23511
rect 19993 23477 20027 23511
rect 20027 23477 20036 23511
rect 19984 23468 20036 23477
rect 21088 23468 21140 23520
rect 21640 23468 21692 23520
rect 22468 23468 22520 23520
rect 26332 23511 26384 23520
rect 26332 23477 26341 23511
rect 26341 23477 26375 23511
rect 26375 23477 26384 23511
rect 26332 23468 26384 23477
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 2964 23264 3016 23316
rect 5632 23264 5684 23316
rect 7196 23264 7248 23316
rect 2136 23196 2188 23248
rect 2596 23196 2648 23248
rect 6920 23196 6972 23248
rect 1584 23128 1636 23180
rect 1860 23060 1912 23112
rect 2964 23060 3016 23112
rect 8484 23264 8536 23316
rect 9496 23264 9548 23316
rect 10232 23264 10284 23316
rect 10508 23307 10560 23316
rect 10508 23273 10517 23307
rect 10517 23273 10551 23307
rect 10551 23273 10560 23307
rect 10508 23264 10560 23273
rect 11244 23307 11296 23316
rect 11244 23273 11253 23307
rect 11253 23273 11287 23307
rect 11287 23273 11296 23307
rect 11244 23264 11296 23273
rect 13912 23264 13964 23316
rect 15476 23264 15528 23316
rect 18788 23307 18840 23316
rect 18788 23273 18797 23307
rect 18797 23273 18831 23307
rect 18831 23273 18840 23307
rect 18788 23264 18840 23273
rect 8392 23239 8444 23248
rect 8392 23205 8401 23239
rect 8401 23205 8435 23239
rect 8435 23205 8444 23239
rect 8392 23196 8444 23205
rect 9956 23196 10008 23248
rect 10876 23196 10928 23248
rect 19340 23264 19392 23316
rect 19432 23307 19484 23316
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 20628 23264 20680 23316
rect 21272 23264 21324 23316
rect 23940 23264 23992 23316
rect 18972 23196 19024 23248
rect 20168 23239 20220 23248
rect 20168 23205 20177 23239
rect 20177 23205 20211 23239
rect 20211 23205 20220 23239
rect 20168 23196 20220 23205
rect 22836 23196 22888 23248
rect 23388 23196 23440 23248
rect 1952 22992 2004 23044
rect 2688 22992 2740 23044
rect 2504 22924 2556 22976
rect 3424 23060 3476 23112
rect 4988 23060 5040 23112
rect 5540 22924 5592 22976
rect 6644 23060 6696 23112
rect 7748 23060 7800 23112
rect 7840 23060 7892 23112
rect 9036 23128 9088 23180
rect 9864 23128 9916 23180
rect 6092 23035 6144 23044
rect 6092 23001 6101 23035
rect 6101 23001 6135 23035
rect 6135 23001 6144 23035
rect 6092 22992 6144 23001
rect 6828 22924 6880 22976
rect 7564 22924 7616 22976
rect 10048 23103 10100 23112
rect 10048 23069 10057 23103
rect 10057 23069 10091 23103
rect 10091 23069 10100 23103
rect 10048 23060 10100 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10324 23060 10376 23069
rect 10968 23128 11020 23180
rect 9680 22992 9732 23044
rect 8668 22924 8720 22976
rect 9036 22924 9088 22976
rect 12900 22992 12952 23044
rect 12992 22992 13044 23044
rect 14648 23060 14700 23112
rect 11520 22924 11572 22976
rect 11612 22924 11664 22976
rect 16856 23128 16908 23180
rect 15292 23060 15344 23112
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 15200 22924 15252 22976
rect 17040 23060 17092 23112
rect 17408 23060 17460 23112
rect 19340 23060 19392 23112
rect 22192 23060 22244 23112
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 22376 23103 22428 23112
rect 22376 23069 22386 23103
rect 22386 23069 22420 23103
rect 22420 23069 22428 23103
rect 22376 23060 22428 23069
rect 22652 23128 22704 23180
rect 22836 23060 22888 23112
rect 18604 23035 18656 23044
rect 18604 23001 18613 23035
rect 18613 23001 18647 23035
rect 18647 23001 18656 23035
rect 18604 22992 18656 23001
rect 16396 22967 16448 22976
rect 16396 22933 16405 22967
rect 16405 22933 16439 22967
rect 16439 22933 16448 22967
rect 16396 22924 16448 22933
rect 17408 22924 17460 22976
rect 18144 22924 18196 22976
rect 19816 23035 19868 23044
rect 19816 23001 19843 23035
rect 19843 23001 19868 23035
rect 19816 22992 19868 23001
rect 20536 22992 20588 23044
rect 21272 23035 21324 23044
rect 21272 23001 21281 23035
rect 21281 23001 21315 23035
rect 21315 23001 21324 23035
rect 21272 22992 21324 23001
rect 23020 22992 23072 23044
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 23480 23060 23532 23112
rect 24400 23103 24452 23112
rect 24400 23069 24409 23103
rect 24409 23069 24443 23103
rect 24443 23069 24452 23103
rect 24400 23060 24452 23069
rect 24952 23060 25004 23112
rect 18788 22967 18840 22976
rect 18788 22933 18813 22967
rect 18813 22933 18840 22967
rect 18788 22924 18840 22933
rect 18972 22967 19024 22976
rect 18972 22933 18981 22967
rect 18981 22933 19015 22967
rect 19015 22933 19024 22967
rect 18972 22924 19024 22933
rect 19432 22967 19484 22976
rect 19432 22933 19459 22967
rect 19459 22933 19484 22967
rect 19432 22924 19484 22933
rect 20720 22924 20772 22976
rect 22192 22924 22244 22976
rect 23940 22992 23992 23044
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 1768 22720 1820 22772
rect 2320 22720 2372 22772
rect 2596 22763 2648 22772
rect 2596 22729 2605 22763
rect 2605 22729 2639 22763
rect 2639 22729 2648 22763
rect 2596 22720 2648 22729
rect 2780 22720 2832 22772
rect 3700 22720 3752 22772
rect 4252 22720 4304 22772
rect 5540 22720 5592 22772
rect 6000 22720 6052 22772
rect 6368 22720 6420 22772
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2872 22652 2924 22704
rect 7472 22720 7524 22772
rect 8392 22720 8444 22772
rect 2228 22516 2280 22568
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 3332 22627 3384 22636
rect 3332 22593 3341 22627
rect 3341 22593 3375 22627
rect 3375 22593 3384 22627
rect 3332 22584 3384 22593
rect 3056 22516 3108 22568
rect 3884 22584 3936 22636
rect 4804 22584 4856 22636
rect 5356 22627 5408 22636
rect 5356 22593 5365 22627
rect 5365 22593 5399 22627
rect 5399 22593 5408 22627
rect 5356 22584 5408 22593
rect 7748 22652 7800 22704
rect 2964 22448 3016 22500
rect 4344 22448 4396 22500
rect 1952 22423 2004 22432
rect 1952 22389 1961 22423
rect 1961 22389 1995 22423
rect 1995 22389 2004 22423
rect 1952 22380 2004 22389
rect 2136 22423 2188 22432
rect 2136 22389 2145 22423
rect 2145 22389 2179 22423
rect 2179 22389 2188 22423
rect 2136 22380 2188 22389
rect 4252 22380 4304 22432
rect 4896 22380 4948 22432
rect 6000 22584 6052 22636
rect 6460 22380 6512 22432
rect 7012 22627 7064 22636
rect 7012 22593 7057 22627
rect 7057 22593 7064 22627
rect 7012 22584 7064 22593
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 8024 22584 8076 22636
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 8392 22516 8444 22568
rect 7472 22380 7524 22432
rect 8668 22448 8720 22500
rect 9312 22720 9364 22772
rect 11520 22763 11572 22772
rect 11520 22729 11529 22763
rect 11529 22729 11563 22763
rect 11563 22729 11572 22763
rect 11520 22720 11572 22729
rect 11704 22720 11756 22772
rect 12900 22763 12952 22772
rect 12900 22729 12909 22763
rect 12909 22729 12943 22763
rect 12943 22729 12952 22763
rect 12900 22720 12952 22729
rect 15476 22720 15528 22772
rect 16764 22720 16816 22772
rect 17224 22720 17276 22772
rect 9036 22516 9088 22568
rect 11888 22584 11940 22636
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 10876 22516 10928 22568
rect 11244 22516 11296 22568
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 11796 22516 11848 22568
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12716 22627 12768 22636
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 13360 22627 13412 22636
rect 13360 22593 13369 22627
rect 13369 22593 13403 22627
rect 13403 22593 13412 22627
rect 13360 22584 13412 22593
rect 15752 22652 15804 22704
rect 15476 22584 15528 22636
rect 15384 22516 15436 22568
rect 15660 22516 15712 22568
rect 9128 22448 9180 22500
rect 12072 22380 12124 22432
rect 12256 22380 12308 22432
rect 13176 22491 13228 22500
rect 13176 22457 13185 22491
rect 13185 22457 13219 22491
rect 13219 22457 13228 22491
rect 17776 22584 17828 22636
rect 16120 22516 16172 22568
rect 18144 22516 18196 22568
rect 18972 22652 19024 22704
rect 19616 22720 19668 22772
rect 23940 22763 23992 22772
rect 23940 22729 23949 22763
rect 23949 22729 23983 22763
rect 23983 22729 23992 22763
rect 23940 22720 23992 22729
rect 25780 22720 25832 22772
rect 18696 22584 18748 22636
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 20720 22652 20772 22704
rect 22284 22652 22336 22704
rect 24492 22695 24544 22704
rect 19524 22627 19576 22636
rect 19524 22593 19533 22627
rect 19533 22593 19567 22627
rect 19567 22593 19576 22627
rect 19524 22584 19576 22593
rect 24492 22661 24501 22695
rect 24501 22661 24535 22695
rect 24535 22661 24544 22695
rect 24492 22652 24544 22661
rect 25136 22652 25188 22704
rect 18972 22559 19024 22568
rect 18972 22525 18981 22559
rect 18981 22525 19015 22559
rect 19015 22525 19024 22559
rect 18972 22516 19024 22525
rect 13176 22448 13228 22457
rect 13084 22380 13136 22432
rect 14740 22380 14792 22432
rect 17040 22380 17092 22432
rect 18052 22380 18104 22432
rect 19432 22448 19484 22500
rect 22744 22516 22796 22568
rect 26332 22448 26384 22500
rect 18788 22380 18840 22432
rect 19984 22380 20036 22432
rect 20444 22380 20496 22432
rect 24952 22423 25004 22432
rect 24952 22389 24961 22423
rect 24961 22389 24995 22423
rect 24995 22389 25004 22423
rect 24952 22380 25004 22389
rect 25688 22423 25740 22432
rect 25688 22389 25697 22423
rect 25697 22389 25731 22423
rect 25731 22389 25740 22423
rect 25688 22380 25740 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 1676 22176 1728 22228
rect 1952 22176 2004 22228
rect 3976 22176 4028 22228
rect 2320 22108 2372 22160
rect 3792 22108 3844 22160
rect 2780 22040 2832 22092
rect 3516 22040 3568 22092
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2136 21972 2188 22024
rect 5724 22176 5776 22228
rect 3424 21904 3476 21956
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 6644 22176 6696 22228
rect 7748 22176 7800 22228
rect 8300 22219 8352 22228
rect 8300 22185 8309 22219
rect 8309 22185 8343 22219
rect 8343 22185 8352 22219
rect 8300 22176 8352 22185
rect 10968 22176 11020 22228
rect 6368 22108 6420 22160
rect 4712 21972 4764 22024
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 6184 22083 6236 22092
rect 6184 22049 6193 22083
rect 6193 22049 6227 22083
rect 6227 22049 6236 22083
rect 6184 22040 6236 22049
rect 6828 22108 6880 22160
rect 8024 22108 8076 22160
rect 8668 22108 8720 22160
rect 11704 22176 11756 22228
rect 11980 22176 12032 22228
rect 12256 22219 12308 22228
rect 12256 22185 12265 22219
rect 12265 22185 12299 22219
rect 12299 22185 12308 22219
rect 12256 22176 12308 22185
rect 15292 22176 15344 22228
rect 5540 21972 5592 21981
rect 5816 22015 5868 22024
rect 5816 21981 5825 22015
rect 5825 21981 5859 22015
rect 5859 21981 5868 22015
rect 5816 21972 5868 21981
rect 5908 21972 5960 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 9312 22040 9364 22092
rect 11612 22108 11664 22160
rect 19340 22176 19392 22228
rect 19616 22219 19668 22228
rect 19616 22185 19625 22219
rect 19625 22185 19659 22219
rect 19659 22185 19668 22219
rect 19616 22176 19668 22185
rect 19984 22176 20036 22228
rect 20812 22176 20864 22228
rect 18696 22108 18748 22160
rect 19156 22108 19208 22160
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6644 21972 6696 21981
rect 8208 21972 8260 22024
rect 6184 21904 6236 21956
rect 6460 21904 6512 21956
rect 7012 21947 7064 21956
rect 7012 21913 7021 21947
rect 7021 21913 7055 21947
rect 7055 21913 7064 21947
rect 7012 21904 7064 21913
rect 9956 21904 10008 21956
rect 2136 21879 2188 21888
rect 2136 21845 2145 21879
rect 2145 21845 2179 21879
rect 2179 21845 2188 21879
rect 2136 21836 2188 21845
rect 4988 21879 5040 21888
rect 4988 21845 4997 21879
rect 4997 21845 5031 21879
rect 5031 21845 5040 21879
rect 4988 21836 5040 21845
rect 5356 21836 5408 21888
rect 6000 21836 6052 21888
rect 6828 21836 6880 21888
rect 7380 21836 7432 21888
rect 10416 21904 10468 21956
rect 10876 21972 10928 22024
rect 10968 22015 11020 22024
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 16028 22083 16080 22092
rect 16028 22049 16037 22083
rect 16037 22049 16071 22083
rect 16071 22049 16080 22083
rect 16028 22040 16080 22049
rect 11244 21947 11296 21956
rect 11244 21913 11279 21947
rect 11279 21913 11296 21947
rect 11704 22015 11756 22024
rect 11704 21981 11713 22015
rect 11713 21981 11747 22015
rect 11747 21981 11756 22015
rect 11704 21972 11756 21981
rect 11796 21972 11848 22024
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 13360 21972 13412 22024
rect 14740 21972 14792 22024
rect 15752 21972 15804 22024
rect 16948 21972 17000 22024
rect 18880 21972 18932 22024
rect 19340 21972 19392 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 20260 22040 20312 22092
rect 19432 21972 19484 21981
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 20444 22108 20496 22160
rect 21088 22040 21140 22092
rect 22744 22219 22796 22228
rect 22744 22185 22753 22219
rect 22753 22185 22787 22219
rect 22787 22185 22796 22219
rect 22744 22176 22796 22185
rect 22836 22219 22888 22228
rect 22836 22185 22845 22219
rect 22845 22185 22879 22219
rect 22879 22185 22888 22219
rect 22836 22176 22888 22185
rect 26332 22176 26384 22228
rect 23572 22108 23624 22160
rect 19892 21972 19944 21981
rect 11244 21904 11296 21913
rect 12532 21904 12584 21956
rect 13176 21947 13228 21956
rect 13176 21913 13185 21947
rect 13185 21913 13219 21947
rect 13219 21913 13228 21947
rect 13176 21904 13228 21913
rect 11060 21836 11112 21888
rect 11612 21836 11664 21888
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 16672 21904 16724 21956
rect 17776 21904 17828 21956
rect 18328 21904 18380 21956
rect 19524 21904 19576 21956
rect 19616 21904 19668 21956
rect 22928 21972 22980 22024
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 23296 21972 23348 22024
rect 14648 21879 14700 21888
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 15292 21836 15344 21888
rect 16304 21836 16356 21888
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 17592 21836 17644 21888
rect 17960 21836 18012 21888
rect 19984 21836 20036 21888
rect 20536 21836 20588 21888
rect 20628 21879 20680 21888
rect 20628 21845 20637 21879
rect 20637 21845 20671 21879
rect 20671 21845 20680 21879
rect 20628 21836 20680 21845
rect 21456 21904 21508 21956
rect 22652 21836 22704 21888
rect 23480 21879 23532 21888
rect 23480 21845 23497 21879
rect 23497 21845 23532 21879
rect 23480 21836 23532 21845
rect 24952 21972 25004 22024
rect 24860 21879 24912 21888
rect 24860 21845 24869 21879
rect 24869 21845 24903 21879
rect 24903 21845 24912 21879
rect 24860 21836 24912 21845
rect 26332 22015 26384 22024
rect 26332 21981 26341 22015
rect 26341 21981 26375 22015
rect 26375 21981 26384 22015
rect 26332 21972 26384 21981
rect 26148 21904 26200 21956
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 2596 21632 2648 21684
rect 3056 21632 3108 21684
rect 3332 21632 3384 21684
rect 2228 21564 2280 21616
rect 2780 21607 2832 21616
rect 2780 21573 2812 21607
rect 2812 21573 2832 21607
rect 2780 21564 2832 21573
rect 2136 21428 2188 21480
rect 4160 21632 4212 21684
rect 4344 21632 4396 21684
rect 5448 21632 5500 21684
rect 5264 21564 5316 21616
rect 6460 21675 6512 21684
rect 6460 21641 6469 21675
rect 6469 21641 6503 21675
rect 6503 21641 6512 21675
rect 6460 21632 6512 21641
rect 7472 21632 7524 21684
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4160 21428 4212 21480
rect 4344 21539 4396 21548
rect 4344 21505 4353 21539
rect 4353 21505 4387 21539
rect 4387 21505 4396 21539
rect 4344 21496 4396 21505
rect 1308 21360 1360 21412
rect 4252 21360 4304 21412
rect 4804 21496 4856 21548
rect 5448 21496 5500 21548
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 4896 21471 4948 21480
rect 4896 21437 4905 21471
rect 4905 21437 4939 21471
rect 4939 21437 4948 21471
rect 4896 21428 4948 21437
rect 5356 21428 5408 21480
rect 6184 21607 6236 21616
rect 6184 21573 6193 21607
rect 6193 21573 6227 21607
rect 6227 21573 6236 21607
rect 6184 21564 6236 21573
rect 6736 21607 6788 21616
rect 6736 21573 6745 21607
rect 6745 21573 6779 21607
rect 6779 21573 6788 21607
rect 6736 21564 6788 21573
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 7288 21496 7340 21548
rect 7472 21539 7524 21582
rect 7472 21530 7481 21539
rect 7481 21530 7515 21539
rect 7515 21530 7524 21539
rect 8484 21632 8536 21684
rect 8300 21564 8352 21616
rect 5540 21360 5592 21412
rect 2320 21292 2372 21344
rect 3240 21292 3292 21344
rect 4804 21335 4856 21344
rect 4804 21301 4813 21335
rect 4813 21301 4847 21335
rect 4847 21301 4856 21335
rect 4804 21292 4856 21301
rect 5908 21360 5960 21412
rect 7196 21428 7248 21480
rect 6920 21292 6972 21344
rect 7564 21428 7616 21480
rect 8484 21539 8536 21548
rect 8484 21505 8493 21539
rect 8493 21505 8527 21539
rect 8527 21505 8536 21539
rect 8484 21496 8536 21505
rect 9404 21632 9456 21684
rect 9772 21632 9824 21684
rect 9864 21564 9916 21616
rect 8392 21428 8444 21480
rect 9588 21471 9640 21480
rect 9588 21437 9597 21471
rect 9597 21437 9631 21471
rect 9631 21437 9640 21471
rect 9588 21428 9640 21437
rect 9956 21496 10008 21548
rect 9772 21360 9824 21412
rect 9864 21403 9916 21412
rect 9864 21369 9873 21403
rect 9873 21369 9907 21403
rect 9907 21369 9916 21403
rect 9864 21360 9916 21369
rect 10968 21632 11020 21684
rect 12532 21632 12584 21684
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 17960 21632 18012 21684
rect 19432 21632 19484 21684
rect 19524 21632 19576 21684
rect 20260 21632 20312 21684
rect 23480 21632 23532 21684
rect 26148 21632 26200 21684
rect 11060 21496 11112 21548
rect 11888 21428 11940 21480
rect 12808 21496 12860 21548
rect 13176 21539 13228 21548
rect 13176 21505 13210 21539
rect 13210 21505 13228 21539
rect 13176 21496 13228 21505
rect 14648 21564 14700 21616
rect 15660 21564 15712 21616
rect 12532 21428 12584 21480
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 16304 21496 16356 21548
rect 17224 21496 17276 21548
rect 17684 21496 17736 21548
rect 19892 21496 19944 21548
rect 20628 21564 20680 21616
rect 22284 21564 22336 21616
rect 7564 21292 7616 21344
rect 7656 21292 7708 21344
rect 9128 21292 9180 21344
rect 10784 21292 10836 21344
rect 11796 21292 11848 21344
rect 12900 21292 12952 21344
rect 13636 21292 13688 21344
rect 14832 21292 14884 21344
rect 16580 21292 16632 21344
rect 18328 21428 18380 21480
rect 19156 21428 19208 21480
rect 19800 21428 19852 21480
rect 18144 21292 18196 21344
rect 18880 21292 18932 21344
rect 19340 21335 19392 21344
rect 19340 21301 19349 21335
rect 19349 21301 19383 21335
rect 19383 21301 19392 21335
rect 19340 21292 19392 21301
rect 19432 21292 19484 21344
rect 19892 21292 19944 21344
rect 21272 21292 21324 21344
rect 22560 21428 22612 21480
rect 22744 21496 22796 21548
rect 23204 21607 23256 21616
rect 23204 21573 23213 21607
rect 23213 21573 23247 21607
rect 23247 21573 23256 21607
rect 23204 21564 23256 21573
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 24860 21428 24912 21480
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 22652 21335 22704 21344
rect 22652 21301 22661 21335
rect 22661 21301 22695 21335
rect 22695 21301 22704 21335
rect 22652 21292 22704 21301
rect 22836 21335 22888 21344
rect 22836 21301 22845 21335
rect 22845 21301 22879 21335
rect 22879 21301 22888 21335
rect 22836 21292 22888 21301
rect 23112 21360 23164 21412
rect 23204 21292 23256 21344
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 2412 21088 2464 21140
rect 2780 21088 2832 21140
rect 4896 21088 4948 21140
rect 3056 21020 3108 21072
rect 3516 21020 3568 21072
rect 2688 20995 2740 21004
rect 2688 20961 2697 20995
rect 2697 20961 2731 20995
rect 2731 20961 2740 20995
rect 2688 20952 2740 20961
rect 3240 20995 3292 21004
rect 3240 20961 3249 20995
rect 3249 20961 3283 20995
rect 3283 20961 3292 20995
rect 3240 20952 3292 20961
rect 3148 20884 3200 20936
rect 4160 20884 4212 20936
rect 5172 20884 5224 20936
rect 5540 21088 5592 21140
rect 6276 21088 6328 21140
rect 7104 21088 7156 21140
rect 7196 21088 7248 21140
rect 6184 20884 6236 20936
rect 6644 20927 6696 20936
rect 6644 20893 6650 20927
rect 6650 20893 6684 20927
rect 6684 20893 6696 20927
rect 6644 20884 6696 20893
rect 6920 20952 6972 21004
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 7656 20927 7708 20936
rect 8760 21131 8812 21140
rect 8760 21097 8769 21131
rect 8769 21097 8803 21131
rect 8803 21097 8812 21131
rect 8760 21088 8812 21097
rect 9128 21131 9180 21140
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 8852 21020 8904 21072
rect 9496 21020 9548 21072
rect 9864 21020 9916 21072
rect 9404 20952 9456 21004
rect 7656 20893 7701 20927
rect 7701 20893 7708 20927
rect 7656 20884 7708 20893
rect 9220 20884 9272 20936
rect 9588 20884 9640 20936
rect 4712 20816 4764 20868
rect 2320 20748 2372 20800
rect 4620 20748 4672 20800
rect 5816 20748 5868 20800
rect 6552 20748 6604 20800
rect 8760 20816 8812 20868
rect 8852 20816 8904 20868
rect 13176 21088 13228 21140
rect 14740 21088 14792 21140
rect 15200 21131 15252 21140
rect 15200 21097 15209 21131
rect 15209 21097 15243 21131
rect 15243 21097 15252 21131
rect 15200 21088 15252 21097
rect 12808 21020 12860 21072
rect 14832 21020 14884 21072
rect 17500 21088 17552 21140
rect 18696 21131 18748 21140
rect 18696 21097 18705 21131
rect 18705 21097 18739 21131
rect 18739 21097 18748 21131
rect 18696 21088 18748 21097
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 19156 21088 19208 21140
rect 19340 21088 19392 21140
rect 21180 21088 21232 21140
rect 21456 21131 21508 21140
rect 21456 21097 21465 21131
rect 21465 21097 21499 21131
rect 21499 21097 21508 21131
rect 21456 21088 21508 21097
rect 22836 21131 22888 21140
rect 22836 21097 22845 21131
rect 22845 21097 22879 21131
rect 22879 21097 22888 21131
rect 22836 21088 22888 21097
rect 23112 21088 23164 21140
rect 23664 21088 23716 21140
rect 24860 21088 24912 21140
rect 19248 21020 19300 21072
rect 20444 21020 20496 21072
rect 10784 20884 10836 20936
rect 11244 20927 11296 20936
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 7380 20748 7432 20800
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 9772 20748 9824 20800
rect 11704 20816 11756 20868
rect 13360 20816 13412 20868
rect 14832 20884 14884 20936
rect 14372 20816 14424 20868
rect 14648 20816 14700 20868
rect 15476 20884 15528 20936
rect 16580 20884 16632 20936
rect 19984 20952 20036 21004
rect 20352 20952 20404 21004
rect 16120 20816 16172 20868
rect 16488 20816 16540 20868
rect 18972 20884 19024 20936
rect 11060 20748 11112 20800
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 14004 20748 14056 20800
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 14740 20748 14792 20800
rect 15200 20748 15252 20800
rect 16764 20748 16816 20800
rect 18696 20816 18748 20868
rect 19340 20884 19392 20936
rect 19524 20816 19576 20868
rect 20904 20816 20956 20868
rect 21088 20816 21140 20868
rect 17684 20748 17736 20800
rect 19064 20748 19116 20800
rect 19984 20791 20036 20800
rect 19984 20757 19993 20791
rect 19993 20757 20027 20791
rect 20027 20757 20036 20791
rect 19984 20748 20036 20757
rect 20076 20748 20128 20800
rect 21180 20748 21232 20800
rect 22284 20952 22336 21004
rect 22836 20952 22888 21004
rect 22560 20884 22612 20936
rect 22928 20884 22980 20936
rect 23112 20816 23164 20868
rect 24492 20952 24544 21004
rect 23020 20791 23072 20800
rect 23020 20757 23037 20791
rect 23037 20757 23072 20791
rect 23020 20748 23072 20757
rect 23756 20791 23808 20800
rect 23756 20757 23765 20791
rect 23765 20757 23799 20791
rect 23799 20757 23808 20791
rect 23756 20748 23808 20757
rect 25136 20748 25188 20800
rect 26240 20748 26292 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 3148 20544 3200 20596
rect 3608 20544 3660 20596
rect 4344 20544 4396 20596
rect 3148 20340 3200 20392
rect 3240 20340 3292 20392
rect 3332 20340 3384 20392
rect 4160 20476 4212 20528
rect 4988 20544 5040 20596
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 6092 20544 6144 20596
rect 7104 20544 7156 20596
rect 11244 20544 11296 20596
rect 6184 20519 6236 20528
rect 6184 20485 6193 20519
rect 6193 20485 6227 20519
rect 6227 20485 6236 20519
rect 6184 20476 6236 20485
rect 4712 20451 4764 20460
rect 4712 20417 4721 20451
rect 4721 20417 4755 20451
rect 4755 20417 4764 20451
rect 4712 20408 4764 20417
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 3240 20204 3292 20256
rect 3608 20204 3660 20256
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4896 20340 4948 20392
rect 4252 20272 4304 20324
rect 5264 20408 5316 20460
rect 6828 20476 6880 20528
rect 7840 20476 7892 20528
rect 13268 20544 13320 20596
rect 16488 20544 16540 20596
rect 17960 20544 18012 20596
rect 12992 20476 13044 20528
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 6552 20408 6604 20460
rect 6736 20408 6788 20460
rect 7380 20408 7432 20460
rect 7472 20408 7524 20460
rect 6184 20340 6236 20392
rect 8484 20340 8536 20392
rect 9404 20408 9456 20460
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 9772 20272 9824 20324
rect 13176 20408 13228 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 14648 20476 14700 20528
rect 13452 20340 13504 20392
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 14096 20408 14148 20460
rect 14740 20408 14792 20460
rect 15200 20476 15252 20528
rect 15660 20408 15712 20460
rect 16212 20476 16264 20528
rect 18144 20476 18196 20528
rect 19340 20544 19392 20596
rect 22100 20476 22152 20528
rect 13636 20340 13688 20392
rect 15568 20340 15620 20392
rect 13820 20272 13872 20324
rect 14280 20315 14332 20324
rect 14280 20281 14289 20315
rect 14289 20281 14323 20315
rect 14323 20281 14332 20315
rect 14280 20272 14332 20281
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17868 20408 17920 20460
rect 18696 20408 18748 20460
rect 19984 20408 20036 20460
rect 20720 20408 20772 20460
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 26332 20544 26384 20596
rect 23756 20476 23808 20528
rect 26240 20476 26292 20528
rect 22284 20408 22336 20460
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 6092 20204 6144 20256
rect 7656 20204 7708 20256
rect 9220 20204 9272 20256
rect 10968 20204 11020 20256
rect 14924 20247 14976 20256
rect 14924 20213 14933 20247
rect 14933 20213 14967 20247
rect 14967 20213 14976 20247
rect 14924 20204 14976 20213
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15384 20204 15436 20213
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 16488 20247 16540 20256
rect 16488 20213 16497 20247
rect 16497 20213 16531 20247
rect 16531 20213 16540 20247
rect 16488 20204 16540 20213
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 17132 20204 17184 20256
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 22928 20408 22980 20460
rect 24952 20408 25004 20460
rect 19156 20272 19208 20324
rect 18972 20204 19024 20256
rect 20076 20204 20128 20256
rect 20628 20204 20680 20256
rect 22100 20204 22152 20256
rect 22744 20204 22796 20256
rect 22928 20204 22980 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 2596 20000 2648 20052
rect 2688 20000 2740 20052
rect 3148 20000 3200 20052
rect 3424 20000 3476 20052
rect 6920 20000 6972 20052
rect 7656 20000 7708 20052
rect 8392 20000 8444 20052
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 9036 20000 9088 20052
rect 9864 20000 9916 20052
rect 10324 20043 10376 20052
rect 10324 20009 10333 20043
rect 10333 20009 10367 20043
rect 10367 20009 10376 20043
rect 10324 20000 10376 20009
rect 10876 20000 10928 20052
rect 11060 20000 11112 20052
rect 11704 20000 11756 20052
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 2964 19932 3016 19984
rect 3240 19932 3292 19984
rect 3884 19932 3936 19984
rect 2320 19864 2372 19916
rect 756 19728 808 19780
rect 2504 19796 2556 19848
rect 4068 19864 4120 19916
rect 5632 19932 5684 19984
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3240 19796 3292 19805
rect 3424 19796 3476 19848
rect 3884 19839 3936 19848
rect 3884 19805 3893 19839
rect 3893 19805 3927 19839
rect 3927 19805 3936 19839
rect 3884 19796 3936 19805
rect 4344 19839 4396 19848
rect 4344 19805 4353 19839
rect 4353 19805 4387 19839
rect 4387 19805 4396 19839
rect 4344 19796 4396 19805
rect 5816 19907 5868 19916
rect 5816 19873 5825 19907
rect 5825 19873 5859 19907
rect 5859 19873 5868 19907
rect 5816 19864 5868 19873
rect 6000 19932 6052 19984
rect 6184 19932 6236 19984
rect 8300 19932 8352 19984
rect 8484 19864 8536 19916
rect 5080 19796 5132 19848
rect 5264 19839 5316 19848
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 7748 19796 7800 19848
rect 9220 19864 9272 19916
rect 10324 19864 10376 19916
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 14096 19864 14148 19916
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 4712 19728 4764 19780
rect 5908 19728 5960 19780
rect 9772 19728 9824 19780
rect 10600 19796 10652 19848
rect 11336 19839 11388 19848
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 12992 19796 13044 19848
rect 13268 19796 13320 19848
rect 13820 19796 13872 19848
rect 14188 19796 14240 19848
rect 13728 19728 13780 19780
rect 14648 19796 14700 19848
rect 15384 20000 15436 20052
rect 16764 20000 16816 20052
rect 17316 20000 17368 20052
rect 17960 20043 18012 20052
rect 17960 20009 17969 20043
rect 17969 20009 18003 20043
rect 18003 20009 18012 20043
rect 17960 20000 18012 20009
rect 18788 20000 18840 20052
rect 19248 20000 19300 20052
rect 19984 20000 20036 20052
rect 18972 19932 19024 19984
rect 20996 20000 21048 20052
rect 21364 20000 21416 20052
rect 22284 20000 22336 20052
rect 22560 20000 22612 20052
rect 17132 19864 17184 19916
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17500 19796 17552 19805
rect 19156 19864 19208 19916
rect 19892 19864 19944 19916
rect 17960 19796 18012 19848
rect 2228 19660 2280 19712
rect 2412 19660 2464 19712
rect 2872 19660 2924 19712
rect 3148 19660 3200 19712
rect 4804 19660 4856 19712
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 5540 19660 5592 19712
rect 5816 19660 5868 19712
rect 6092 19660 6144 19712
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 9864 19660 9916 19712
rect 10140 19660 10192 19712
rect 14556 19660 14608 19712
rect 15568 19728 15620 19780
rect 16028 19728 16080 19780
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 18512 19796 18564 19848
rect 18696 19796 18748 19848
rect 19340 19796 19392 19848
rect 19064 19728 19116 19780
rect 19984 19728 20036 19780
rect 22928 19839 22980 19848
rect 22928 19805 22946 19839
rect 22946 19805 22980 19839
rect 22928 19796 22980 19805
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 24952 19796 25004 19848
rect 25964 19796 26016 19848
rect 26332 19796 26384 19848
rect 16120 19660 16172 19712
rect 17316 19660 17368 19712
rect 17776 19660 17828 19712
rect 18328 19660 18380 19712
rect 19248 19660 19300 19712
rect 20628 19771 20680 19780
rect 20628 19737 20662 19771
rect 20662 19737 20680 19771
rect 20628 19728 20680 19737
rect 20996 19728 21048 19780
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 25412 19728 25464 19780
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 2044 19456 2096 19508
rect 2504 19456 2556 19508
rect 5264 19456 5316 19508
rect 6828 19456 6880 19508
rect 8392 19456 8444 19508
rect 9312 19456 9364 19508
rect 9680 19499 9732 19508
rect 9680 19465 9682 19499
rect 9682 19465 9716 19499
rect 9716 19465 9732 19499
rect 9680 19456 9732 19465
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 11060 19456 11112 19508
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 14740 19456 14792 19508
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3148 19320 3200 19372
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 4160 19363 4212 19372
rect 4160 19329 4169 19363
rect 4169 19329 4203 19363
rect 4203 19329 4212 19363
rect 4160 19320 4212 19329
rect 4436 19363 4488 19372
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 6736 19388 6788 19440
rect 2780 19184 2832 19236
rect 5080 19363 5132 19372
rect 5080 19329 5125 19363
rect 5125 19329 5132 19363
rect 5080 19320 5132 19329
rect 5540 19320 5592 19372
rect 5172 19184 5224 19236
rect 6552 19320 6604 19372
rect 8944 19388 8996 19440
rect 7748 19320 7800 19372
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 7656 19252 7708 19304
rect 9036 19320 9088 19372
rect 10968 19431 11020 19440
rect 10968 19397 10977 19431
rect 10977 19397 11011 19431
rect 11011 19397 11020 19431
rect 10968 19388 11020 19397
rect 11428 19388 11480 19440
rect 15200 19388 15252 19440
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 6460 19184 6512 19236
rect 9588 19184 9640 19236
rect 2688 19116 2740 19168
rect 2872 19116 2924 19168
rect 3976 19116 4028 19168
rect 4896 19116 4948 19168
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10416 19252 10468 19304
rect 11244 19320 11296 19372
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12992 19320 13044 19372
rect 13728 19320 13780 19372
rect 13820 19320 13872 19372
rect 11796 19184 11848 19236
rect 14648 19252 14700 19304
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 10968 19116 11020 19168
rect 11244 19116 11296 19168
rect 12348 19116 12400 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 12716 19116 12768 19168
rect 13360 19116 13412 19168
rect 14280 19116 14332 19168
rect 15476 19320 15528 19372
rect 17500 19499 17552 19508
rect 17500 19465 17509 19499
rect 17509 19465 17543 19499
rect 17543 19465 17552 19499
rect 17500 19456 17552 19465
rect 18604 19499 18656 19508
rect 18604 19465 18613 19499
rect 18613 19465 18647 19499
rect 18647 19465 18656 19499
rect 18604 19456 18656 19465
rect 18696 19456 18748 19508
rect 19524 19456 19576 19508
rect 16028 19431 16080 19440
rect 16028 19397 16037 19431
rect 16037 19397 16071 19431
rect 16071 19397 16080 19431
rect 16028 19388 16080 19397
rect 17776 19388 17828 19440
rect 17960 19388 18012 19440
rect 18144 19388 18196 19440
rect 18236 19431 18288 19440
rect 18236 19397 18245 19431
rect 18245 19397 18279 19431
rect 18279 19397 18288 19431
rect 18236 19388 18288 19397
rect 19248 19388 19300 19440
rect 19616 19388 19668 19440
rect 19984 19456 20036 19508
rect 23572 19456 23624 19508
rect 20444 19388 20496 19440
rect 24492 19388 24544 19440
rect 15384 19252 15436 19304
rect 15292 19184 15344 19236
rect 16672 19252 16724 19304
rect 16304 19184 16356 19236
rect 15108 19116 15160 19168
rect 19340 19252 19392 19304
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 18512 19116 18564 19168
rect 18788 19184 18840 19236
rect 19892 19184 19944 19236
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 25412 19499 25464 19508
rect 25412 19465 25421 19499
rect 25421 19465 25455 19499
rect 25455 19465 25464 19499
rect 25412 19456 25464 19465
rect 20260 19252 20312 19304
rect 21640 19252 21692 19304
rect 25872 19320 25924 19372
rect 24492 19252 24544 19304
rect 20628 19184 20680 19236
rect 20996 19184 21048 19236
rect 21732 19184 21784 19236
rect 23940 19116 23992 19168
rect 24584 19159 24636 19168
rect 24584 19125 24593 19159
rect 24593 19125 24627 19159
rect 24627 19125 24636 19159
rect 24584 19116 24636 19125
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 1676 18912 1728 18964
rect 2688 18912 2740 18964
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 4160 18844 4212 18896
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 2412 18776 2464 18828
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 3056 18708 3108 18760
rect 3884 18708 3936 18760
rect 6184 18708 6236 18760
rect 7288 18912 7340 18964
rect 9588 18912 9640 18964
rect 11796 18955 11848 18964
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 9312 18844 9364 18896
rect 13360 18912 13412 18964
rect 16304 18912 16356 18964
rect 12532 18887 12584 18896
rect 12532 18853 12541 18887
rect 12541 18853 12575 18887
rect 12575 18853 12584 18887
rect 12532 18844 12584 18853
rect 19156 18912 19208 18964
rect 19248 18955 19300 18964
rect 19248 18921 19257 18955
rect 19257 18921 19291 18955
rect 19291 18921 19300 18955
rect 19248 18912 19300 18921
rect 19616 18912 19668 18964
rect 20168 18955 20220 18964
rect 20168 18921 20177 18955
rect 20177 18921 20211 18955
rect 20211 18921 20220 18955
rect 20168 18912 20220 18921
rect 22376 18955 22428 18964
rect 22376 18921 22385 18955
rect 22385 18921 22419 18955
rect 22419 18921 22428 18955
rect 22376 18912 22428 18921
rect 23756 18955 23808 18964
rect 23756 18921 23765 18955
rect 23765 18921 23799 18955
rect 23799 18921 23808 18955
rect 23756 18912 23808 18921
rect 23940 18912 23992 18964
rect 24584 18912 24636 18964
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 20444 18844 20496 18896
rect 10048 18776 10100 18828
rect 7012 18708 7064 18760
rect 3516 18572 3568 18624
rect 3608 18572 3660 18624
rect 6736 18640 6788 18692
rect 7748 18708 7800 18760
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 9956 18708 10008 18760
rect 10048 18640 10100 18692
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 10968 18776 11020 18828
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 13820 18776 13872 18828
rect 11152 18640 11204 18692
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13728 18708 13780 18760
rect 14004 18708 14056 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 14188 18708 14240 18760
rect 13176 18683 13228 18692
rect 13176 18649 13185 18683
rect 13185 18649 13219 18683
rect 13219 18649 13228 18683
rect 14740 18708 14792 18760
rect 15476 18708 15528 18760
rect 15660 18708 15712 18760
rect 17960 18776 18012 18828
rect 19432 18819 19484 18828
rect 19432 18785 19450 18819
rect 19450 18785 19484 18819
rect 19432 18776 19484 18785
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 20812 18776 20864 18828
rect 20996 18776 21048 18828
rect 17408 18708 17460 18760
rect 13176 18640 13228 18649
rect 15384 18683 15436 18692
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 18880 18640 18932 18692
rect 19156 18640 19208 18692
rect 19800 18640 19852 18692
rect 20168 18683 20220 18692
rect 10416 18572 10468 18624
rect 12992 18572 13044 18624
rect 13544 18572 13596 18624
rect 13912 18572 13964 18624
rect 14648 18572 14700 18624
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 16028 18572 16080 18624
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 16764 18572 16816 18624
rect 17040 18572 17092 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 18144 18572 18196 18624
rect 19064 18572 19116 18624
rect 19524 18615 19576 18624
rect 19524 18581 19533 18615
rect 19533 18581 19567 18615
rect 19567 18581 19576 18615
rect 19524 18572 19576 18581
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 19616 18572 19668 18581
rect 19892 18572 19944 18624
rect 20168 18649 20195 18683
rect 20195 18649 20220 18683
rect 20168 18640 20220 18649
rect 20536 18708 20588 18760
rect 20996 18572 21048 18624
rect 21732 18844 21784 18896
rect 22284 18776 22336 18828
rect 22836 18776 22888 18828
rect 23572 18887 23624 18896
rect 23572 18853 23581 18887
rect 23581 18853 23615 18887
rect 23615 18853 23624 18887
rect 23572 18844 23624 18853
rect 25688 18776 25740 18828
rect 25964 18819 26016 18828
rect 25964 18785 25973 18819
rect 25973 18785 26007 18819
rect 26007 18785 26016 18819
rect 25964 18776 26016 18785
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 23664 18708 23716 18760
rect 26240 18751 26292 18760
rect 21824 18615 21876 18624
rect 21824 18581 21833 18615
rect 21833 18581 21867 18615
rect 21867 18581 21876 18615
rect 21824 18572 21876 18581
rect 21916 18572 21968 18624
rect 23480 18640 23532 18692
rect 24124 18640 24176 18692
rect 24216 18683 24268 18692
rect 24216 18649 24225 18683
rect 24225 18649 24259 18683
rect 24259 18649 24268 18683
rect 24216 18640 24268 18649
rect 26240 18717 26274 18751
rect 26274 18717 26292 18751
rect 26240 18708 26292 18717
rect 26700 18640 26752 18692
rect 22284 18572 22336 18624
rect 22744 18572 22796 18624
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 24032 18615 24084 18624
rect 24032 18581 24059 18615
rect 24059 18581 24084 18615
rect 24032 18572 24084 18581
rect 25964 18572 26016 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 2320 18411 2372 18420
rect 2320 18377 2329 18411
rect 2329 18377 2363 18411
rect 2363 18377 2372 18411
rect 2320 18368 2372 18377
rect 3240 18368 3292 18420
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 4804 18368 4856 18420
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 2596 18300 2648 18352
rect 1768 18232 1820 18284
rect 2320 18232 2372 18284
rect 2504 18275 2556 18284
rect 2504 18241 2513 18275
rect 2513 18241 2547 18275
rect 2547 18241 2556 18275
rect 2504 18232 2556 18241
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 4436 18300 4488 18352
rect 5448 18300 5500 18352
rect 4344 18275 4396 18284
rect 2688 18096 2740 18148
rect 3332 18096 3384 18148
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 5264 18232 5316 18284
rect 6920 18368 6972 18420
rect 9312 18368 9364 18420
rect 9496 18368 9548 18420
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 5908 18275 5960 18284
rect 5908 18241 5917 18275
rect 5917 18241 5951 18275
rect 5951 18241 5960 18275
rect 5908 18232 5960 18241
rect 6736 18232 6788 18284
rect 7748 18232 7800 18284
rect 6000 18164 6052 18216
rect 6184 18207 6236 18216
rect 6184 18173 6193 18207
rect 6193 18173 6227 18207
rect 6227 18173 6236 18207
rect 6184 18164 6236 18173
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 4804 18096 4856 18148
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 9128 18275 9180 18284
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 9496 18275 9548 18284
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 9680 18368 9732 18420
rect 11244 18368 11296 18420
rect 12164 18368 12216 18420
rect 12992 18368 13044 18420
rect 9956 18300 10008 18352
rect 10048 18232 10100 18284
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 11980 18232 12032 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 13912 18232 13964 18284
rect 14188 18232 14240 18284
rect 16764 18368 16816 18420
rect 17408 18368 17460 18420
rect 22560 18411 22612 18420
rect 22560 18377 22569 18411
rect 22569 18377 22603 18411
rect 22603 18377 22612 18411
rect 22560 18368 22612 18377
rect 14648 18343 14700 18352
rect 14648 18309 14657 18343
rect 14657 18309 14691 18343
rect 14691 18309 14700 18343
rect 14648 18300 14700 18309
rect 15108 18232 15160 18284
rect 15200 18232 15252 18284
rect 15936 18300 15988 18352
rect 15752 18232 15804 18284
rect 14832 18207 14884 18216
rect 14832 18173 14841 18207
rect 14841 18173 14875 18207
rect 14875 18173 14884 18207
rect 14832 18164 14884 18173
rect 15476 18164 15528 18216
rect 16028 18164 16080 18216
rect 17132 18343 17184 18352
rect 16304 18164 16356 18216
rect 4252 18028 4304 18080
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 8576 18028 8628 18037
rect 9680 18028 9732 18080
rect 13176 18096 13228 18148
rect 13452 18028 13504 18080
rect 15384 18096 15436 18148
rect 17132 18309 17155 18343
rect 17155 18309 17184 18343
rect 17132 18300 17184 18309
rect 17316 18300 17368 18352
rect 14740 18028 14792 18080
rect 15292 18028 15344 18080
rect 15660 18028 15712 18080
rect 15936 18028 15988 18080
rect 16764 18028 16816 18080
rect 16948 18232 17000 18284
rect 17960 18232 18012 18284
rect 18696 18300 18748 18352
rect 20904 18343 20956 18352
rect 19248 18232 19300 18284
rect 20904 18309 20931 18343
rect 20931 18309 20956 18343
rect 20904 18300 20956 18309
rect 20996 18300 21048 18352
rect 22376 18343 22428 18352
rect 22376 18309 22385 18343
rect 22385 18309 22419 18343
rect 22419 18309 22428 18343
rect 22376 18300 22428 18309
rect 25964 18411 26016 18420
rect 25964 18377 25973 18411
rect 25973 18377 26007 18411
rect 26007 18377 26016 18411
rect 25964 18368 26016 18377
rect 18236 18164 18288 18216
rect 19064 18164 19116 18216
rect 21916 18164 21968 18216
rect 20536 18096 20588 18148
rect 21456 18096 21508 18148
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 22376 18164 22428 18216
rect 22928 18164 22980 18216
rect 23204 18232 23256 18284
rect 23848 18232 23900 18284
rect 24308 18275 24360 18284
rect 24308 18241 24317 18275
rect 24317 18241 24351 18275
rect 24351 18241 24360 18275
rect 24308 18232 24360 18241
rect 24584 18207 24636 18216
rect 24584 18173 24593 18207
rect 24593 18173 24627 18207
rect 24627 18173 24636 18207
rect 24584 18164 24636 18173
rect 17776 18028 17828 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 19524 18028 19576 18080
rect 21364 18028 21416 18080
rect 22468 18028 22520 18080
rect 22928 18071 22980 18080
rect 22928 18037 22937 18071
rect 22937 18037 22971 18071
rect 22971 18037 22980 18071
rect 22928 18028 22980 18037
rect 26700 18275 26752 18284
rect 26700 18241 26709 18275
rect 26709 18241 26743 18275
rect 26743 18241 26752 18275
rect 26700 18232 26752 18241
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 26516 18028 26568 18080
rect 26884 18028 26936 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 1768 17824 1820 17876
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 3792 17824 3844 17876
rect 4804 17824 4856 17876
rect 10324 17824 10376 17876
rect 10784 17824 10836 17876
rect 5908 17756 5960 17808
rect 7656 17756 7708 17808
rect 8576 17799 8628 17808
rect 8576 17765 8585 17799
rect 8585 17765 8619 17799
rect 8619 17765 8628 17799
rect 8576 17756 8628 17765
rect 9404 17756 9456 17808
rect 4160 17688 4212 17740
rect 1676 17595 1728 17604
rect 1676 17561 1685 17595
rect 1685 17561 1719 17595
rect 1719 17561 1728 17595
rect 1676 17552 1728 17561
rect 2504 17552 2556 17604
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 3332 17663 3384 17672
rect 3332 17629 3341 17663
rect 3341 17629 3375 17663
rect 3375 17629 3384 17663
rect 3332 17620 3384 17629
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 4252 17620 4304 17672
rect 5172 17688 5224 17740
rect 8852 17688 8904 17740
rect 9680 17756 9732 17808
rect 4896 17663 4948 17672
rect 4896 17629 4905 17663
rect 4905 17629 4939 17663
rect 4939 17629 4948 17663
rect 4896 17620 4948 17629
rect 5264 17620 5316 17672
rect 1584 17484 1636 17536
rect 6368 17552 6420 17604
rect 7104 17620 7156 17672
rect 8576 17620 8628 17672
rect 5080 17484 5132 17536
rect 5632 17484 5684 17536
rect 9404 17620 9456 17672
rect 10508 17620 10560 17672
rect 12624 17824 12676 17876
rect 13820 17824 13872 17876
rect 15844 17824 15896 17876
rect 16580 17824 16632 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 16856 17824 16908 17876
rect 19349 17824 19401 17876
rect 11704 17756 11756 17808
rect 13176 17756 13228 17808
rect 14280 17756 14332 17808
rect 22284 17824 22336 17876
rect 23572 17756 23624 17808
rect 23940 17799 23992 17808
rect 23940 17765 23949 17799
rect 23949 17765 23983 17799
rect 23983 17765 23992 17799
rect 23940 17756 23992 17765
rect 13268 17688 13320 17740
rect 12164 17595 12216 17604
rect 12164 17561 12198 17595
rect 12198 17561 12216 17595
rect 12164 17552 12216 17561
rect 14556 17688 14608 17740
rect 16304 17688 16356 17740
rect 13176 17552 13228 17604
rect 14740 17620 14792 17672
rect 16212 17620 16264 17672
rect 14004 17552 14056 17604
rect 9956 17484 10008 17536
rect 11796 17484 11848 17536
rect 13084 17484 13136 17536
rect 15384 17552 15436 17604
rect 19892 17688 19944 17740
rect 23112 17688 23164 17740
rect 24308 17824 24360 17876
rect 25136 17824 25188 17876
rect 26516 17756 26568 17808
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 16948 17552 17000 17604
rect 19524 17620 19576 17672
rect 19616 17595 19668 17604
rect 19616 17561 19625 17595
rect 19625 17561 19659 17595
rect 19659 17561 19668 17595
rect 19616 17552 19668 17561
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20996 17620 21048 17672
rect 20628 17552 20680 17604
rect 23204 17663 23256 17672
rect 23204 17629 23208 17663
rect 23208 17629 23242 17663
rect 23242 17629 23256 17663
rect 23204 17620 23256 17629
rect 23388 17595 23440 17604
rect 23388 17561 23397 17595
rect 23397 17561 23431 17595
rect 23431 17561 23440 17595
rect 23388 17552 23440 17561
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 25136 17620 25188 17672
rect 26884 17663 26936 17672
rect 24768 17595 24820 17604
rect 24768 17561 24777 17595
rect 24777 17561 24811 17595
rect 24811 17561 24820 17595
rect 24768 17552 24820 17561
rect 14832 17484 14884 17536
rect 16304 17527 16356 17536
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 16580 17484 16632 17536
rect 20260 17484 20312 17536
rect 21364 17484 21416 17536
rect 24584 17484 24636 17536
rect 26884 17629 26893 17663
rect 26893 17629 26927 17663
rect 26927 17629 26936 17663
rect 26884 17620 26936 17629
rect 26976 17620 27028 17672
rect 25504 17595 25556 17604
rect 25504 17561 25538 17595
rect 25538 17561 25556 17595
rect 25504 17552 25556 17561
rect 26240 17552 26292 17604
rect 26700 17595 26752 17604
rect 26700 17561 26709 17595
rect 26709 17561 26743 17595
rect 26743 17561 26752 17595
rect 26700 17552 26752 17561
rect 27436 17595 27488 17604
rect 27436 17561 27470 17595
rect 27470 17561 27488 17595
rect 27436 17552 27488 17561
rect 27068 17527 27120 17536
rect 27068 17493 27077 17527
rect 27077 17493 27111 17527
rect 27111 17493 27120 17527
rect 27068 17484 27120 17493
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 1676 17212 1728 17264
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 3884 17280 3936 17332
rect 5356 17280 5408 17332
rect 5540 17280 5592 17332
rect 12072 17280 12124 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 6092 17212 6144 17264
rect 7748 17212 7800 17264
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 1768 16940 1820 16992
rect 4896 17076 4948 17128
rect 6920 17144 6972 17196
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 8668 17144 8720 17196
rect 11704 17212 11756 17264
rect 12256 17144 12308 17196
rect 12532 17144 12584 17196
rect 14280 17280 14332 17332
rect 14648 17280 14700 17332
rect 15200 17280 15252 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 21088 17280 21140 17332
rect 21548 17280 21600 17332
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13360 17144 13412 17196
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 14096 17212 14148 17264
rect 23204 17323 23256 17332
rect 23204 17289 23213 17323
rect 23213 17289 23247 17323
rect 23247 17289 23256 17323
rect 23204 17280 23256 17289
rect 23572 17280 23624 17332
rect 23940 17280 23992 17332
rect 24676 17280 24728 17332
rect 25504 17323 25556 17332
rect 25504 17289 25513 17323
rect 25513 17289 25547 17323
rect 25547 17289 25556 17323
rect 25504 17280 25556 17289
rect 27436 17323 27488 17332
rect 27436 17289 27445 17323
rect 27445 17289 27479 17323
rect 27479 17289 27488 17323
rect 27436 17280 27488 17289
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 5908 17051 5960 17060
rect 5908 17017 5917 17051
rect 5917 17017 5951 17051
rect 5951 17017 5960 17051
rect 5908 17008 5960 17017
rect 6000 17008 6052 17060
rect 9128 17008 9180 17060
rect 17776 17144 17828 17196
rect 17960 17144 18012 17196
rect 18604 17144 18656 17196
rect 18788 17187 18840 17196
rect 18788 17153 18822 17187
rect 18822 17153 18840 17187
rect 18788 17144 18840 17153
rect 20260 17187 20312 17196
rect 20260 17153 20283 17187
rect 20283 17153 20312 17187
rect 20260 17144 20312 17153
rect 21548 17144 21600 17196
rect 22100 17144 22152 17196
rect 24032 17144 24084 17196
rect 26240 17212 26292 17264
rect 25596 17144 25648 17196
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9956 16940 10008 16992
rect 10876 16940 10928 16992
rect 12256 16940 12308 16992
rect 15752 16940 15804 16992
rect 18696 16940 18748 16992
rect 19432 16940 19484 16992
rect 19892 16983 19944 16992
rect 19892 16949 19901 16983
rect 19901 16949 19935 16983
rect 19935 16949 19944 16983
rect 19892 16940 19944 16949
rect 20996 17008 21048 17060
rect 22468 17076 22520 17128
rect 23112 17076 23164 17128
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 6000 16736 6052 16788
rect 9128 16736 9180 16788
rect 9864 16736 9916 16788
rect 11980 16736 12032 16788
rect 9404 16711 9456 16720
rect 9404 16677 9413 16711
rect 9413 16677 9447 16711
rect 9447 16677 9456 16711
rect 9404 16668 9456 16677
rect 10232 16668 10284 16720
rect 3516 16576 3568 16584
rect 3516 16542 3534 16576
rect 3534 16542 3568 16576
rect 3516 16532 3568 16542
rect 2044 16464 2096 16516
rect 4160 16532 4212 16584
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 4896 16532 4948 16584
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 5172 16532 5224 16584
rect 3792 16396 3844 16448
rect 3976 16396 4028 16448
rect 4804 16396 4856 16448
rect 7380 16575 7432 16584
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 7656 16507 7708 16516
rect 7656 16473 7690 16507
rect 7690 16473 7708 16507
rect 7656 16464 7708 16473
rect 8760 16464 8812 16516
rect 10784 16600 10836 16652
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 12072 16668 12124 16720
rect 12532 16736 12584 16788
rect 16856 16779 16908 16788
rect 16856 16745 16865 16779
rect 16865 16745 16899 16779
rect 16899 16745 16908 16779
rect 16856 16736 16908 16745
rect 18052 16736 18104 16788
rect 18788 16779 18840 16788
rect 18788 16745 18797 16779
rect 18797 16745 18831 16779
rect 18831 16745 18840 16779
rect 18788 16736 18840 16745
rect 14188 16668 14240 16720
rect 14648 16668 14700 16720
rect 10968 16507 11020 16516
rect 10968 16473 10977 16507
rect 10977 16473 11011 16507
rect 11011 16473 11020 16507
rect 10968 16464 11020 16473
rect 6184 16396 6236 16448
rect 6736 16396 6788 16448
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 12256 16643 12308 16652
rect 12256 16609 12265 16643
rect 12265 16609 12299 16643
rect 12299 16609 12308 16643
rect 12256 16600 12308 16609
rect 18328 16668 18380 16720
rect 18880 16668 18932 16720
rect 12716 16532 12768 16584
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16580 16532 16632 16541
rect 16672 16532 16724 16584
rect 18236 16532 18288 16584
rect 18972 16600 19024 16652
rect 19156 16600 19208 16652
rect 19524 16600 19576 16652
rect 19984 16736 20036 16788
rect 21088 16736 21140 16788
rect 22468 16736 22520 16788
rect 23204 16736 23256 16788
rect 23388 16736 23440 16788
rect 23756 16736 23808 16788
rect 25596 16736 25648 16788
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 18696 16532 18748 16584
rect 19432 16532 19484 16584
rect 12808 16507 12860 16516
rect 12808 16473 12817 16507
rect 12817 16473 12851 16507
rect 12851 16473 12860 16507
rect 12808 16464 12860 16473
rect 11980 16396 12032 16448
rect 12440 16396 12492 16448
rect 13268 16464 13320 16516
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 14280 16396 14332 16448
rect 14556 16396 14608 16448
rect 16856 16507 16908 16516
rect 16856 16473 16865 16507
rect 16865 16473 16899 16507
rect 16899 16473 16908 16507
rect 16856 16464 16908 16473
rect 17500 16464 17552 16516
rect 17960 16464 18012 16516
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 19892 16532 19944 16541
rect 21088 16575 21140 16584
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 17224 16396 17276 16448
rect 17776 16396 17828 16448
rect 18420 16396 18472 16448
rect 19708 16507 19760 16516
rect 19708 16473 19717 16507
rect 19717 16473 19751 16507
rect 19751 16473 19760 16507
rect 19708 16464 19760 16473
rect 19800 16464 19852 16516
rect 20260 16464 20312 16516
rect 19432 16439 19484 16448
rect 19432 16405 19459 16439
rect 19459 16405 19484 16439
rect 19432 16396 19484 16405
rect 19524 16396 19576 16448
rect 20536 16439 20588 16448
rect 20536 16405 20558 16439
rect 20558 16405 20588 16439
rect 22100 16532 22152 16584
rect 23848 16711 23900 16720
rect 23848 16677 23857 16711
rect 23857 16677 23891 16711
rect 23891 16677 23900 16711
rect 23848 16668 23900 16677
rect 25136 16711 25188 16720
rect 25136 16677 25145 16711
rect 25145 16677 25179 16711
rect 25179 16677 25188 16711
rect 25136 16668 25188 16677
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 24584 16600 24636 16652
rect 20536 16396 20588 16405
rect 23572 16507 23624 16516
rect 23572 16473 23581 16507
rect 23581 16473 23615 16507
rect 23615 16473 23624 16507
rect 23572 16464 23624 16473
rect 23848 16464 23900 16516
rect 24860 16507 24912 16516
rect 24860 16473 24869 16507
rect 24869 16473 24903 16507
rect 24903 16473 24912 16507
rect 24860 16464 24912 16473
rect 27068 16532 27120 16584
rect 26424 16464 26476 16516
rect 27160 16396 27212 16448
rect 27528 16439 27580 16448
rect 27528 16405 27537 16439
rect 27537 16405 27571 16439
rect 27571 16405 27580 16439
rect 27528 16396 27580 16405
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 2872 16192 2924 16244
rect 3792 16192 3844 16244
rect 4068 16192 4120 16244
rect 1676 16167 1728 16176
rect 1676 16133 1685 16167
rect 1685 16133 1719 16167
rect 1719 16133 1728 16167
rect 1676 16124 1728 16133
rect 2964 16124 3016 16176
rect 756 16056 808 16108
rect 3332 16056 3384 16108
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 4896 16124 4948 16176
rect 5816 16192 5868 16244
rect 6184 16192 6236 16244
rect 7196 16192 7248 16244
rect 7656 16192 7708 16244
rect 9404 16192 9456 16244
rect 10968 16235 11020 16244
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 7104 16056 7156 16108
rect 8668 16124 8720 16176
rect 12072 16192 12124 16244
rect 12716 16192 12768 16244
rect 9864 16099 9916 16108
rect 9864 16065 9898 16099
rect 9898 16065 9916 16099
rect 3148 15988 3200 16040
rect 3976 15988 4028 16040
rect 9864 16056 9916 16065
rect 14004 16192 14056 16244
rect 14188 16192 14240 16244
rect 14740 16192 14792 16244
rect 15936 16192 15988 16244
rect 16120 16192 16172 16244
rect 17040 16235 17092 16244
rect 14280 16124 14332 16176
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 12164 16056 12216 16108
rect 12808 16056 12860 16108
rect 13176 16056 13228 16108
rect 15108 16056 15160 16108
rect 16120 16056 16172 16108
rect 5264 15920 5316 15972
rect 6092 15963 6144 15972
rect 6092 15929 6101 15963
rect 6101 15929 6135 15963
rect 6135 15929 6144 15963
rect 6092 15920 6144 15929
rect 6736 15963 6788 15972
rect 6736 15929 6745 15963
rect 6745 15929 6779 15963
rect 6779 15929 6788 15963
rect 6736 15920 6788 15929
rect 7380 15920 7432 15972
rect 2136 15852 2188 15904
rect 4344 15852 4396 15904
rect 14648 15988 14700 16040
rect 15476 15988 15528 16040
rect 16304 16056 16356 16108
rect 16396 16099 16448 16108
rect 16396 16065 16405 16099
rect 16405 16065 16439 16099
rect 16439 16065 16448 16099
rect 16396 16056 16448 16065
rect 19708 16192 19760 16244
rect 20352 16192 20404 16244
rect 20628 16192 20680 16244
rect 21088 16192 21140 16244
rect 21364 16192 21416 16244
rect 21640 16192 21692 16244
rect 18328 16124 18380 16176
rect 22836 16192 22888 16244
rect 22376 16124 22428 16176
rect 24768 16192 24820 16244
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 18512 16056 18564 16108
rect 19524 15988 19576 16040
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 20444 16056 20496 16108
rect 20996 16056 21048 16108
rect 24308 16056 24360 16108
rect 25688 16124 25740 16176
rect 26148 16192 26200 16244
rect 26424 16235 26476 16244
rect 26424 16201 26433 16235
rect 26433 16201 26467 16235
rect 26467 16201 26476 16235
rect 26424 16192 26476 16201
rect 27528 16192 27580 16244
rect 24584 16056 24636 16108
rect 24768 16099 24820 16108
rect 24768 16065 24802 16099
rect 24802 16065 24820 16099
rect 24768 16056 24820 16065
rect 26976 16056 27028 16108
rect 11244 15852 11296 15904
rect 13084 15852 13136 15904
rect 15016 15895 15068 15904
rect 15016 15861 15025 15895
rect 15025 15861 15059 15895
rect 15059 15861 15068 15895
rect 15016 15852 15068 15861
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 15568 15852 15620 15904
rect 17408 15852 17460 15904
rect 20720 15852 20772 15904
rect 21088 15852 21140 15904
rect 21824 15895 21876 15904
rect 21824 15861 21833 15895
rect 21833 15861 21867 15895
rect 21867 15861 21876 15895
rect 21824 15852 21876 15861
rect 23204 15920 23256 15972
rect 24124 15920 24176 15972
rect 23112 15852 23164 15904
rect 25872 15895 25924 15904
rect 25872 15861 25881 15895
rect 25881 15861 25915 15895
rect 25915 15861 25924 15895
rect 25872 15852 25924 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 3332 15648 3384 15700
rect 4344 15648 4396 15700
rect 4804 15648 4856 15700
rect 9496 15648 9548 15700
rect 9864 15648 9916 15700
rect 10508 15648 10560 15700
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 12716 15648 12768 15700
rect 13636 15648 13688 15700
rect 14372 15648 14424 15700
rect 4160 15580 4212 15632
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 3240 15444 3292 15496
rect 3792 15444 3844 15496
rect 5724 15512 5776 15564
rect 6000 15512 6052 15564
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 9312 15512 9364 15564
rect 3976 15376 4028 15428
rect 4160 15419 4212 15428
rect 4160 15385 4169 15419
rect 4169 15385 4203 15419
rect 4203 15385 4212 15419
rect 4160 15376 4212 15385
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 15936 15648 15988 15700
rect 17040 15648 17092 15700
rect 13084 15623 13136 15632
rect 13084 15589 13093 15623
rect 13093 15589 13127 15623
rect 13127 15589 13136 15623
rect 13084 15580 13136 15589
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 12900 15512 12952 15564
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 14280 15444 14332 15496
rect 15016 15580 15068 15632
rect 15108 15623 15160 15632
rect 15108 15589 15117 15623
rect 15117 15589 15151 15623
rect 15151 15589 15160 15623
rect 15108 15580 15160 15589
rect 16120 15580 16172 15632
rect 14924 15444 14976 15496
rect 15292 15460 15344 15512
rect 11152 15376 11204 15428
rect 1676 15308 1728 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 5724 15308 5776 15360
rect 7380 15308 7432 15360
rect 8300 15308 8352 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 9312 15308 9364 15360
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 13820 15419 13872 15428
rect 13820 15385 13829 15419
rect 13829 15385 13863 15419
rect 13863 15385 13872 15419
rect 13820 15376 13872 15385
rect 14556 15419 14608 15428
rect 14556 15385 14565 15419
rect 14565 15385 14599 15419
rect 14599 15385 14608 15419
rect 14556 15376 14608 15385
rect 16304 15512 16356 15564
rect 16948 15444 17000 15496
rect 17592 15691 17644 15700
rect 17592 15657 17601 15691
rect 17601 15657 17635 15691
rect 17635 15657 17644 15691
rect 17592 15648 17644 15657
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 21824 15648 21876 15700
rect 23112 15691 23164 15700
rect 23112 15657 23121 15691
rect 23121 15657 23155 15691
rect 23155 15657 23164 15691
rect 23112 15648 23164 15657
rect 15936 15419 15988 15428
rect 15936 15385 15945 15419
rect 15945 15385 15979 15419
rect 15979 15385 15988 15419
rect 15936 15376 15988 15385
rect 17224 15376 17276 15428
rect 17592 15376 17644 15428
rect 18052 15580 18104 15632
rect 20536 15580 20588 15632
rect 23756 15623 23808 15632
rect 23756 15589 23765 15623
rect 23765 15589 23799 15623
rect 23799 15589 23808 15623
rect 23756 15580 23808 15589
rect 24308 15648 24360 15700
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 25688 15648 25740 15700
rect 25136 15580 25188 15632
rect 25872 15580 25924 15632
rect 18236 15512 18288 15564
rect 19064 15444 19116 15496
rect 19156 15444 19208 15496
rect 20628 15444 20680 15496
rect 18328 15419 18380 15428
rect 18328 15385 18337 15419
rect 18337 15385 18371 15419
rect 18371 15385 18380 15419
rect 18328 15376 18380 15385
rect 21088 15444 21140 15496
rect 21272 15444 21324 15496
rect 24768 15444 24820 15496
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 28448 15487 28500 15496
rect 28448 15453 28457 15487
rect 28457 15453 28491 15487
rect 28491 15453 28500 15487
rect 28448 15444 28500 15453
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16120 15308 16172 15360
rect 16948 15308 17000 15360
rect 17408 15308 17460 15360
rect 18604 15308 18656 15360
rect 20996 15376 21048 15428
rect 22192 15376 22244 15428
rect 22928 15376 22980 15428
rect 24032 15376 24084 15428
rect 24124 15419 24176 15428
rect 24124 15385 24133 15419
rect 24133 15385 24167 15419
rect 24167 15385 24176 15419
rect 24124 15376 24176 15385
rect 27436 15376 27488 15428
rect 20352 15308 20404 15360
rect 20444 15308 20496 15360
rect 21640 15308 21692 15360
rect 22560 15308 22612 15360
rect 22836 15308 22888 15360
rect 23388 15308 23440 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 1676 15079 1728 15088
rect 1676 15045 1710 15079
rect 1710 15045 1728 15079
rect 5448 15104 5500 15156
rect 5632 15104 5684 15156
rect 6000 15104 6052 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8300 15104 8352 15156
rect 1676 15036 1728 15045
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 4344 14968 4396 15020
rect 4620 15011 4672 15020
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 4804 15036 4856 15088
rect 9404 15104 9456 15156
rect 11152 15147 11204 15156
rect 11152 15113 11161 15147
rect 11161 15113 11195 15147
rect 11195 15113 11204 15147
rect 11152 15104 11204 15113
rect 11244 15104 11296 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 12900 15104 12952 15156
rect 14556 15104 14608 15156
rect 15752 15104 15804 15156
rect 3516 14900 3568 14952
rect 6092 14968 6144 15020
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 11704 14968 11756 15020
rect 13820 15036 13872 15088
rect 7104 14900 7156 14952
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 11152 14900 11204 14952
rect 14004 14968 14056 15020
rect 17776 15104 17828 15156
rect 18052 15147 18104 15156
rect 18052 15113 18061 15147
rect 18061 15113 18095 15147
rect 18095 15113 18104 15147
rect 18052 15104 18104 15113
rect 18328 15104 18380 15156
rect 20260 15036 20312 15088
rect 21732 15104 21784 15156
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 27436 15147 27488 15156
rect 27436 15113 27445 15147
rect 27445 15113 27479 15147
rect 27479 15113 27488 15147
rect 27436 15104 27488 15113
rect 17316 14968 17368 15020
rect 2136 14764 2188 14816
rect 2688 14764 2740 14816
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 9312 14764 9364 14816
rect 11980 14832 12032 14884
rect 15752 14832 15804 14884
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 16580 14764 16632 14816
rect 21640 15036 21692 15088
rect 21364 14968 21416 15020
rect 22560 14968 22612 15020
rect 23756 15011 23808 15020
rect 23756 14977 23790 15011
rect 23790 14977 23808 15011
rect 23756 14968 23808 14977
rect 24860 15036 24912 15088
rect 17868 14900 17920 14952
rect 20260 14900 20312 14952
rect 20812 14900 20864 14952
rect 21640 14900 21692 14952
rect 25596 14943 25648 14952
rect 25596 14909 25605 14943
rect 25605 14909 25639 14943
rect 25639 14909 25648 14943
rect 25596 14900 25648 14909
rect 17684 14832 17736 14884
rect 17776 14832 17828 14884
rect 20628 14832 20680 14884
rect 20996 14832 21048 14884
rect 21456 14832 21508 14884
rect 25688 14832 25740 14884
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 26976 14832 27028 14884
rect 19156 14764 19208 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 20720 14807 20772 14816
rect 20720 14773 20729 14807
rect 20729 14773 20763 14807
rect 20763 14773 20772 14807
rect 20720 14764 20772 14773
rect 21272 14764 21324 14816
rect 23480 14764 23532 14816
rect 24860 14807 24912 14816
rect 24860 14773 24869 14807
rect 24869 14773 24903 14807
rect 24903 14773 24912 14807
rect 24860 14764 24912 14773
rect 26332 14807 26384 14816
rect 26332 14773 26341 14807
rect 26341 14773 26375 14807
rect 26375 14773 26384 14807
rect 26332 14764 26384 14773
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 2504 14560 2556 14612
rect 3148 14560 3200 14612
rect 3332 14560 3384 14612
rect 4344 14560 4396 14612
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 13544 14560 13596 14612
rect 15476 14560 15528 14612
rect 17316 14560 17368 14612
rect 18052 14560 18104 14612
rect 19708 14560 19760 14612
rect 20168 14560 20220 14612
rect 3424 14424 3476 14476
rect 4252 14492 4304 14544
rect 4988 14492 5040 14544
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2872 14356 2924 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 8116 14424 8168 14476
rect 14372 14424 14424 14476
rect 3056 14288 3108 14340
rect 2688 14220 2740 14272
rect 2964 14220 3016 14272
rect 4896 14288 4948 14340
rect 5172 14356 5224 14408
rect 5724 14356 5776 14408
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 7380 14399 7432 14408
rect 7380 14365 7414 14399
rect 7414 14365 7432 14399
rect 7380 14356 7432 14365
rect 9220 14399 9272 14408
rect 9220 14365 9254 14399
rect 9254 14365 9272 14399
rect 9220 14356 9272 14365
rect 9772 14356 9824 14408
rect 10876 14399 10928 14408
rect 10876 14365 10910 14399
rect 10910 14365 10928 14399
rect 10876 14356 10928 14365
rect 12808 14356 12860 14408
rect 12992 14288 13044 14340
rect 14188 14288 14240 14340
rect 14372 14288 14424 14340
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 10324 14263 10376 14272
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 11704 14220 11756 14272
rect 13176 14220 13228 14272
rect 13820 14220 13872 14272
rect 14464 14220 14516 14272
rect 17592 14492 17644 14544
rect 16396 14424 16448 14476
rect 17684 14424 17736 14476
rect 17868 14424 17920 14476
rect 19524 14424 19576 14476
rect 22192 14560 22244 14612
rect 23756 14560 23808 14612
rect 27252 14560 27304 14612
rect 23480 14535 23532 14544
rect 23480 14501 23489 14535
rect 23489 14501 23523 14535
rect 23523 14501 23532 14535
rect 23480 14492 23532 14501
rect 19340 14356 19392 14408
rect 15200 14220 15252 14272
rect 17316 14220 17368 14272
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 17776 14220 17828 14272
rect 18328 14263 18380 14272
rect 18328 14229 18337 14263
rect 18337 14229 18371 14263
rect 18371 14229 18380 14263
rect 18328 14220 18380 14229
rect 20168 14356 20220 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 27528 14535 27580 14544
rect 27528 14501 27537 14535
rect 27537 14501 27571 14535
rect 27571 14501 27580 14535
rect 27528 14492 27580 14501
rect 24952 14424 25004 14476
rect 23848 14356 23900 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 20352 14288 20404 14340
rect 20904 14288 20956 14340
rect 26332 14356 26384 14408
rect 26976 14356 27028 14408
rect 27344 14288 27396 14340
rect 20168 14263 20220 14272
rect 20168 14229 20177 14263
rect 20177 14229 20211 14263
rect 20211 14229 20220 14263
rect 20168 14220 20220 14229
rect 20628 14263 20680 14272
rect 20628 14229 20637 14263
rect 20637 14229 20671 14263
rect 20671 14229 20680 14263
rect 20628 14220 20680 14229
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 25596 14220 25648 14272
rect 25688 14263 25740 14272
rect 25688 14229 25697 14263
rect 25697 14229 25731 14263
rect 25731 14229 25740 14263
rect 25688 14220 25740 14229
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 3424 14016 3476 14068
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 4252 14016 4304 14068
rect 4988 14016 5040 14068
rect 10692 14016 10744 14068
rect 12532 14016 12584 14068
rect 2688 13991 2740 14000
rect 2688 13957 2697 13991
rect 2697 13957 2731 13991
rect 2731 13957 2740 13991
rect 2688 13948 2740 13957
rect 2872 13991 2924 14000
rect 2872 13957 2881 13991
rect 2881 13957 2915 13991
rect 2915 13957 2924 13991
rect 2872 13948 2924 13957
rect 6276 13948 6328 14000
rect 8760 13948 8812 14000
rect 756 13880 808 13932
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 3976 13676 4028 13728
rect 4988 13812 5040 13864
rect 6460 13812 6512 13864
rect 11152 13948 11204 14000
rect 9680 13880 9732 13932
rect 10324 13880 10376 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 13544 13880 13596 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 13820 13880 13872 13932
rect 14188 13948 14240 14000
rect 15936 14016 15988 14068
rect 17776 14016 17828 14068
rect 17960 14016 18012 14068
rect 18328 14016 18380 14068
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 20444 14059 20496 14068
rect 20444 14025 20453 14059
rect 20453 14025 20487 14059
rect 20487 14025 20496 14059
rect 20444 14016 20496 14025
rect 20628 14016 20680 14068
rect 20904 14016 20956 14068
rect 21456 14016 21508 14068
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14832 13880 14884 13932
rect 15016 13923 15068 13932
rect 15016 13889 15050 13923
rect 15050 13889 15068 13923
rect 15016 13880 15068 13889
rect 15476 13880 15528 13932
rect 16396 13880 16448 13932
rect 17592 13880 17644 13932
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 18236 13880 18288 13889
rect 19984 13948 20036 14000
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 22376 14016 22428 14068
rect 24952 14016 25004 14068
rect 20904 13880 20956 13932
rect 21364 13880 21416 13932
rect 6092 13676 6144 13728
rect 7748 13676 7800 13728
rect 8300 13676 8352 13728
rect 9220 13787 9272 13796
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 9220 13744 9272 13753
rect 9772 13744 9824 13796
rect 13452 13787 13504 13796
rect 13452 13753 13461 13787
rect 13461 13753 13495 13787
rect 13495 13753 13504 13787
rect 13452 13744 13504 13753
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 17040 13812 17092 13864
rect 18052 13812 18104 13864
rect 19524 13812 19576 13864
rect 20352 13812 20404 13864
rect 20444 13812 20496 13864
rect 22008 13812 22060 13864
rect 28448 13948 28500 14000
rect 23756 13923 23808 13932
rect 23756 13889 23765 13923
rect 23765 13889 23799 13923
rect 23799 13889 23808 13923
rect 23756 13880 23808 13889
rect 26976 13880 27028 13932
rect 28264 13923 28316 13932
rect 28264 13889 28282 13923
rect 28282 13889 28316 13923
rect 28264 13880 28316 13889
rect 22836 13812 22888 13864
rect 25596 13812 25648 13864
rect 16948 13787 17000 13796
rect 16948 13753 16957 13787
rect 16957 13753 16991 13787
rect 16991 13753 17000 13787
rect 16948 13744 17000 13753
rect 14464 13676 14516 13728
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 17224 13744 17276 13796
rect 17316 13744 17368 13796
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 18972 13676 19024 13728
rect 19248 13676 19300 13728
rect 19800 13719 19852 13728
rect 19800 13685 19809 13719
rect 19809 13685 19843 13719
rect 19843 13685 19852 13719
rect 19800 13676 19852 13685
rect 22376 13719 22428 13728
rect 22376 13685 22385 13719
rect 22385 13685 22419 13719
rect 22419 13685 22428 13719
rect 22376 13676 22428 13685
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 1400 13472 1452 13524
rect 2044 13472 2096 13524
rect 2504 13472 2556 13524
rect 3332 13472 3384 13524
rect 5448 13472 5500 13524
rect 6276 13472 6328 13524
rect 2872 13268 2924 13320
rect 3608 13200 3660 13252
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 7104 13336 7156 13388
rect 6184 13268 6236 13320
rect 2596 13175 2648 13184
rect 2596 13141 2605 13175
rect 2605 13141 2639 13175
rect 2639 13141 2648 13175
rect 2596 13132 2648 13141
rect 4436 13132 4488 13184
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9220 13472 9272 13524
rect 9680 13404 9732 13456
rect 9496 13268 9548 13320
rect 7656 13243 7708 13252
rect 7656 13209 7690 13243
rect 7690 13209 7708 13243
rect 7656 13200 7708 13209
rect 9128 13200 9180 13252
rect 11152 13404 11204 13456
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 14188 13472 14240 13524
rect 15016 13515 15068 13524
rect 15016 13481 15025 13515
rect 15025 13481 15059 13515
rect 15059 13481 15068 13515
rect 15016 13472 15068 13481
rect 15752 13472 15804 13524
rect 16672 13515 16724 13524
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 17592 13472 17644 13524
rect 19708 13472 19760 13524
rect 19800 13472 19852 13524
rect 19984 13472 20036 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20996 13472 21048 13524
rect 22008 13515 22060 13524
rect 22008 13481 22017 13515
rect 22017 13481 22051 13515
rect 22051 13481 22060 13515
rect 22008 13472 22060 13481
rect 23756 13472 23808 13524
rect 26976 13472 27028 13524
rect 14464 13404 14516 13456
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 11060 13268 11112 13320
rect 11152 13268 11204 13320
rect 11428 13311 11480 13320
rect 11428 13277 11438 13311
rect 11438 13277 11472 13311
rect 11472 13277 11480 13311
rect 11428 13268 11480 13277
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 12532 13311 12584 13320
rect 9772 13200 9824 13252
rect 11244 13200 11296 13252
rect 10048 13132 10100 13184
rect 10416 13132 10468 13184
rect 11060 13132 11112 13184
rect 11336 13132 11388 13184
rect 12532 13277 12555 13311
rect 12555 13277 12584 13311
rect 12532 13268 12584 13277
rect 13268 13268 13320 13320
rect 14372 13268 14424 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 14832 13200 14884 13252
rect 17500 13336 17552 13388
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 19984 13336 20036 13388
rect 17684 13268 17736 13320
rect 17960 13268 18012 13320
rect 18144 13268 18196 13320
rect 12348 13132 12400 13184
rect 14648 13132 14700 13184
rect 17500 13243 17552 13252
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 18972 13311 19024 13320
rect 18972 13277 18981 13311
rect 18981 13277 19015 13311
rect 19015 13277 19024 13311
rect 18972 13268 19024 13277
rect 19524 13268 19576 13320
rect 19156 13200 19208 13252
rect 19432 13243 19484 13252
rect 19432 13209 19441 13243
rect 19441 13209 19475 13243
rect 19475 13209 19484 13243
rect 19432 13200 19484 13209
rect 19708 13243 19760 13252
rect 19708 13209 19717 13243
rect 19717 13209 19751 13243
rect 19751 13209 19760 13243
rect 19708 13200 19760 13209
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 22100 13404 22152 13456
rect 23940 13447 23992 13456
rect 23940 13413 23949 13447
rect 23949 13413 23983 13447
rect 23983 13413 23992 13447
rect 23940 13404 23992 13413
rect 28264 13472 28316 13524
rect 27620 13447 27672 13456
rect 27620 13413 27629 13447
rect 27629 13413 27663 13447
rect 27663 13413 27672 13447
rect 27620 13404 27672 13413
rect 27344 13379 27396 13388
rect 27344 13345 27353 13379
rect 27353 13345 27387 13379
rect 27387 13345 27396 13379
rect 27344 13336 27396 13345
rect 20076 13243 20128 13252
rect 20076 13209 20085 13243
rect 20085 13209 20119 13243
rect 20119 13209 20128 13243
rect 20076 13200 20128 13209
rect 16580 13132 16632 13184
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 17316 13175 17368 13184
rect 17316 13141 17343 13175
rect 17343 13141 17368 13175
rect 17316 13132 17368 13141
rect 17408 13132 17460 13184
rect 17684 13132 17736 13184
rect 21364 13200 21416 13252
rect 22376 13243 22428 13252
rect 22376 13209 22410 13243
rect 22410 13209 22428 13243
rect 22376 13200 22428 13209
rect 24952 13268 25004 13320
rect 23020 13132 23072 13184
rect 23388 13132 23440 13184
rect 24400 13175 24452 13184
rect 24400 13141 24409 13175
rect 24409 13141 24443 13175
rect 24443 13141 24452 13175
rect 24400 13132 24452 13141
rect 25964 13200 26016 13252
rect 26240 13200 26292 13252
rect 24952 13132 25004 13184
rect 25136 13132 25188 13184
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 2872 12928 2924 12980
rect 2136 12860 2188 12912
rect 4436 12928 4488 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 7656 12928 7708 12980
rect 7748 12928 7800 12980
rect 1676 12835 1728 12844
rect 1676 12801 1710 12835
rect 1710 12801 1728 12835
rect 1676 12792 1728 12801
rect 3332 12792 3384 12844
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 6644 12903 6696 12912
rect 4160 12792 4212 12844
rect 6644 12869 6667 12903
rect 6667 12869 6696 12903
rect 6644 12860 6696 12869
rect 6276 12792 6328 12844
rect 6092 12724 6144 12776
rect 6368 12767 6420 12776
rect 6368 12733 6377 12767
rect 6377 12733 6411 12767
rect 6411 12733 6420 12767
rect 6368 12724 6420 12733
rect 4988 12699 5040 12708
rect 4988 12665 4997 12699
rect 4997 12665 5031 12699
rect 5031 12665 5040 12699
rect 4988 12656 5040 12665
rect 9312 12928 9364 12980
rect 9404 12928 9456 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 10968 12928 11020 12980
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 4344 12588 4396 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 8300 12588 8352 12640
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 14648 12928 14700 12980
rect 12256 12860 12308 12912
rect 11428 12792 11480 12844
rect 11796 12792 11848 12844
rect 12808 12792 12860 12844
rect 9496 12724 9548 12776
rect 11336 12724 11388 12776
rect 11244 12656 11296 12708
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13084 12792 13136 12844
rect 13820 12792 13872 12844
rect 17316 12928 17368 12980
rect 9220 12588 9272 12640
rect 10876 12588 10928 12640
rect 12440 12656 12492 12708
rect 12164 12588 12216 12640
rect 14740 12656 14792 12708
rect 15936 12792 15988 12844
rect 16488 12792 16540 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17684 12860 17736 12912
rect 17592 12835 17644 12844
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 16488 12699 16540 12708
rect 16488 12665 16497 12699
rect 16497 12665 16531 12699
rect 16531 12665 16540 12699
rect 16488 12656 16540 12665
rect 16580 12656 16632 12708
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 17132 12656 17184 12708
rect 17316 12656 17368 12708
rect 19432 12928 19484 12980
rect 19984 12928 20036 12980
rect 20076 12928 20128 12980
rect 21364 12928 21416 12980
rect 25044 12928 25096 12980
rect 25596 12928 25648 12980
rect 20444 12860 20496 12912
rect 21640 12860 21692 12912
rect 17960 12792 18012 12844
rect 19156 12792 19208 12844
rect 20076 12724 20128 12776
rect 20996 12835 21048 12844
rect 20996 12801 21008 12835
rect 21008 12801 21042 12835
rect 21042 12801 21048 12835
rect 20996 12792 21048 12801
rect 21180 12792 21232 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 20536 12699 20588 12708
rect 20536 12665 20545 12699
rect 20545 12665 20579 12699
rect 20579 12665 20588 12699
rect 20536 12656 20588 12665
rect 22284 12835 22336 12844
rect 22284 12801 22319 12835
rect 22319 12801 22336 12835
rect 23020 12903 23072 12912
rect 23020 12869 23029 12903
rect 23029 12869 23063 12903
rect 23063 12869 23072 12903
rect 23020 12860 23072 12869
rect 25136 12860 25188 12912
rect 26148 12928 26200 12980
rect 26240 12971 26292 12980
rect 26240 12937 26249 12971
rect 26249 12937 26283 12971
rect 26283 12937 26292 12971
rect 26240 12928 26292 12937
rect 27620 12928 27672 12980
rect 22284 12792 22336 12801
rect 20720 12588 20772 12640
rect 21272 12631 21324 12640
rect 21272 12597 21281 12631
rect 21281 12597 21315 12631
rect 21315 12597 21324 12631
rect 21272 12588 21324 12597
rect 21640 12588 21692 12640
rect 23848 12792 23900 12844
rect 24952 12792 25004 12844
rect 22192 12656 22244 12708
rect 23020 12724 23072 12776
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 23940 12724 23992 12776
rect 23388 12699 23440 12708
rect 23388 12665 23397 12699
rect 23397 12665 23431 12699
rect 23431 12665 23440 12699
rect 23388 12656 23440 12665
rect 23572 12656 23624 12708
rect 26976 12792 27028 12844
rect 27436 12835 27488 12844
rect 27436 12801 27470 12835
rect 27470 12801 27488 12835
rect 27436 12792 27488 12801
rect 24400 12588 24452 12640
rect 25228 12631 25280 12640
rect 25228 12597 25237 12631
rect 25237 12597 25271 12631
rect 25271 12597 25280 12631
rect 25228 12588 25280 12597
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 1676 12384 1728 12436
rect 1768 12316 1820 12368
rect 756 12180 808 12232
rect 3332 12384 3384 12436
rect 13084 12384 13136 12436
rect 14372 12384 14424 12436
rect 15844 12384 15896 12436
rect 17040 12384 17092 12436
rect 17592 12384 17644 12436
rect 18236 12427 18288 12436
rect 18236 12393 18245 12427
rect 18245 12393 18279 12427
rect 18279 12393 18288 12427
rect 18236 12384 18288 12393
rect 18880 12384 18932 12436
rect 19708 12384 19760 12436
rect 16488 12316 16540 12368
rect 21364 12384 21416 12436
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 27436 12384 27488 12436
rect 19984 12359 20036 12368
rect 19984 12325 19993 12359
rect 19993 12325 20027 12359
rect 20027 12325 20036 12359
rect 19984 12316 20036 12325
rect 20812 12316 20864 12368
rect 20996 12316 21048 12368
rect 22560 12316 22612 12368
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 7380 12248 7432 12300
rect 11980 12248 12032 12300
rect 2228 12180 2280 12232
rect 2596 12180 2648 12232
rect 3240 12180 3292 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 13820 12248 13872 12300
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 15292 12248 15344 12300
rect 2044 12044 2096 12096
rect 14648 12112 14700 12164
rect 9588 12044 9640 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 15108 12112 15160 12164
rect 15476 12180 15528 12232
rect 17408 12248 17460 12300
rect 16028 12044 16080 12096
rect 17316 12180 17368 12232
rect 17776 12112 17828 12164
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 19616 12248 19668 12300
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 19156 12180 19208 12232
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 19984 12180 20036 12232
rect 21456 12248 21508 12300
rect 17500 12044 17552 12096
rect 19248 12112 19300 12164
rect 20168 12112 20220 12164
rect 21180 12180 21232 12232
rect 23480 12180 23532 12232
rect 25044 12223 25096 12232
rect 25044 12189 25053 12223
rect 25053 12189 25087 12223
rect 25087 12189 25096 12223
rect 25044 12180 25096 12189
rect 26700 12223 26752 12232
rect 26700 12189 26709 12223
rect 26709 12189 26743 12223
rect 26743 12189 26752 12223
rect 26700 12180 26752 12189
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 20444 12044 20496 12096
rect 20904 12044 20956 12096
rect 22192 12044 22244 12096
rect 25412 12044 25464 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 3516 11840 3568 11892
rect 4160 11840 4212 11892
rect 6092 11840 6144 11892
rect 3608 11772 3660 11824
rect 2964 11704 3016 11756
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 7380 11772 7432 11824
rect 10048 11840 10100 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 14188 11840 14240 11892
rect 18604 11840 18656 11892
rect 19248 11883 19300 11892
rect 19248 11849 19273 11883
rect 19273 11849 19300 11883
rect 19248 11840 19300 11849
rect 19892 11840 19944 11892
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 2596 11636 2648 11688
rect 2136 11568 2188 11620
rect 8668 11568 8720 11620
rect 9036 11611 9088 11620
rect 9036 11577 9045 11611
rect 9045 11577 9079 11611
rect 9079 11577 9088 11611
rect 9036 11568 9088 11577
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 5724 11500 5776 11552
rect 6828 11500 6880 11552
rect 7656 11500 7708 11552
rect 11796 11772 11848 11824
rect 15292 11772 15344 11824
rect 16120 11772 16172 11824
rect 16304 11772 16356 11824
rect 11888 11704 11940 11756
rect 12164 11704 12216 11756
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 14372 11636 14424 11688
rect 17132 11636 17184 11688
rect 19248 11704 19300 11756
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 20352 11704 20404 11756
rect 21088 11747 21140 11756
rect 21088 11713 21098 11747
rect 21098 11713 21132 11747
rect 21132 11713 21140 11747
rect 21088 11704 21140 11713
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 19984 11636 20036 11688
rect 20904 11636 20956 11688
rect 21916 11840 21968 11892
rect 22468 11840 22520 11892
rect 22008 11772 22060 11824
rect 23020 11815 23072 11824
rect 23020 11781 23055 11815
rect 23055 11781 23072 11815
rect 23020 11772 23072 11781
rect 24952 11772 25004 11824
rect 21640 11704 21692 11756
rect 21916 11747 21968 11756
rect 21916 11713 21926 11747
rect 21926 11713 21960 11747
rect 21960 11713 21968 11747
rect 21916 11704 21968 11713
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 11704 11568 11756 11620
rect 13820 11568 13872 11620
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 18788 11500 18840 11552
rect 20352 11543 20404 11552
rect 20352 11509 20361 11543
rect 20361 11509 20395 11543
rect 20395 11509 20404 11543
rect 20352 11500 20404 11509
rect 21640 11611 21692 11620
rect 21640 11577 21649 11611
rect 21649 11577 21683 11611
rect 21683 11577 21692 11611
rect 21640 11568 21692 11577
rect 22100 11568 22152 11620
rect 22376 11568 22428 11620
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 23388 11704 23440 11756
rect 27436 11747 27488 11756
rect 27436 11713 27470 11747
rect 27470 11713 27488 11747
rect 27436 11704 27488 11713
rect 26240 11636 26292 11688
rect 26700 11636 26752 11688
rect 25412 11568 25464 11620
rect 21364 11500 21416 11552
rect 21548 11500 21600 11552
rect 23664 11500 23716 11552
rect 23940 11500 23992 11552
rect 25596 11543 25648 11552
rect 25596 11509 25605 11543
rect 25605 11509 25639 11543
rect 25639 11509 25648 11543
rect 25596 11500 25648 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 2504 11296 2556 11348
rect 5632 11296 5684 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 9772 11296 9824 11348
rect 10140 11296 10192 11348
rect 10692 11296 10744 11348
rect 12532 11296 12584 11348
rect 5172 11271 5224 11280
rect 5172 11237 5181 11271
rect 5181 11237 5215 11271
rect 5215 11237 5224 11271
rect 5172 11228 5224 11237
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 5724 11135 5776 11144
rect 5724 11101 5758 11135
rect 5758 11101 5776 11135
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 3148 11024 3200 11033
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 5724 11092 5776 11101
rect 6460 11092 6512 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7656 11135 7708 11144
rect 7656 11101 7690 11135
rect 7690 11101 7708 11135
rect 7656 11092 7708 11101
rect 8852 11092 8904 11144
rect 9680 11228 9732 11280
rect 11336 11228 11388 11280
rect 13728 11228 13780 11280
rect 14464 11296 14516 11348
rect 9312 11160 9364 11212
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 10600 11160 10652 11212
rect 9588 11092 9640 11144
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14188 11160 14240 11212
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 12992 11092 13044 11144
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 9680 10956 9732 11008
rect 13820 11024 13872 11076
rect 14372 11024 14424 11076
rect 14648 11160 14700 11212
rect 17960 11160 18012 11212
rect 20352 11228 20404 11280
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 10508 10956 10560 11008
rect 11980 10956 12032 11008
rect 14556 10999 14608 11008
rect 14556 10965 14565 10999
rect 14565 10965 14599 10999
rect 14599 10965 14608 10999
rect 14556 10956 14608 10965
rect 16028 11024 16080 11076
rect 16764 11092 16816 11144
rect 17500 11092 17552 11144
rect 16212 11067 16264 11076
rect 16212 11033 16246 11067
rect 16246 11033 16264 11067
rect 16212 11024 16264 11033
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 21364 11092 21416 11144
rect 23664 11228 23716 11280
rect 27344 11339 27396 11348
rect 27344 11305 27353 11339
rect 27353 11305 27387 11339
rect 27387 11305 27396 11339
rect 27344 11296 27396 11305
rect 27436 11339 27488 11348
rect 27436 11305 27445 11339
rect 27445 11305 27479 11339
rect 27479 11305 27488 11339
rect 27436 11296 27488 11305
rect 23204 11160 23256 11212
rect 23848 11160 23900 11212
rect 22560 11092 22612 11144
rect 23296 11135 23348 11144
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 24860 11160 24912 11212
rect 15752 10956 15804 11008
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 16948 10956 17000 11008
rect 17684 10956 17736 11008
rect 17776 10956 17828 11008
rect 19248 10956 19300 11008
rect 20536 10956 20588 11008
rect 21916 11024 21968 11076
rect 23480 11024 23532 11076
rect 24216 11135 24268 11144
rect 24216 11101 24225 11135
rect 24225 11101 24259 11135
rect 24259 11101 24268 11135
rect 24216 11092 24268 11101
rect 25596 11092 25648 11144
rect 26240 11092 26292 11144
rect 27436 11092 27488 11144
rect 24400 11024 24452 11076
rect 26884 11067 26936 11076
rect 26884 11033 26893 11067
rect 26893 11033 26927 11067
rect 26927 11033 26936 11067
rect 26884 11024 26936 11033
rect 21088 10956 21140 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 1952 10752 2004 10804
rect 1860 10684 1912 10736
rect 756 10616 808 10668
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 3976 10684 4028 10736
rect 5080 10684 5132 10736
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 7104 10684 7156 10736
rect 8852 10727 8904 10736
rect 8852 10693 8869 10727
rect 8869 10693 8904 10727
rect 8852 10684 8904 10693
rect 9036 10752 9088 10804
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6460 10616 6512 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 9588 10752 9640 10804
rect 9956 10752 10008 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 10784 10752 10836 10804
rect 11888 10752 11940 10804
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 12808 10752 12860 10804
rect 9496 10684 9548 10736
rect 11336 10684 11388 10736
rect 16028 10752 16080 10804
rect 16212 10795 16264 10804
rect 16212 10761 16221 10795
rect 16221 10761 16255 10795
rect 16255 10761 16264 10795
rect 16212 10752 16264 10761
rect 16856 10752 16908 10804
rect 17960 10752 18012 10804
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 19984 10752 20036 10804
rect 20168 10752 20220 10804
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 7748 10480 7800 10532
rect 10232 10659 10284 10668
rect 10232 10625 10241 10659
rect 10241 10625 10275 10659
rect 10275 10625 10284 10659
rect 10232 10616 10284 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 11244 10616 11296 10668
rect 11704 10659 11756 10668
rect 11704 10625 11711 10659
rect 11711 10625 11756 10659
rect 11704 10616 11756 10625
rect 15200 10684 15252 10736
rect 16948 10684 17000 10736
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 5172 10412 5224 10464
rect 5632 10412 5684 10464
rect 9312 10548 9364 10600
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 12348 10616 12400 10668
rect 12992 10616 13044 10668
rect 13176 10616 13228 10668
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 13544 10616 13596 10668
rect 13636 10616 13688 10668
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 15844 10616 15896 10668
rect 16304 10616 16356 10668
rect 17592 10616 17644 10668
rect 11888 10480 11940 10532
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 17132 10548 17184 10600
rect 15752 10480 15804 10532
rect 19064 10684 19116 10736
rect 19616 10684 19668 10736
rect 20536 10684 20588 10736
rect 22652 10752 22704 10804
rect 23388 10752 23440 10804
rect 23848 10752 23900 10804
rect 27436 10795 27488 10804
rect 27436 10761 27445 10795
rect 27445 10761 27479 10795
rect 27479 10761 27488 10795
rect 27436 10752 27488 10761
rect 21088 10727 21140 10736
rect 21088 10693 21097 10727
rect 21097 10693 21131 10727
rect 21131 10693 21140 10727
rect 21088 10684 21140 10693
rect 21272 10684 21324 10736
rect 23112 10684 23164 10736
rect 24676 10684 24728 10736
rect 24952 10684 25004 10736
rect 26884 10684 26936 10736
rect 18236 10616 18288 10668
rect 23020 10616 23072 10668
rect 23480 10659 23532 10668
rect 23480 10625 23484 10659
rect 23484 10625 23518 10659
rect 23518 10625 23532 10659
rect 23480 10616 23532 10625
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 23756 10659 23808 10668
rect 23756 10625 23801 10659
rect 23801 10625 23808 10659
rect 23756 10616 23808 10625
rect 18328 10548 18380 10600
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 23020 10480 23072 10532
rect 23388 10548 23440 10600
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 24032 10480 24084 10532
rect 24492 10480 24544 10532
rect 25688 10523 25740 10532
rect 25688 10489 25697 10523
rect 25697 10489 25731 10523
rect 25731 10489 25740 10523
rect 25688 10480 25740 10489
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 22192 10412 22244 10464
rect 22468 10455 22520 10464
rect 22468 10421 22477 10455
rect 22477 10421 22511 10455
rect 22511 10421 22520 10455
rect 22468 10412 22520 10421
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 23940 10412 23992 10464
rect 25872 10455 25924 10464
rect 25872 10421 25881 10455
rect 25881 10421 25915 10455
rect 25915 10421 25924 10455
rect 25872 10412 25924 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1584 10208 1636 10260
rect 1860 10140 1912 10192
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 2688 10072 2740 10124
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 5264 10208 5316 10260
rect 6184 10208 6236 10260
rect 7288 10208 7340 10260
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 9312 10208 9364 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 5632 10183 5684 10192
rect 5632 10149 5641 10183
rect 5641 10149 5675 10183
rect 5675 10149 5684 10183
rect 5632 10140 5684 10149
rect 5816 10183 5868 10192
rect 5816 10149 5825 10183
rect 5825 10149 5859 10183
rect 5859 10149 5868 10183
rect 5816 10140 5868 10149
rect 7656 10140 7708 10192
rect 5172 10072 5224 10124
rect 2780 9936 2832 9988
rect 4896 9936 4948 9988
rect 5724 10004 5776 10056
rect 8760 10004 8812 10056
rect 3056 9868 3108 9920
rect 7380 9936 7432 9988
rect 9036 9979 9088 9988
rect 9036 9945 9045 9979
rect 9045 9945 9079 9979
rect 9079 9945 9088 9979
rect 9036 9936 9088 9945
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 11244 10208 11296 10260
rect 12992 10208 13044 10260
rect 14280 10208 14332 10260
rect 15384 10208 15436 10260
rect 15568 10208 15620 10260
rect 15844 10208 15896 10260
rect 18236 10208 18288 10260
rect 20352 10208 20404 10260
rect 20628 10251 20680 10260
rect 20628 10217 20637 10251
rect 20637 10217 20671 10251
rect 20671 10217 20680 10251
rect 20628 10208 20680 10217
rect 22192 10251 22244 10260
rect 22192 10217 22201 10251
rect 22201 10217 22235 10251
rect 22235 10217 22244 10251
rect 22192 10208 22244 10217
rect 23204 10208 23256 10260
rect 23664 10208 23716 10260
rect 23848 10208 23900 10260
rect 24216 10208 24268 10260
rect 11980 10183 12032 10192
rect 11980 10149 11989 10183
rect 11989 10149 12023 10183
rect 12023 10149 12032 10183
rect 11980 10140 12032 10149
rect 14464 10183 14516 10192
rect 14464 10149 14473 10183
rect 14473 10149 14507 10183
rect 14507 10149 14516 10183
rect 14464 10140 14516 10149
rect 16580 10072 16632 10124
rect 17776 10072 17828 10124
rect 23756 10140 23808 10192
rect 24952 10140 25004 10192
rect 26240 10208 26292 10260
rect 13360 10004 13412 10056
rect 9588 9936 9640 9988
rect 10968 9936 11020 9988
rect 12072 9936 12124 9988
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 16120 10004 16172 10056
rect 17132 10004 17184 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 17684 9936 17736 9988
rect 19340 9936 19392 9988
rect 19616 9979 19668 9988
rect 19616 9945 19625 9979
rect 19625 9945 19659 9979
rect 19659 9945 19668 9979
rect 19616 9936 19668 9945
rect 19892 9936 19944 9988
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 16948 9868 17000 9920
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 20444 9911 20496 9920
rect 20444 9877 20469 9911
rect 20469 9877 20496 9911
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 21180 9936 21232 9988
rect 22652 9936 22704 9988
rect 20444 9868 20496 9877
rect 21640 9868 21692 9920
rect 22192 9868 22244 9920
rect 22376 9911 22428 9920
rect 22376 9877 22393 9911
rect 22393 9877 22428 9911
rect 22376 9868 22428 9877
rect 22836 9868 22888 9920
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23940 10004 23992 10056
rect 24492 10072 24544 10124
rect 24032 9868 24084 9920
rect 25872 10047 25924 10056
rect 25872 10013 25906 10047
rect 25906 10013 25924 10047
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 24584 9868 24636 9920
rect 25872 10004 25924 10013
rect 27528 9936 27580 9988
rect 27252 9868 27304 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 1860 9664 1912 9716
rect 10876 9664 10928 9716
rect 14464 9664 14516 9716
rect 1492 9596 1544 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 2044 9596 2096 9648
rect 5816 9596 5868 9648
rect 8760 9596 8812 9648
rect 2136 9528 2188 9580
rect 2688 9528 2740 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 2504 9392 2556 9444
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 2136 9324 2188 9376
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3608 9324 3660 9376
rect 3792 9392 3844 9444
rect 5908 9528 5960 9580
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7748 9528 7800 9580
rect 9864 9528 9916 9580
rect 13176 9596 13228 9648
rect 13452 9596 13504 9648
rect 16120 9664 16172 9716
rect 6092 9460 6144 9512
rect 10600 9528 10652 9580
rect 11244 9528 11296 9580
rect 6644 9392 6696 9444
rect 12532 9528 12584 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 12900 9528 12952 9580
rect 14188 9528 14240 9580
rect 14464 9528 14516 9580
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 14648 9460 14700 9512
rect 15292 9639 15344 9648
rect 15292 9605 15319 9639
rect 15319 9605 15344 9639
rect 15292 9596 15344 9605
rect 16580 9664 16632 9716
rect 17224 9664 17276 9716
rect 17960 9664 18012 9716
rect 20352 9664 20404 9716
rect 20720 9664 20772 9716
rect 21180 9707 21232 9716
rect 21180 9673 21189 9707
rect 21189 9673 21223 9707
rect 21223 9673 21232 9707
rect 21180 9664 21232 9673
rect 21272 9664 21324 9716
rect 22468 9664 22520 9716
rect 22928 9664 22980 9716
rect 24768 9664 24820 9716
rect 27528 9707 27580 9716
rect 27528 9673 27537 9707
rect 27537 9673 27571 9707
rect 27571 9673 27580 9707
rect 27528 9664 27580 9673
rect 17040 9596 17092 9648
rect 17776 9596 17828 9648
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16212 9460 16264 9512
rect 11980 9392 12032 9444
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7932 9367 7984 9376
rect 7932 9333 7941 9367
rect 7941 9333 7975 9367
rect 7975 9333 7984 9367
rect 7932 9324 7984 9333
rect 9588 9324 9640 9376
rect 9680 9324 9732 9376
rect 10692 9324 10744 9376
rect 10968 9324 11020 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 14188 9324 14240 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 14556 9324 14608 9376
rect 16028 9324 16080 9376
rect 18972 9528 19024 9580
rect 19524 9528 19576 9580
rect 21732 9596 21784 9648
rect 22008 9639 22060 9648
rect 22008 9605 22033 9639
rect 22033 9605 22060 9639
rect 22008 9596 22060 9605
rect 22376 9596 22428 9648
rect 24124 9596 24176 9648
rect 26884 9596 26936 9648
rect 22652 9528 22704 9580
rect 21088 9392 21140 9444
rect 22836 9392 22888 9444
rect 27252 9435 27304 9444
rect 27252 9401 27261 9435
rect 27261 9401 27295 9435
rect 27295 9401 27304 9435
rect 27252 9392 27304 9401
rect 20628 9324 20680 9376
rect 21180 9324 21232 9376
rect 21456 9324 21508 9376
rect 21640 9324 21692 9376
rect 24952 9324 25004 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 1952 9120 2004 9172
rect 2596 9120 2648 9172
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2872 9120 2924 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 3700 8984 3752 9036
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 9864 9120 9916 9172
rect 10324 9120 10376 9172
rect 10232 9052 10284 9104
rect 10508 9052 10560 9104
rect 12256 9120 12308 9172
rect 12532 9052 12584 9104
rect 12900 9163 12952 9172
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 14280 9120 14332 9172
rect 14740 9120 14792 9172
rect 15200 9163 15252 9172
rect 15200 9129 15209 9163
rect 15209 9129 15243 9163
rect 15243 9129 15252 9163
rect 15200 9120 15252 9129
rect 15292 9120 15344 9172
rect 15936 9120 15988 9172
rect 16028 9120 16080 9172
rect 16212 9120 16264 9172
rect 16672 9120 16724 9172
rect 18144 9120 18196 9172
rect 18972 9163 19024 9172
rect 18972 9129 18981 9163
rect 18981 9129 19015 9163
rect 19015 9129 19024 9163
rect 18972 9120 19024 9129
rect 19524 9120 19576 9172
rect 22468 9120 22520 9172
rect 23020 9163 23072 9172
rect 23020 9129 23029 9163
rect 23029 9129 23063 9163
rect 23063 9129 23072 9163
rect 23020 9120 23072 9129
rect 14188 9052 14240 9104
rect 14556 9052 14608 9104
rect 17224 9052 17276 9104
rect 17960 9095 18012 9104
rect 17960 9061 17969 9095
rect 17969 9061 18003 9095
rect 18003 9061 18012 9095
rect 17960 9052 18012 9061
rect 9864 8984 9916 9036
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 5816 8848 5868 8900
rect 6552 8916 6604 8968
rect 7932 8916 7984 8968
rect 10600 8916 10652 8968
rect 9128 8848 9180 8900
rect 9680 8848 9732 8900
rect 9864 8848 9916 8900
rect 10692 8891 10744 8900
rect 10692 8857 10701 8891
rect 10701 8857 10735 8891
rect 10735 8857 10744 8891
rect 10692 8848 10744 8857
rect 12440 8916 12492 8968
rect 12808 8984 12860 9036
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13268 8984 13320 9036
rect 22376 9052 22428 9104
rect 23756 9163 23808 9172
rect 23756 9129 23765 9163
rect 23765 9129 23799 9163
rect 23799 9129 23808 9163
rect 23756 9120 23808 9129
rect 27620 9120 27672 9172
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 13912 8916 13964 8968
rect 5448 8780 5500 8832
rect 10508 8780 10560 8832
rect 10600 8780 10652 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11980 8780 12032 8832
rect 13084 8891 13136 8900
rect 13084 8857 13093 8891
rect 13093 8857 13127 8891
rect 13127 8857 13136 8891
rect 13084 8848 13136 8857
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 12716 8780 12768 8832
rect 13360 8780 13412 8832
rect 14740 8780 14792 8832
rect 15384 8848 15436 8900
rect 15476 8891 15528 8900
rect 15476 8857 15485 8891
rect 15485 8857 15519 8891
rect 15519 8857 15528 8891
rect 15476 8848 15528 8857
rect 17132 8916 17184 8968
rect 19248 8916 19300 8968
rect 20720 8916 20772 8968
rect 22744 8916 22796 8968
rect 23296 8916 23348 8968
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 24952 8916 25004 8968
rect 26608 8959 26660 8968
rect 26608 8925 26617 8959
rect 26617 8925 26651 8959
rect 26651 8925 26660 8959
rect 26608 8916 26660 8925
rect 15844 8780 15896 8832
rect 16120 8823 16172 8832
rect 16120 8789 16147 8823
rect 16147 8789 16172 8823
rect 16120 8780 16172 8789
rect 16580 8848 16632 8900
rect 16764 8891 16816 8900
rect 16764 8857 16773 8891
rect 16773 8857 16807 8891
rect 16807 8857 16816 8891
rect 16764 8848 16816 8857
rect 17500 8848 17552 8900
rect 17776 8848 17828 8900
rect 19616 8848 19668 8900
rect 17132 8780 17184 8832
rect 19340 8780 19392 8832
rect 21456 8848 21508 8900
rect 22652 8891 22704 8900
rect 22652 8857 22661 8891
rect 22661 8857 22695 8891
rect 22695 8857 22704 8891
rect 22652 8848 22704 8857
rect 23756 8848 23808 8900
rect 21548 8823 21600 8832
rect 21548 8789 21557 8823
rect 21557 8789 21591 8823
rect 21591 8789 21600 8823
rect 21548 8780 21600 8789
rect 21640 8780 21692 8832
rect 22836 8823 22888 8832
rect 22836 8789 22861 8823
rect 22861 8789 22888 8823
rect 22836 8780 22888 8789
rect 23940 8780 23992 8832
rect 24860 8848 24912 8900
rect 26332 8891 26384 8900
rect 26332 8857 26341 8891
rect 26341 8857 26375 8891
rect 26375 8857 26384 8891
rect 26332 8848 26384 8857
rect 25872 8823 25924 8832
rect 25872 8789 25881 8823
rect 25881 8789 25915 8823
rect 25915 8789 25924 8823
rect 25872 8780 25924 8789
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1492 8576 1544 8628
rect 2780 8576 2832 8628
rect 3148 8576 3200 8628
rect 5448 8576 5500 8628
rect 6644 8576 6696 8628
rect 6736 8576 6788 8628
rect 7748 8576 7800 8628
rect 8760 8576 8812 8628
rect 9128 8576 9180 8628
rect 9312 8576 9364 8628
rect 10232 8576 10284 8628
rect 10416 8576 10468 8628
rect 10876 8619 10928 8628
rect 10876 8585 10901 8619
rect 10901 8585 10928 8619
rect 10876 8576 10928 8585
rect 14648 8619 14700 8628
rect 14648 8585 14657 8619
rect 14657 8585 14691 8619
rect 14691 8585 14700 8619
rect 14648 8576 14700 8585
rect 14740 8576 14792 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 4160 8551 4212 8560
rect 4160 8517 4169 8551
rect 4169 8517 4203 8551
rect 4203 8517 4212 8551
rect 4160 8508 4212 8517
rect 3424 8440 3476 8492
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 5356 8304 5408 8356
rect 7564 8440 7616 8492
rect 8852 8551 8904 8560
rect 8852 8517 8886 8551
rect 8886 8517 8904 8551
rect 8852 8508 8904 8517
rect 9680 8508 9732 8560
rect 10600 8508 10652 8560
rect 10784 8508 10836 8560
rect 12072 8508 12124 8560
rect 16396 8576 16448 8628
rect 10968 8440 11020 8492
rect 11060 8440 11112 8492
rect 11704 8483 11756 8492
rect 11704 8449 11711 8483
rect 11711 8449 11756 8483
rect 11704 8440 11756 8449
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9864 8372 9916 8424
rect 11244 8372 11296 8424
rect 13452 8440 13504 8492
rect 15936 8508 15988 8560
rect 16488 8508 16540 8560
rect 16580 8508 16632 8560
rect 16948 8551 17000 8560
rect 16948 8517 16973 8551
rect 16973 8517 17000 8551
rect 17408 8576 17460 8628
rect 17592 8576 17644 8628
rect 16948 8508 17000 8517
rect 17684 8508 17736 8560
rect 13360 8372 13412 8424
rect 14648 8440 14700 8492
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 17960 8508 18012 8560
rect 19064 8508 19116 8560
rect 19984 8576 20036 8628
rect 21180 8619 21232 8628
rect 21180 8585 21205 8619
rect 21205 8585 21232 8619
rect 21180 8576 21232 8585
rect 22652 8576 22704 8628
rect 5632 8236 5684 8288
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 6828 8236 6880 8288
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 11152 8304 11204 8356
rect 12164 8347 12216 8356
rect 12164 8313 12173 8347
rect 12173 8313 12207 8347
rect 12207 8313 12216 8347
rect 12164 8304 12216 8313
rect 12256 8304 12308 8356
rect 12716 8304 12768 8356
rect 13636 8304 13688 8356
rect 16212 8372 16264 8424
rect 16396 8372 16448 8424
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20720 8440 20772 8492
rect 20996 8551 21048 8560
rect 20996 8517 21031 8551
rect 21031 8517 21048 8551
rect 20996 8508 21048 8517
rect 21548 8508 21600 8560
rect 21732 8508 21784 8560
rect 22008 8508 22060 8560
rect 20996 8372 21048 8424
rect 21640 8372 21692 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 23296 8619 23348 8628
rect 23296 8585 23305 8619
rect 23305 8585 23339 8619
rect 23339 8585 23348 8619
rect 23296 8576 23348 8585
rect 23572 8576 23624 8628
rect 23480 8551 23532 8560
rect 23480 8517 23491 8551
rect 23491 8517 23532 8551
rect 23480 8508 23532 8517
rect 23664 8551 23716 8560
rect 23664 8517 23673 8551
rect 23673 8517 23707 8551
rect 23707 8517 23716 8551
rect 23664 8508 23716 8517
rect 23848 8508 23900 8560
rect 24032 8576 24084 8628
rect 24860 8576 24912 8628
rect 25872 8576 25924 8628
rect 26608 8576 26660 8628
rect 26332 8508 26384 8560
rect 24492 8372 24544 8424
rect 10968 8236 11020 8288
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 17960 8304 18012 8356
rect 20444 8347 20496 8356
rect 20444 8313 20453 8347
rect 20453 8313 20487 8347
rect 20487 8313 20496 8347
rect 20444 8304 20496 8313
rect 15292 8236 15344 8288
rect 16028 8279 16080 8288
rect 16028 8245 16037 8279
rect 16037 8245 16071 8279
rect 16071 8245 16080 8279
rect 16028 8236 16080 8245
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 18236 8279 18288 8288
rect 18236 8245 18245 8279
rect 18245 8245 18279 8279
rect 18279 8245 18288 8279
rect 18236 8236 18288 8245
rect 19984 8279 20036 8288
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 23664 8236 23716 8288
rect 24124 8279 24176 8288
rect 24124 8245 24133 8279
rect 24133 8245 24167 8279
rect 24167 8245 24176 8279
rect 24124 8236 24176 8245
rect 24584 8347 24636 8356
rect 24584 8313 24593 8347
rect 24593 8313 24627 8347
rect 24627 8313 24636 8347
rect 24584 8304 24636 8313
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 3424 8032 3476 8084
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 3424 7828 3476 7880
rect 4804 8032 4856 8084
rect 8852 8032 8904 8084
rect 13084 8032 13136 8084
rect 14464 8032 14516 8084
rect 6644 7896 6696 7948
rect 9956 7964 10008 8016
rect 3792 7760 3844 7812
rect 1676 7692 1728 7744
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 4896 7760 4948 7812
rect 5632 7760 5684 7812
rect 6644 7760 6696 7812
rect 10232 7896 10284 7948
rect 8484 7828 8536 7880
rect 11060 7964 11112 8016
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16212 8032 16264 8084
rect 16304 8075 16356 8084
rect 16304 8041 16313 8075
rect 16313 8041 16347 8075
rect 16347 8041 16356 8075
rect 16304 8032 16356 8041
rect 17132 7964 17184 8016
rect 12532 7896 12584 7948
rect 12716 7896 12768 7948
rect 20076 8032 20128 8084
rect 21180 8032 21232 8084
rect 20720 7964 20772 8016
rect 20996 7964 21048 8016
rect 11796 7828 11848 7880
rect 12440 7828 12492 7880
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13360 7828 13412 7880
rect 14096 7871 14148 7880
rect 6736 7735 6788 7744
rect 6736 7701 6745 7735
rect 6745 7701 6779 7735
rect 6779 7701 6788 7735
rect 6736 7692 6788 7701
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 10600 7692 10652 7744
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 12256 7803 12308 7812
rect 12256 7769 12281 7803
rect 12281 7769 12308 7803
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 16304 7828 16356 7880
rect 16488 7828 16540 7880
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 17040 7828 17092 7880
rect 12256 7760 12308 7769
rect 13820 7760 13872 7812
rect 17224 7828 17276 7880
rect 17408 7828 17460 7880
rect 19156 7828 19208 7880
rect 19984 7871 20036 7880
rect 19984 7837 20018 7871
rect 20018 7837 20036 7871
rect 18696 7760 18748 7812
rect 12808 7692 12860 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 16212 7692 16264 7744
rect 19340 7760 19392 7812
rect 19984 7828 20036 7837
rect 20720 7828 20772 7880
rect 22560 8032 22612 8084
rect 23480 8032 23532 8084
rect 23572 8032 23624 8084
rect 24400 8032 24452 8084
rect 21456 7896 21508 7948
rect 19892 7692 19944 7744
rect 21548 7803 21600 7812
rect 21548 7769 21557 7803
rect 21557 7769 21591 7803
rect 21591 7769 21600 7803
rect 21548 7760 21600 7769
rect 22192 7828 22244 7880
rect 22744 7828 22796 7880
rect 24584 7896 24636 7948
rect 25780 7896 25832 7948
rect 25872 7896 25924 7948
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 23296 7760 23348 7812
rect 24308 7760 24360 7812
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 21364 7692 21416 7744
rect 23848 7692 23900 7744
rect 24768 7692 24820 7744
rect 26976 7735 27028 7744
rect 26976 7701 26985 7735
rect 26985 7701 27019 7735
rect 27019 7701 27028 7735
rect 26976 7692 27028 7701
rect 28356 7692 28408 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 2320 7488 2372 7540
rect 2780 7488 2832 7540
rect 2872 7488 2924 7540
rect 3424 7531 3476 7540
rect 3424 7497 3433 7531
rect 3433 7497 3467 7531
rect 3467 7497 3476 7531
rect 3424 7488 3476 7497
rect 4436 7488 4488 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 5540 7488 5592 7540
rect 6552 7488 6604 7540
rect 6736 7488 6788 7540
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 5724 7420 5776 7472
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 7564 7352 7616 7404
rect 8024 7352 8076 7404
rect 10968 7488 11020 7540
rect 11244 7488 11296 7540
rect 11612 7488 11664 7540
rect 8208 7420 8260 7472
rect 12716 7488 12768 7540
rect 12808 7488 12860 7540
rect 12532 7420 12584 7472
rect 12992 7488 13044 7540
rect 13360 7420 13412 7472
rect 10232 7395 10284 7404
rect 10232 7361 10266 7395
rect 10266 7361 10284 7395
rect 10232 7352 10284 7361
rect 10600 7352 10652 7404
rect 11612 7352 11664 7404
rect 1676 7216 1728 7268
rect 9864 7284 9916 7336
rect 15292 7488 15344 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 16396 7488 16448 7540
rect 17132 7488 17184 7540
rect 17224 7488 17276 7540
rect 17500 7488 17552 7540
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 19800 7488 19852 7540
rect 21180 7488 21232 7540
rect 22100 7488 22152 7540
rect 23296 7531 23348 7540
rect 23296 7497 23305 7531
rect 23305 7497 23339 7531
rect 23339 7497 23348 7531
rect 23296 7488 23348 7497
rect 24124 7488 24176 7540
rect 24860 7488 24912 7540
rect 25780 7531 25832 7540
rect 25780 7497 25789 7531
rect 25789 7497 25823 7531
rect 25823 7497 25832 7531
rect 25780 7488 25832 7497
rect 26792 7531 26844 7540
rect 26792 7497 26801 7531
rect 26801 7497 26835 7531
rect 26835 7497 26844 7531
rect 26792 7488 26844 7497
rect 26976 7488 27028 7540
rect 28356 7531 28408 7540
rect 28356 7497 28365 7531
rect 28365 7497 28399 7531
rect 28399 7497 28408 7531
rect 28356 7488 28408 7497
rect 12992 7352 13044 7404
rect 13636 7352 13688 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 15568 7420 15620 7472
rect 16488 7420 16540 7472
rect 16672 7420 16724 7472
rect 16856 7352 16908 7404
rect 14280 7284 14332 7336
rect 17684 7352 17736 7404
rect 18604 7420 18656 7472
rect 23572 7420 23624 7472
rect 23848 7463 23900 7472
rect 23848 7429 23857 7463
rect 23857 7429 23891 7463
rect 23891 7429 23900 7463
rect 23848 7420 23900 7429
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 24400 7420 24452 7472
rect 26332 7463 26384 7472
rect 26332 7429 26341 7463
rect 26341 7429 26375 7463
rect 26375 7429 26384 7463
rect 26332 7420 26384 7429
rect 24492 7352 24544 7404
rect 5816 7148 5868 7200
rect 6092 7148 6144 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8208 7148 8260 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 16212 7216 16264 7268
rect 17684 7259 17736 7268
rect 17684 7225 17693 7259
rect 17693 7225 17727 7259
rect 17727 7225 17736 7259
rect 17684 7216 17736 7225
rect 18144 7216 18196 7268
rect 18972 7148 19024 7200
rect 19156 7148 19208 7200
rect 22100 7216 22152 7268
rect 24308 7216 24360 7268
rect 26608 7259 26660 7268
rect 26608 7225 26617 7259
rect 26617 7225 26651 7259
rect 26651 7225 26660 7259
rect 26608 7216 26660 7225
rect 22192 7148 22244 7200
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 3792 6944 3844 6996
rect 7012 6944 7064 6996
rect 7748 6944 7800 6996
rect 8024 6944 8076 6996
rect 2228 6740 2280 6792
rect 3148 6740 3200 6792
rect 1676 6672 1728 6724
rect 6644 6672 6696 6724
rect 9220 6808 9272 6860
rect 10232 6944 10284 6996
rect 10416 6944 10468 6996
rect 11244 6876 11296 6928
rect 11796 6944 11848 6996
rect 14188 6944 14240 6996
rect 16948 6944 17000 6996
rect 8392 6740 8444 6792
rect 8484 6740 8536 6792
rect 9956 6740 10008 6792
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 14740 6876 14792 6928
rect 18236 6944 18288 6996
rect 21456 6944 21508 6996
rect 22192 6944 22244 6996
rect 22560 6944 22612 6996
rect 24400 6944 24452 6996
rect 26700 6944 26752 6996
rect 15476 6808 15528 6860
rect 18144 6808 18196 6860
rect 23112 6876 23164 6928
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 13912 6740 13964 6792
rect 14096 6740 14148 6792
rect 8576 6672 8628 6724
rect 9128 6715 9180 6724
rect 9128 6681 9145 6715
rect 9145 6681 9180 6715
rect 9128 6672 9180 6681
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 3884 6604 3936 6656
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 10048 6715 10100 6724
rect 10048 6681 10057 6715
rect 10057 6681 10091 6715
rect 10091 6681 10100 6715
rect 10048 6672 10100 6681
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 13820 6672 13872 6724
rect 20720 6740 20772 6792
rect 21272 6740 21324 6792
rect 22284 6740 22336 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 25780 6783 25832 6792
rect 25780 6749 25789 6783
rect 25789 6749 25823 6783
rect 25823 6749 25832 6783
rect 25780 6740 25832 6749
rect 14464 6604 14516 6656
rect 17224 6672 17276 6724
rect 18052 6672 18104 6724
rect 18696 6672 18748 6724
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 21640 6672 21692 6724
rect 23756 6672 23808 6724
rect 26148 6672 26200 6724
rect 23020 6604 23072 6656
rect 23296 6604 23348 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1860 6400 1912 6452
rect 2228 6400 2280 6452
rect 756 6264 808 6316
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 4712 6400 4764 6452
rect 3240 6307 3292 6316
rect 3240 6273 3258 6307
rect 3258 6273 3292 6307
rect 3240 6264 3292 6273
rect 4804 6264 4856 6316
rect 6092 6443 6144 6452
rect 6092 6409 6101 6443
rect 6101 6409 6135 6443
rect 6135 6409 6144 6443
rect 6092 6400 6144 6409
rect 6552 6400 6604 6452
rect 8484 6400 8536 6452
rect 9680 6400 9732 6452
rect 9864 6400 9916 6452
rect 10508 6400 10560 6452
rect 12440 6400 12492 6452
rect 8576 6264 8628 6316
rect 13636 6400 13688 6452
rect 12716 6375 12768 6384
rect 12716 6341 12746 6375
rect 12746 6341 12768 6375
rect 12716 6332 12768 6341
rect 14004 6332 14056 6384
rect 14464 6375 14516 6384
rect 14464 6341 14473 6375
rect 14473 6341 14507 6375
rect 14507 6341 14516 6375
rect 14464 6332 14516 6341
rect 16120 6332 16172 6384
rect 17592 6400 17644 6452
rect 20260 6400 20312 6452
rect 21088 6400 21140 6452
rect 21640 6400 21692 6452
rect 23480 6400 23532 6452
rect 16764 6332 16816 6384
rect 9864 6264 9916 6316
rect 12348 6264 12400 6316
rect 12440 6264 12492 6316
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 19432 6332 19484 6384
rect 20904 6332 20956 6384
rect 4252 6196 4304 6248
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 11888 6196 11940 6248
rect 14280 6196 14332 6248
rect 3792 6128 3844 6180
rect 17132 6196 17184 6248
rect 17224 6196 17276 6248
rect 17500 6196 17552 6248
rect 18696 6264 18748 6316
rect 20536 6196 20588 6248
rect 4068 6060 4120 6112
rect 6736 6060 6788 6112
rect 14740 6128 14792 6180
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 14648 6060 14700 6112
rect 16120 6128 16172 6180
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 18236 6128 18288 6180
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 21364 6264 21416 6316
rect 22376 6332 22428 6384
rect 22744 6332 22796 6384
rect 23296 6264 23348 6316
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22192 6128 22244 6180
rect 23756 6375 23808 6384
rect 23756 6341 23765 6375
rect 23765 6341 23799 6375
rect 23799 6341 23808 6375
rect 24768 6400 24820 6452
rect 26148 6443 26200 6452
rect 26148 6409 26157 6443
rect 26157 6409 26191 6443
rect 26191 6409 26200 6443
rect 26148 6400 26200 6409
rect 23756 6332 23808 6341
rect 24860 6264 24912 6316
rect 24952 6128 25004 6180
rect 19340 6060 19392 6112
rect 20352 6103 20404 6112
rect 20352 6069 20361 6103
rect 20361 6069 20395 6103
rect 20395 6069 20404 6103
rect 20352 6060 20404 6069
rect 20444 6060 20496 6112
rect 20720 6060 20772 6112
rect 23388 6060 23440 6112
rect 24400 6060 24452 6112
rect 24492 6103 24544 6112
rect 24492 6069 24501 6103
rect 24501 6069 24535 6103
rect 24535 6069 24544 6103
rect 24492 6060 24544 6069
rect 25044 6103 25096 6112
rect 25044 6069 25053 6103
rect 25053 6069 25087 6103
rect 25087 6069 25096 6103
rect 25044 6060 25096 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6736 5856 6788 5908
rect 8484 5856 8536 5908
rect 9864 5856 9916 5908
rect 9956 5856 10008 5908
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 4160 5652 4212 5704
rect 6644 5652 6696 5704
rect 9772 5788 9824 5840
rect 9680 5720 9732 5772
rect 9220 5652 9272 5704
rect 7012 5584 7064 5636
rect 9128 5584 9180 5636
rect 12624 5856 12676 5908
rect 13176 5899 13228 5908
rect 13176 5865 13185 5899
rect 13185 5865 13219 5899
rect 13219 5865 13228 5899
rect 13176 5856 13228 5865
rect 13360 5856 13412 5908
rect 13728 5856 13780 5908
rect 14280 5856 14332 5908
rect 10140 5788 10192 5840
rect 11980 5831 12032 5840
rect 11980 5797 11989 5831
rect 11989 5797 12023 5831
rect 12023 5797 12032 5831
rect 11980 5788 12032 5797
rect 10508 5720 10560 5772
rect 10232 5652 10284 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 11888 5652 11940 5704
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 12532 5788 12584 5840
rect 14372 5788 14424 5840
rect 15660 5788 15712 5840
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 12900 5652 12952 5704
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 11704 5584 11756 5636
rect 14096 5652 14148 5704
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14280 5516 14332 5568
rect 15384 5652 15436 5704
rect 16120 5652 16172 5704
rect 16580 5856 16632 5908
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 17132 5856 17184 5908
rect 17316 5856 17368 5908
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 17960 5899 18012 5908
rect 17960 5865 17969 5899
rect 17969 5865 18003 5899
rect 18003 5865 18012 5899
rect 17960 5856 18012 5865
rect 18052 5856 18104 5908
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 14740 5584 14792 5636
rect 16856 5584 16908 5636
rect 17500 5627 17552 5636
rect 17500 5593 17509 5627
rect 17509 5593 17543 5627
rect 17543 5593 17552 5627
rect 17500 5584 17552 5593
rect 17868 5652 17920 5704
rect 19156 5856 19208 5908
rect 19432 5856 19484 5908
rect 20352 5856 20404 5908
rect 20812 5856 20864 5908
rect 20444 5720 20496 5772
rect 22192 5856 22244 5908
rect 24400 5899 24452 5908
rect 24400 5865 24409 5899
rect 24409 5865 24443 5899
rect 24443 5865 24452 5899
rect 24400 5856 24452 5865
rect 24492 5856 24544 5908
rect 25044 5856 25096 5908
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 16488 5516 16540 5568
rect 19340 5652 19392 5704
rect 18420 5516 18472 5568
rect 20720 5516 20772 5568
rect 21088 5627 21140 5636
rect 21088 5593 21097 5627
rect 21097 5593 21131 5627
rect 21131 5593 21140 5627
rect 21088 5584 21140 5593
rect 21364 5584 21416 5636
rect 25780 5695 25832 5704
rect 25780 5661 25789 5695
rect 25789 5661 25823 5695
rect 25823 5661 25832 5695
rect 25780 5652 25832 5661
rect 24952 5584 25004 5636
rect 23020 5516 23072 5568
rect 23756 5516 23808 5568
rect 25044 5516 25096 5568
rect 26056 5559 26108 5568
rect 26056 5525 26065 5559
rect 26065 5525 26099 5559
rect 26099 5525 26108 5559
rect 26056 5516 26108 5525
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 4160 5312 4212 5364
rect 4804 5312 4856 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7656 5312 7708 5364
rect 5264 5176 5316 5228
rect 6644 5244 6696 5296
rect 6828 5244 6880 5296
rect 5632 5108 5684 5160
rect 7288 5176 7340 5228
rect 10324 5312 10376 5364
rect 10416 5287 10468 5296
rect 10416 5253 10425 5287
rect 10425 5253 10459 5287
rect 10459 5253 10468 5287
rect 10416 5244 10468 5253
rect 12348 5312 12400 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 7656 5108 7708 5160
rect 8576 5176 8628 5228
rect 10048 5176 10100 5228
rect 11980 5244 12032 5296
rect 12624 5244 12676 5296
rect 9772 5108 9824 5160
rect 10876 5108 10928 5160
rect 14096 5244 14148 5296
rect 14556 5312 14608 5364
rect 14740 5355 14792 5364
rect 14740 5321 14749 5355
rect 14749 5321 14783 5355
rect 14783 5321 14792 5355
rect 14740 5312 14792 5321
rect 15384 5312 15436 5364
rect 15936 5312 15988 5364
rect 16672 5312 16724 5364
rect 16856 5312 16908 5364
rect 17684 5312 17736 5364
rect 18512 5355 18564 5364
rect 18512 5321 18534 5355
rect 18534 5321 18564 5355
rect 18512 5312 18564 5321
rect 14280 5176 14332 5228
rect 14648 5176 14700 5228
rect 17592 5244 17644 5296
rect 20536 5355 20588 5364
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 17224 5176 17276 5228
rect 14372 5108 14424 5160
rect 7472 4972 7524 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 11980 5015 12032 5024
rect 11980 4981 11989 5015
rect 11989 4981 12023 5015
rect 12023 4981 12032 5015
rect 11980 4972 12032 4981
rect 12624 5040 12676 5092
rect 17500 5108 17552 5160
rect 20260 5176 20312 5228
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 20996 5176 21048 5228
rect 22744 5244 22796 5296
rect 13636 4972 13688 5024
rect 17408 5040 17460 5092
rect 18880 5040 18932 5092
rect 19156 5040 19208 5092
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 16488 4972 16540 5024
rect 16580 4972 16632 5024
rect 17776 4972 17828 5024
rect 19064 4972 19116 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 20812 4972 20864 5024
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 22652 5176 22704 5228
rect 22744 5108 22796 5160
rect 23020 5244 23072 5296
rect 23388 5312 23440 5364
rect 23480 5176 23532 5228
rect 23756 5176 23808 5228
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 22928 5083 22980 5092
rect 22928 5049 22937 5083
rect 22937 5049 22971 5083
rect 22971 5049 22980 5083
rect 22928 5040 22980 5049
rect 23388 5151 23440 5160
rect 23388 5117 23397 5151
rect 23397 5117 23431 5151
rect 23431 5117 23440 5151
rect 23388 5108 23440 5117
rect 24676 5312 24728 5364
rect 24952 5355 25004 5364
rect 24952 5321 24961 5355
rect 24961 5321 24995 5355
rect 24995 5321 25004 5355
rect 24952 5312 25004 5321
rect 26056 5287 26108 5296
rect 26056 5253 26074 5287
rect 26074 5253 26108 5287
rect 26056 5244 26108 5253
rect 25780 5176 25832 5228
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 4804 4768 4856 4820
rect 7656 4768 7708 4820
rect 8944 4768 8996 4820
rect 10048 4768 10100 4820
rect 16580 4768 16632 4820
rect 17500 4768 17552 4820
rect 17776 4768 17828 4820
rect 18696 4768 18748 4820
rect 7288 4700 7340 4752
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 8484 4564 8536 4616
rect 9772 4632 9824 4684
rect 11704 4700 11756 4752
rect 12716 4743 12768 4752
rect 12716 4709 12725 4743
rect 12725 4709 12759 4743
rect 12759 4709 12768 4743
rect 12716 4700 12768 4709
rect 20260 4768 20312 4820
rect 20444 4768 20496 4820
rect 22652 4768 22704 4820
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 23388 4768 23440 4820
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 11152 4632 11204 4684
rect 14004 4632 14056 4684
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 11060 4564 11112 4616
rect 11980 4564 12032 4616
rect 756 4496 808 4548
rect 2136 4496 2188 4548
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 7288 4539 7340 4548
rect 7288 4505 7297 4539
rect 7297 4505 7331 4539
rect 7331 4505 7340 4539
rect 7288 4496 7340 4505
rect 9404 4496 9456 4548
rect 9588 4539 9640 4548
rect 9588 4505 9597 4539
rect 9597 4505 9631 4539
rect 9631 4505 9640 4539
rect 9588 4496 9640 4505
rect 9772 4539 9824 4548
rect 9772 4505 9807 4539
rect 9807 4505 9824 4539
rect 9772 4496 9824 4505
rect 13544 4564 13596 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17040 4564 17092 4616
rect 17132 4564 17184 4616
rect 12256 4496 12308 4548
rect 13912 4496 13964 4548
rect 18604 4564 18656 4616
rect 20076 4564 20128 4616
rect 22560 4632 22612 4684
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 11612 4428 11664 4480
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 19708 4496 19760 4548
rect 20996 4539 21048 4548
rect 20996 4505 21030 4539
rect 21030 4505 21048 4539
rect 20996 4496 21048 4505
rect 22836 4539 22888 4548
rect 22836 4505 22845 4539
rect 22845 4505 22879 4539
rect 22879 4505 22888 4539
rect 22836 4496 22888 4505
rect 23112 4496 23164 4548
rect 23296 4539 23348 4548
rect 23296 4505 23305 4539
rect 23305 4505 23339 4539
rect 23339 4505 23348 4539
rect 23296 4496 23348 4505
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23480 4564 23532 4573
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24860 4428 24912 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 6828 4224 6880 4276
rect 6920 4224 6972 4276
rect 8484 4224 8536 4276
rect 5632 4156 5684 4208
rect 9312 4224 9364 4276
rect 13452 4224 13504 4276
rect 9772 4156 9824 4208
rect 9864 4199 9916 4208
rect 9864 4165 9873 4199
rect 9873 4165 9907 4199
rect 9907 4165 9916 4199
rect 9864 4156 9916 4165
rect 10140 4156 10192 4208
rect 11152 4156 11204 4208
rect 11612 4156 11664 4208
rect 12256 4156 12308 4208
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 7932 4131 7984 4140
rect 7932 4097 7966 4131
rect 7966 4097 7984 4131
rect 7932 4088 7984 4097
rect 9036 4088 9088 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10508 4088 10560 4140
rect 12532 4156 12584 4208
rect 12900 4088 12952 4140
rect 14096 4156 14148 4208
rect 16488 4267 16540 4276
rect 16488 4233 16497 4267
rect 16497 4233 16531 4267
rect 16531 4233 16540 4267
rect 16488 4224 16540 4233
rect 15476 4156 15528 4208
rect 15844 4156 15896 4208
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 20812 4224 20864 4276
rect 20996 4224 21048 4276
rect 22560 4224 22612 4276
rect 23296 4224 23348 4276
rect 23480 4224 23532 4276
rect 17132 4156 17184 4208
rect 18696 4156 18748 4208
rect 15200 4088 15252 4140
rect 17500 4088 17552 4140
rect 18604 4088 18656 4140
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 9680 4020 9732 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 4068 3884 4120 3936
rect 6552 3884 6604 3936
rect 14740 4020 14792 4072
rect 23756 4156 23808 4208
rect 21640 4020 21692 4072
rect 22284 4088 22336 4140
rect 23848 4088 23900 4140
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 9220 3884 9272 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 10784 3884 10836 3936
rect 11244 3884 11296 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 19432 3995 19484 4004
rect 19432 3961 19441 3995
rect 19441 3961 19475 3995
rect 19475 3961 19484 3995
rect 19432 3952 19484 3961
rect 23572 3884 23624 3936
rect 25872 3952 25924 4004
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 5816 3680 5868 3732
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 6644 3680 6696 3732
rect 7656 3680 7708 3732
rect 7932 3680 7984 3732
rect 6552 3519 6604 3528
rect 6552 3485 6586 3519
rect 6586 3485 6604 3519
rect 6552 3476 6604 3485
rect 10600 3680 10652 3732
rect 11612 3680 11664 3732
rect 12164 3680 12216 3732
rect 12532 3680 12584 3732
rect 12716 3680 12768 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 14280 3680 14332 3732
rect 15660 3680 15712 3732
rect 17040 3680 17092 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 19432 3680 19484 3732
rect 23572 3680 23624 3732
rect 23848 3723 23900 3732
rect 23848 3689 23857 3723
rect 23857 3689 23891 3723
rect 23891 3689 23900 3723
rect 23848 3680 23900 3689
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 11704 3519 11756 3528
rect 11704 3485 11738 3519
rect 11738 3485 11756 3519
rect 9588 3408 9640 3460
rect 10232 3451 10284 3460
rect 10232 3417 10266 3451
rect 10266 3417 10284 3451
rect 10232 3408 10284 3417
rect 11704 3476 11756 3485
rect 13544 3612 13596 3664
rect 14004 3544 14056 3596
rect 12808 3476 12860 3528
rect 15844 3612 15896 3664
rect 16488 3612 16540 3664
rect 21272 3612 21324 3664
rect 17316 3476 17368 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 17500 3476 17552 3528
rect 10048 3340 10100 3392
rect 11244 3340 11296 3392
rect 11980 3340 12032 3392
rect 16672 3451 16724 3460
rect 13636 3340 13688 3392
rect 16672 3417 16681 3451
rect 16681 3417 16715 3451
rect 16715 3417 16724 3451
rect 16672 3408 16724 3417
rect 15844 3383 15896 3392
rect 15844 3349 15853 3383
rect 15853 3349 15887 3383
rect 15887 3349 15896 3383
rect 15844 3340 15896 3349
rect 19248 3451 19300 3460
rect 19248 3417 19257 3451
rect 19257 3417 19291 3451
rect 19291 3417 19300 3451
rect 19248 3408 19300 3417
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 23204 3544 23256 3596
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 10232 3136 10284 3188
rect 10324 3136 10376 3188
rect 10784 3136 10836 3188
rect 15200 3136 15252 3188
rect 9680 3068 9732 3120
rect 10048 3068 10100 3120
rect 16028 3068 16080 3120
rect 17408 3136 17460 3188
rect 22468 3179 22520 3188
rect 22468 3145 22477 3179
rect 22477 3145 22511 3179
rect 22511 3145 22520 3179
rect 22468 3136 22520 3145
rect 22836 3136 22888 3188
rect 19248 3068 19300 3120
rect 22284 3068 22336 3120
rect 11612 3000 11664 3052
rect 12256 3000 12308 3052
rect 15384 3000 15436 3052
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 11796 2796 11848 2848
rect 14740 2932 14792 2984
rect 18052 2864 18104 2916
rect 19708 2907 19760 2916
rect 19708 2873 19717 2907
rect 19717 2873 19751 2907
rect 19751 2873 19760 2907
rect 19708 2864 19760 2873
rect 21640 2864 21692 2916
rect 13452 2796 13504 2848
rect 19524 2839 19576 2848
rect 19524 2805 19533 2839
rect 19533 2805 19567 2839
rect 19567 2805 19576 2839
rect 19524 2796 19576 2805
rect 20812 2839 20864 2848
rect 20812 2805 20821 2839
rect 20821 2805 20855 2839
rect 20855 2805 20864 2839
rect 20812 2796 20864 2805
rect 25044 2932 25096 2984
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 7748 2592 7800 2644
rect 11980 2592 12032 2644
rect 13268 2592 13320 2644
rect 6644 2456 6696 2508
rect 9680 2524 9732 2576
rect 9772 2524 9824 2576
rect 11244 2499 11296 2508
rect 11244 2465 11253 2499
rect 11253 2465 11287 2499
rect 11287 2465 11296 2499
rect 11244 2456 11296 2465
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 15384 2635 15436 2644
rect 15384 2601 15393 2635
rect 15393 2601 15427 2635
rect 15427 2601 15436 2635
rect 15384 2592 15436 2601
rect 18052 2592 18104 2644
rect 18880 2592 18932 2644
rect 19708 2592 19760 2644
rect 20352 2592 20404 2644
rect 22652 2592 22704 2644
rect 23020 2524 23072 2576
rect 7196 2320 7248 2372
rect 9036 2320 9088 2372
rect 9496 2295 9548 2304
rect 9496 2261 9505 2295
rect 9505 2261 9539 2295
rect 9539 2261 9548 2295
rect 9496 2252 9548 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 13452 2363 13504 2372
rect 13452 2329 13461 2363
rect 13461 2329 13495 2363
rect 13495 2329 13504 2363
rect 13452 2320 13504 2329
rect 15844 2388 15896 2440
rect 17500 2388 17552 2440
rect 19892 2388 19944 2440
rect 20812 2388 20864 2440
rect 14372 2252 14424 2304
rect 16488 2320 16540 2372
rect 19616 2320 19668 2372
rect 22284 2363 22336 2372
rect 22284 2329 22293 2363
rect 22293 2329 22327 2363
rect 22327 2329 22336 2363
rect 22284 2320 22336 2329
rect 18696 2252 18748 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 7196 2091 7248 2100
rect 7196 2057 7205 2091
rect 7205 2057 7239 2091
rect 7239 2057 7248 2091
rect 7196 2048 7248 2057
rect 6644 1912 6696 1964
rect 9036 2048 9088 2100
rect 9772 2048 9824 2100
rect 10048 2048 10100 2100
rect 8484 1980 8536 2032
rect 9680 1980 9732 2032
rect 10232 2023 10284 2032
rect 10232 1989 10266 2023
rect 10266 1989 10284 2023
rect 10232 1980 10284 1989
rect 11244 1980 11296 2032
rect 9956 1955 10008 1964
rect 9956 1921 9965 1955
rect 9965 1921 9999 1955
rect 9999 1921 10008 1955
rect 9956 1912 10008 1921
rect 11980 1912 12032 1964
rect 12164 1912 12216 1964
rect 13452 1980 13504 2032
rect 16488 2091 16540 2100
rect 16488 2057 16497 2091
rect 16497 2057 16531 2091
rect 16531 2057 16540 2091
rect 16488 2048 16540 2057
rect 17500 2048 17552 2100
rect 18696 2091 18748 2100
rect 18696 2057 18705 2091
rect 18705 2057 18739 2091
rect 18739 2057 18748 2091
rect 18696 2048 18748 2057
rect 19524 2048 19576 2100
rect 19616 2091 19668 2100
rect 19616 2057 19625 2091
rect 19625 2057 19659 2091
rect 19659 2057 19668 2091
rect 19616 2048 19668 2057
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 7932 1887 7984 1896
rect 7932 1853 7941 1887
rect 7941 1853 7975 1887
rect 7975 1853 7984 1887
rect 7932 1844 7984 1853
rect 14464 1844 14516 1896
rect 17408 1912 17460 1964
rect 9864 1776 9916 1828
rect 11888 1819 11940 1828
rect 11888 1785 11897 1819
rect 11897 1785 11931 1819
rect 11931 1785 11940 1819
rect 11888 1776 11940 1785
rect 16396 1776 16448 1828
rect 11980 1751 12032 1760
rect 11980 1717 11989 1751
rect 11989 1717 12023 1751
rect 12023 1717 12032 1751
rect 11980 1708 12032 1717
rect 13728 1708 13780 1760
rect 17040 1708 17092 1760
rect 19248 1912 19300 1964
rect 23020 2048 23072 2100
rect 19616 1912 19668 1964
rect 21456 1955 21508 1964
rect 21456 1921 21465 1955
rect 21465 1921 21499 1955
rect 21499 1921 21508 1955
rect 21456 1912 21508 1921
rect 21640 1912 21692 1964
rect 19892 1887 19944 1896
rect 19892 1853 19901 1887
rect 19901 1853 19935 1887
rect 19935 1853 19944 1887
rect 19892 1844 19944 1853
rect 18880 1776 18932 1828
rect 19248 1751 19300 1760
rect 19248 1717 19257 1751
rect 19257 1717 19291 1751
rect 19291 1717 19300 1751
rect 19248 1708 19300 1717
rect 22192 1708 22244 1760
rect 4423 1606 4475 1658
rect 4487 1606 4539 1658
rect 4551 1606 4603 1658
rect 4615 1606 4667 1658
rect 4679 1606 4731 1658
rect 11369 1606 11421 1658
rect 11433 1606 11485 1658
rect 11497 1606 11549 1658
rect 11561 1606 11613 1658
rect 11625 1606 11677 1658
rect 18315 1606 18367 1658
rect 18379 1606 18431 1658
rect 18443 1606 18495 1658
rect 18507 1606 18559 1658
rect 18571 1606 18623 1658
rect 25261 1606 25313 1658
rect 25325 1606 25377 1658
rect 25389 1606 25441 1658
rect 25453 1606 25505 1658
rect 25517 1606 25569 1658
rect 9864 1504 9916 1556
rect 12164 1547 12216 1556
rect 12164 1513 12173 1547
rect 12173 1513 12207 1547
rect 12207 1513 12216 1547
rect 12164 1504 12216 1513
rect 16396 1504 16448 1556
rect 17408 1547 17460 1556
rect 17408 1513 17417 1547
rect 17417 1513 17451 1547
rect 17451 1513 17460 1547
rect 17408 1504 17460 1513
rect 19156 1504 19208 1556
rect 19616 1547 19668 1556
rect 19616 1513 19625 1547
rect 19625 1513 19659 1547
rect 19659 1513 19668 1547
rect 19616 1504 19668 1513
rect 21456 1504 21508 1556
rect 17040 1479 17092 1488
rect 17040 1445 17049 1479
rect 17049 1445 17083 1479
rect 17083 1445 17092 1479
rect 17040 1436 17092 1445
rect 22192 1436 22244 1488
rect 7932 1368 7984 1420
rect 22284 1411 22336 1420
rect 22284 1377 22293 1411
rect 22293 1377 22327 1411
rect 22327 1377 22336 1411
rect 22284 1368 22336 1377
rect 9496 1300 9548 1352
rect 11980 1343 12032 1352
rect 11980 1309 11989 1343
rect 11989 1309 12023 1343
rect 12023 1309 12032 1343
rect 11980 1300 12032 1309
rect 14372 1343 14424 1352
rect 14372 1309 14406 1343
rect 14406 1309 14424 1343
rect 14372 1300 14424 1309
rect 14740 1300 14792 1352
rect 16672 1343 16724 1352
rect 16672 1309 16681 1343
rect 16681 1309 16715 1343
rect 16715 1309 16724 1343
rect 16672 1300 16724 1309
rect 19248 1300 19300 1352
rect 7896 1062 7948 1114
rect 7960 1062 8012 1114
rect 8024 1062 8076 1114
rect 8088 1062 8140 1114
rect 8152 1062 8204 1114
rect 14842 1062 14894 1114
rect 14906 1062 14958 1114
rect 14970 1062 15022 1114
rect 15034 1062 15086 1114
rect 15098 1062 15150 1114
rect 21788 1062 21840 1114
rect 21852 1062 21904 1114
rect 21916 1062 21968 1114
rect 21980 1062 22032 1114
rect 22044 1062 22096 1114
rect 28734 1062 28786 1114
rect 28798 1062 28850 1114
rect 28862 1062 28914 1114
rect 28926 1062 28978 1114
rect 28990 1062 29042 1114
<< metal2 >>
rect 7896 32668 8204 32677
rect 7896 32666 7902 32668
rect 7958 32666 7982 32668
rect 8038 32666 8062 32668
rect 8118 32666 8142 32668
rect 8198 32666 8204 32668
rect 7958 32614 7960 32666
rect 8140 32614 8142 32666
rect 7896 32612 7902 32614
rect 7958 32612 7982 32614
rect 8038 32612 8062 32614
rect 8118 32612 8142 32614
rect 8198 32612 8204 32614
rect 7896 32603 8204 32612
rect 14842 32668 15150 32677
rect 14842 32666 14848 32668
rect 14904 32666 14928 32668
rect 14984 32666 15008 32668
rect 15064 32666 15088 32668
rect 15144 32666 15150 32668
rect 14904 32614 14906 32666
rect 15086 32614 15088 32666
rect 14842 32612 14848 32614
rect 14904 32612 14928 32614
rect 14984 32612 15008 32614
rect 15064 32612 15088 32614
rect 15144 32612 15150 32614
rect 14842 32603 15150 32612
rect 21788 32668 22096 32677
rect 21788 32666 21794 32668
rect 21850 32666 21874 32668
rect 21930 32666 21954 32668
rect 22010 32666 22034 32668
rect 22090 32666 22096 32668
rect 21850 32614 21852 32666
rect 22032 32614 22034 32666
rect 21788 32612 21794 32614
rect 21850 32612 21874 32614
rect 21930 32612 21954 32614
rect 22010 32612 22034 32614
rect 22090 32612 22096 32614
rect 21788 32603 22096 32612
rect 28734 32668 29042 32677
rect 28734 32666 28740 32668
rect 28796 32666 28820 32668
rect 28876 32666 28900 32668
rect 28956 32666 28980 32668
rect 29036 32666 29042 32668
rect 28796 32614 28798 32666
rect 28978 32614 28980 32666
rect 28734 32612 28740 32614
rect 28796 32612 28820 32614
rect 28876 32612 28900 32614
rect 28956 32612 28980 32614
rect 29036 32612 29042 32614
rect 28734 32603 29042 32612
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 4252 32360 4304 32366
rect 4252 32302 4304 32308
rect 6460 32360 6512 32366
rect 6460 32302 6512 32308
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 3988 31822 4016 32302
rect 4264 31958 4292 32302
rect 4344 32224 4396 32230
rect 4344 32166 4396 32172
rect 4252 31952 4304 31958
rect 4252 31894 4304 31900
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 2412 31476 2464 31482
rect 2412 31418 2464 31424
rect 2424 31142 2452 31418
rect 3988 31346 4016 31758
rect 4264 31346 4292 31894
rect 4356 31686 4384 32166
rect 4423 32124 4731 32133
rect 4423 32122 4429 32124
rect 4485 32122 4509 32124
rect 4565 32122 4589 32124
rect 4645 32122 4669 32124
rect 4725 32122 4731 32124
rect 4485 32070 4487 32122
rect 4667 32070 4669 32122
rect 4423 32068 4429 32070
rect 4485 32068 4509 32070
rect 4565 32068 4589 32070
rect 4645 32068 4669 32070
rect 4725 32068 4731 32070
rect 4423 32059 4731 32068
rect 6472 31890 6500 32302
rect 7852 31890 7880 32302
rect 9600 31890 9628 32302
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 32026 11100 32166
rect 11369 32124 11677 32133
rect 11369 32122 11375 32124
rect 11431 32122 11455 32124
rect 11511 32122 11535 32124
rect 11591 32122 11615 32124
rect 11671 32122 11677 32124
rect 11431 32070 11433 32122
rect 11613 32070 11615 32122
rect 11369 32068 11375 32070
rect 11431 32068 11455 32070
rect 11511 32068 11535 32070
rect 11591 32068 11615 32070
rect 11671 32068 11677 32070
rect 11369 32059 11677 32068
rect 18315 32124 18623 32133
rect 18315 32122 18321 32124
rect 18377 32122 18401 32124
rect 18457 32122 18481 32124
rect 18537 32122 18561 32124
rect 18617 32122 18623 32124
rect 18377 32070 18379 32122
rect 18559 32070 18561 32122
rect 18315 32068 18321 32070
rect 18377 32068 18401 32070
rect 18457 32068 18481 32070
rect 18537 32068 18561 32070
rect 18617 32068 18623 32070
rect 18315 32059 18623 32068
rect 25261 32124 25569 32133
rect 25261 32122 25267 32124
rect 25323 32122 25347 32124
rect 25403 32122 25427 32124
rect 25483 32122 25507 32124
rect 25563 32122 25569 32124
rect 25323 32070 25325 32122
rect 25505 32070 25507 32122
rect 25261 32068 25267 32070
rect 25323 32068 25347 32070
rect 25403 32068 25427 32070
rect 25483 32068 25507 32070
rect 25563 32068 25569 32070
rect 25261 32059 25569 32068
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 6460 31884 6512 31890
rect 6460 31826 6512 31832
rect 7840 31884 7892 31890
rect 7840 31826 7892 31832
rect 9588 31884 9640 31890
rect 9588 31826 9640 31832
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 8668 31816 8720 31822
rect 8668 31758 8720 31764
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 4344 31680 4396 31686
rect 4344 31622 4396 31628
rect 4356 31482 4384 31622
rect 4344 31476 4396 31482
rect 4344 31418 4396 31424
rect 2504 31340 2556 31346
rect 2504 31282 2556 31288
rect 3976 31340 4028 31346
rect 3976 31282 4028 31288
rect 4252 31340 4304 31346
rect 4252 31282 4304 31288
rect 1860 31136 1912 31142
rect 1030 31104 1086 31113
rect 1860 31078 1912 31084
rect 2412 31136 2464 31142
rect 2412 31078 2464 31084
rect 1030 31039 1086 31048
rect 1044 30938 1072 31039
rect 1032 30932 1084 30938
rect 1032 30874 1084 30880
rect 1872 30734 1900 31078
rect 2516 30802 2544 31282
rect 3056 31204 3108 31210
rect 3056 31146 3108 31152
rect 2780 31136 2832 31142
rect 2780 31078 2832 31084
rect 1952 30796 2004 30802
rect 1952 30738 2004 30744
rect 2504 30796 2556 30802
rect 2504 30738 2556 30744
rect 1860 30728 1912 30734
rect 1860 30670 1912 30676
rect 1860 30592 1912 30598
rect 1860 30534 1912 30540
rect 1872 29714 1900 30534
rect 1964 30190 1992 30738
rect 2792 30734 2820 31078
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2872 30660 2924 30666
rect 2872 30602 2924 30608
rect 1952 30184 2004 30190
rect 1952 30126 2004 30132
rect 2688 30048 2740 30054
rect 2688 29990 2740 29996
rect 1860 29708 1912 29714
rect 1860 29650 1912 29656
rect 2136 29708 2188 29714
rect 2136 29650 2188 29656
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1596 28762 1624 29135
rect 1780 29050 1808 29582
rect 1860 29504 1912 29510
rect 1860 29446 1912 29452
rect 1872 29306 1900 29446
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 2148 29170 2176 29650
rect 2700 29646 2728 29990
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2136 29164 2188 29170
rect 2136 29106 2188 29112
rect 2780 29096 2832 29102
rect 1780 29034 1900 29050
rect 2780 29038 2832 29044
rect 1780 29028 1912 29034
rect 1780 29022 1860 29028
rect 1860 28970 1912 28976
rect 1584 28756 1636 28762
rect 1584 28698 1636 28704
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1780 28218 1808 28494
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1676 27532 1728 27538
rect 1676 27474 1728 27480
rect 1688 27130 1716 27474
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1872 27010 1900 28970
rect 2792 28762 2820 29038
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2044 28552 2096 28558
rect 2044 28494 2096 28500
rect 2056 28082 2084 28494
rect 2136 28416 2188 28422
rect 2136 28358 2188 28364
rect 2148 28218 2176 28358
rect 2136 28212 2188 28218
rect 2136 28154 2188 28160
rect 2596 28144 2648 28150
rect 2596 28086 2648 28092
rect 2044 28076 2096 28082
rect 2044 28018 2096 28024
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2516 27470 2544 28018
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2504 27464 2556 27470
rect 2504 27406 2556 27412
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2136 27328 2188 27334
rect 2136 27270 2188 27276
rect 1688 26982 1900 27010
rect 2056 26994 2084 27270
rect 2148 27130 2176 27270
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 2044 26988 2096 26994
rect 1398 24984 1454 24993
rect 1398 24919 1454 24928
rect 1412 24274 1440 24919
rect 1492 24608 1544 24614
rect 1492 24550 1544 24556
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1306 21584 1362 21593
rect 1306 21519 1362 21528
rect 1320 21418 1348 21519
rect 1308 21412 1360 21418
rect 1308 21354 1360 21360
rect 756 19780 808 19786
rect 756 19722 808 19728
rect 768 19689 796 19722
rect 754 19680 810 19689
rect 754 19615 810 19624
rect 1504 19334 1532 24550
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1596 22642 1624 23122
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1688 22234 1716 26982
rect 2044 26930 2096 26936
rect 2240 26926 2268 27406
rect 2516 27062 2544 27406
rect 2504 27056 2556 27062
rect 2504 26998 2556 27004
rect 2228 26920 2280 26926
rect 2228 26862 2280 26868
rect 2136 26240 2188 26246
rect 2136 26182 2188 26188
rect 2148 26042 2176 26182
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2240 25906 2268 26862
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 2320 25900 2372 25906
rect 2320 25842 2372 25848
rect 2332 25498 2360 25842
rect 2412 25764 2464 25770
rect 2412 25706 2464 25712
rect 2320 25492 2372 25498
rect 2320 25434 2372 25440
rect 2228 24880 2280 24886
rect 2228 24822 2280 24828
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 1964 23730 1992 24142
rect 2240 23866 2268 24822
rect 2320 24676 2372 24682
rect 2320 24618 2372 24624
rect 2332 24342 2360 24618
rect 2320 24336 2372 24342
rect 2320 24278 2372 24284
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2332 23730 2360 24142
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2320 23724 2372 23730
rect 2320 23666 2372 23672
rect 1964 23202 1992 23666
rect 2148 23254 2176 23666
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 1780 23174 1992 23202
rect 2136 23248 2188 23254
rect 2136 23190 2188 23196
rect 1780 22778 1808 23174
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1872 22030 1900 23054
rect 1952 23044 2004 23050
rect 1952 22986 2004 22992
rect 1964 22438 1992 22986
rect 2240 22574 2268 23462
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 2228 22568 2280 22574
rect 2228 22510 2280 22516
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 1964 22094 1992 22170
rect 1964 22066 2084 22094
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 2056 21842 2084 22066
rect 2148 22030 2176 22374
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2136 21888 2188 21894
rect 2056 21836 2136 21842
rect 2056 21830 2188 21836
rect 2056 21814 2176 21830
rect 2148 21486 2176 21814
rect 2240 21622 2268 22510
rect 2332 22166 2360 22714
rect 2320 22160 2372 22166
rect 2320 22102 2372 22108
rect 2228 21616 2280 21622
rect 2228 21558 2280 21564
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2240 19718 2268 21558
rect 2332 21350 2360 22102
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2424 21146 2452 25706
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2516 23594 2544 24754
rect 2608 24410 2636 28086
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2792 27452 2820 27814
rect 2884 27606 2912 30602
rect 3068 30598 3096 31146
rect 3988 30938 4016 31282
rect 4264 30938 4292 31282
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 4252 30932 4304 30938
rect 4252 30874 4304 30880
rect 4356 30734 4384 31418
rect 5000 31346 5028 31758
rect 7300 31346 7328 31758
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 4816 30870 4844 31214
rect 5000 30938 5028 31282
rect 8484 31272 8536 31278
rect 8484 31214 8536 31220
rect 8496 30938 8524 31214
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 4804 30864 4856 30870
rect 4804 30806 4856 30812
rect 8680 30734 8708 31758
rect 9324 31278 9352 31758
rect 9692 31686 9720 31758
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9600 31346 9628 31622
rect 9692 31346 9720 31622
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 8944 31136 8996 31142
rect 8944 31078 8996 31084
rect 8956 30734 8984 31078
rect 9324 30802 9352 31214
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9312 30796 9364 30802
rect 9312 30738 9364 30744
rect 9416 30734 9444 31078
rect 9600 30802 9628 31282
rect 9692 31142 9720 31282
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9956 30864 10008 30870
rect 9956 30806 10008 30812
rect 9588 30796 9640 30802
rect 9588 30738 9640 30744
rect 4344 30728 4396 30734
rect 4344 30670 4396 30676
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 5724 30728 5776 30734
rect 5724 30670 5776 30676
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8944 30728 8996 30734
rect 8944 30670 8996 30676
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 3056 30592 3108 30598
rect 3056 30534 3108 30540
rect 3424 30592 3476 30598
rect 3424 30534 3476 30540
rect 3068 30394 3096 30534
rect 3056 30388 3108 30394
rect 3056 30330 3108 30336
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2976 29170 3004 30126
rect 3068 29510 3096 30330
rect 3436 30190 3464 30534
rect 4816 30394 4844 30670
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4068 30320 4120 30326
rect 4068 30262 4120 30268
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3884 30184 3936 30190
rect 3884 30126 3936 30132
rect 3252 29850 3280 30126
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3056 29504 3108 29510
rect 3056 29446 3108 29452
rect 3068 29306 3096 29446
rect 3056 29300 3108 29306
rect 3056 29242 3108 29248
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2976 28422 3004 29106
rect 3068 29034 3096 29242
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3056 29028 3108 29034
rect 3056 28970 3108 28976
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2872 27600 2924 27606
rect 2872 27542 2924 27548
rect 2792 27424 2912 27452
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2700 23798 2728 26386
rect 2792 25362 2820 27231
rect 2884 26858 2912 27424
rect 2976 26858 3004 28358
rect 3068 27878 3096 28970
rect 3252 28422 3280 29106
rect 3240 28416 3292 28422
rect 3240 28358 3292 28364
rect 3148 28008 3200 28014
rect 3148 27950 3200 27956
rect 3056 27872 3108 27878
rect 3056 27814 3108 27820
rect 3160 27470 3188 27950
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3252 27418 3280 28358
rect 3332 27872 3384 27878
rect 3332 27814 3384 27820
rect 3344 27538 3372 27814
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3252 27390 3372 27418
rect 3344 26994 3372 27390
rect 3056 26988 3108 26994
rect 3056 26930 3108 26936
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2872 26852 2924 26858
rect 2872 26794 2924 26800
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 2872 26580 2924 26586
rect 2872 26522 2924 26528
rect 2884 25974 2912 26522
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2872 25968 2924 25974
rect 2872 25910 2924 25916
rect 2872 25832 2924 25838
rect 2976 25786 3004 26318
rect 3068 25974 3096 26930
rect 3344 26586 3372 26930
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3436 26466 3464 30126
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3528 29238 3556 29446
rect 3516 29232 3568 29238
rect 3516 29174 3568 29180
rect 3896 29170 3924 30126
rect 4080 29238 4108 30262
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 4068 29232 4120 29238
rect 4068 29174 4120 29180
rect 3884 29164 3936 29170
rect 3884 29106 3936 29112
rect 3516 28416 3568 28422
rect 3516 28358 3568 28364
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 3528 28218 3556 28358
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3528 27713 3556 28018
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3252 26438 3464 26466
rect 3056 25968 3108 25974
rect 3056 25910 3108 25916
rect 3068 25838 3096 25910
rect 3148 25900 3200 25906
rect 3148 25842 3200 25848
rect 2924 25780 3004 25786
rect 2872 25774 3004 25780
rect 3056 25832 3108 25838
rect 3056 25774 3108 25780
rect 2884 25758 3004 25774
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2884 24682 2912 25758
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2872 24676 2924 24682
rect 2872 24618 2924 24624
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 24274 2820 24550
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 2964 24132 3016 24138
rect 2964 24074 3016 24080
rect 2792 23866 2820 24074
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2688 23792 2740 23798
rect 2688 23734 2740 23740
rect 2504 23588 2556 23594
rect 2504 23530 2556 23536
rect 2516 22982 2544 23530
rect 2778 23488 2834 23497
rect 2778 23423 2834 23432
rect 2596 23248 2648 23254
rect 2596 23190 2648 23196
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2608 22778 2636 23190
rect 2688 23044 2740 23050
rect 2688 22986 2740 22992
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2608 21690 2636 22714
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2700 21010 2728 22986
rect 2792 22778 2820 23423
rect 2976 23322 3004 24074
rect 2964 23316 3016 23322
rect 2964 23258 3016 23264
rect 2964 23112 3016 23118
rect 3068 23100 3096 25638
rect 3160 24721 3188 25842
rect 3146 24712 3202 24721
rect 3146 24647 3202 24656
rect 3252 24274 3280 26438
rect 3528 26382 3556 26930
rect 3608 26852 3660 26858
rect 3608 26794 3660 26800
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 3332 25288 3384 25294
rect 3332 25230 3384 25236
rect 3344 24410 3372 25230
rect 3436 24614 3464 26250
rect 3620 25702 3648 26794
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3712 25906 3740 26726
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3528 24993 3556 25638
rect 3620 25498 3648 25638
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3514 24984 3570 24993
rect 3514 24919 3570 24928
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 3160 23730 3188 24074
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3148 23588 3200 23594
rect 3148 23530 3200 23536
rect 3016 23072 3096 23100
rect 2964 23054 3016 23060
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2872 22704 2924 22710
rect 2792 22652 2872 22658
rect 2792 22646 2924 22652
rect 2792 22630 2912 22646
rect 3160 22642 3188 23530
rect 3252 22642 3280 24210
rect 3436 23118 3464 24550
rect 3712 24274 3740 25094
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3712 23882 3740 24210
rect 3620 23854 3740 23882
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3148 22636 3200 22642
rect 2792 22098 2820 22630
rect 3148 22578 3200 22584
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 2964 22500 3016 22506
rect 2964 22442 3016 22448
rect 2780 22092 2832 22098
rect 2976 22094 3004 22442
rect 2780 22034 2832 22040
rect 2884 22066 3004 22094
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2792 21146 2820 21558
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2688 21004 2740 21010
rect 2608 20964 2688 20992
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2332 19922 2360 20742
rect 2608 20058 2636 20964
rect 2688 20946 2740 20952
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1412 19306 1532 19334
rect 756 16108 808 16114
rect 756 16050 808 16056
rect 768 15881 796 16050
rect 754 15872 810 15881
rect 754 15807 810 15816
rect 754 13968 810 13977
rect 754 13903 756 13912
rect 808 13903 810 13912
rect 756 13874 808 13880
rect 1412 13530 1440 19306
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1688 18970 1716 19246
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1780 18426 1808 19246
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17882 1808 18226
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 17066 1624 17478
rect 1688 17270 1716 17546
rect 1676 17264 1728 17270
rect 1676 17206 1728 17212
rect 1584 17060 1636 17066
rect 1584 17002 1636 17008
rect 1596 14074 1624 17002
rect 1688 16182 1716 17206
rect 1780 16998 1808 17818
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 15094 1716 15302
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12442 1716 12786
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1780 12374 1808 16934
rect 2056 16522 2084 19450
rect 2424 18834 2452 19654
rect 2516 19514 2544 19790
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2700 19174 2728 19994
rect 2884 19718 2912 22066
rect 3068 21690 3096 22510
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3068 21078 3096 21626
rect 3056 21072 3108 21078
rect 3056 21014 3108 21020
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19372 2832 19378
rect 2976 19360 3004 19926
rect 2832 19332 3004 19360
rect 2780 19314 2832 19320
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18970 2728 19110
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2332 18426 2360 18770
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2332 18290 2360 18362
rect 2608 18358 2636 18702
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2134 18184 2190 18193
rect 2134 18119 2190 18128
rect 2148 17338 2176 18119
rect 2516 17610 2544 18226
rect 2700 18154 2728 18906
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2792 17785 2820 19178
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2884 18766 2912 19110
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 2056 15502 2084 16458
rect 2884 16250 2912 17138
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2976 16182 3004 19332
rect 3068 18766 3096 21014
rect 3160 20942 3188 22578
rect 3344 21690 3372 22578
rect 3516 22092 3568 22098
rect 3516 22034 3568 22040
rect 3424 21956 3476 21962
rect 3424 21898 3476 21904
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3252 21010 3280 21286
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 3160 20602 3188 20878
rect 3148 20596 3200 20602
rect 3200 20556 3280 20584
rect 3148 20538 3200 20544
rect 3252 20398 3280 20556
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3160 20058 3188 20334
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3252 19990 3280 20198
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3252 19854 3280 19926
rect 3240 19848 3292 19854
rect 3344 19836 3372 20334
rect 3436 20058 3464 21898
rect 3528 21078 3556 22034
rect 3516 21072 3568 21078
rect 3516 21014 3568 21020
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3424 19848 3476 19854
rect 3344 19808 3424 19836
rect 3240 19790 3292 19796
rect 3424 19790 3476 19796
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19378 3188 19654
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3054 17504 3110 17513
rect 3054 17439 3110 17448
rect 3068 17338 3096 17439
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 3160 16046 3188 19314
rect 3252 18426 3280 19790
rect 3436 19258 3464 19790
rect 3528 19378 3556 21014
rect 3620 20602 3648 23854
rect 3698 23488 3754 23497
rect 3698 23423 3754 23432
rect 3712 22778 3740 23423
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3620 19378 3648 20198
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3436 19230 3648 19258
rect 3620 18630 3648 19230
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3528 18426 3556 18566
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3252 17678 3280 18362
rect 3514 18320 3570 18329
rect 3332 18284 3384 18290
rect 3620 18290 3648 18566
rect 3514 18255 3570 18264
rect 3608 18284 3660 18290
rect 3332 18226 3384 18232
rect 3344 18154 3372 18226
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3344 17678 3372 18090
rect 3528 17882 3556 18255
rect 3608 18226 3660 18232
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 17338 3372 17614
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3516 16584 3568 16590
rect 3712 16572 3740 22714
rect 3804 22166 3832 28358
rect 4264 28082 4292 29582
rect 4816 29102 4844 29786
rect 5080 29572 5132 29578
rect 5080 29514 5132 29520
rect 5092 29306 5120 29514
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 5448 29232 5500 29238
rect 5448 29174 5500 29180
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4988 29096 5040 29102
rect 4988 29038 5040 29044
rect 4252 28076 4304 28082
rect 4252 28018 4304 28024
rect 4264 27674 4292 28018
rect 4252 27668 4304 27674
rect 4252 27610 4304 27616
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 4252 27328 4304 27334
rect 4252 27270 4304 27276
rect 4172 27062 4200 27270
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4264 26042 4292 27270
rect 4356 26518 4384 29038
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 4816 27606 4844 28018
rect 4804 27600 4856 27606
rect 4804 27542 4856 27548
rect 5000 27538 5028 29038
rect 5184 28762 5212 29106
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5460 28694 5488 29174
rect 5736 29034 5764 30670
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 7196 30252 7248 30258
rect 7196 30194 7248 30200
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6000 29504 6052 29510
rect 6000 29446 6052 29452
rect 6012 29102 6040 29446
rect 6000 29096 6052 29102
rect 6000 29038 6052 29044
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5448 28688 5500 28694
rect 5448 28630 5500 28636
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4816 26568 4844 27406
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4724 26540 4844 26568
rect 4344 26512 4396 26518
rect 4344 26454 4396 26460
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 4344 26240 4396 26246
rect 4344 26182 4396 26188
rect 4356 26042 4384 26182
rect 4252 26036 4304 26042
rect 4252 25978 4304 25984
rect 4344 26036 4396 26042
rect 4344 25978 4396 25984
rect 4356 25922 4384 25978
rect 4540 25974 4568 26318
rect 3976 25900 4028 25906
rect 3896 25860 3976 25888
rect 3896 24274 3924 25860
rect 3976 25842 4028 25848
rect 4264 25894 4384 25922
rect 4528 25968 4580 25974
rect 4528 25910 4580 25916
rect 4264 25378 4292 25894
rect 4540 25770 4568 25910
rect 4724 25906 4752 26540
rect 4802 26480 4858 26489
rect 4802 26415 4858 26424
rect 4816 26382 4844 26415
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4908 25974 4936 27270
rect 5092 26790 5120 27814
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5184 27130 5212 27406
rect 5172 27124 5224 27130
rect 5172 27066 5224 27072
rect 5276 27033 5304 27882
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5262 27024 5318 27033
rect 5262 26959 5318 26968
rect 5276 26926 5304 26959
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 4988 26580 5040 26586
rect 4988 26522 5040 26528
rect 4896 25968 4948 25974
rect 4816 25928 4896 25956
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 4344 25764 4396 25770
rect 4344 25706 4396 25712
rect 4528 25764 4580 25770
rect 4528 25706 4580 25712
rect 4356 25498 4384 25706
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4344 25492 4396 25498
rect 4816 25480 4844 25928
rect 4896 25910 4948 25916
rect 4896 25832 4948 25838
rect 4896 25774 4948 25780
rect 4344 25434 4396 25440
rect 4724 25452 4844 25480
rect 4264 25350 4384 25378
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 4172 24954 4200 25230
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 3884 24268 3936 24274
rect 3884 24210 3936 24216
rect 3896 23730 3924 24210
rect 4080 23798 4108 24550
rect 4264 24154 4292 25230
rect 4356 24256 4384 25350
rect 4724 24614 4752 25452
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4356 24228 4476 24256
rect 4172 24126 4292 24154
rect 4344 24132 4396 24138
rect 4068 23792 4120 23798
rect 3988 23752 4068 23780
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 3988 23610 4016 23752
rect 4068 23734 4120 23740
rect 3896 23582 4016 23610
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 3896 22642 3924 23582
rect 3976 23520 4028 23526
rect 3976 23462 4028 23468
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3988 22234 4016 23462
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 4080 22094 4108 23598
rect 3896 22066 4108 22094
rect 3896 22012 3924 22066
rect 3804 21984 3924 22012
rect 3804 17882 3832 21984
rect 4172 21690 4200 24126
rect 4344 24074 4396 24080
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23866 4292 24006
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4264 22778 4292 23666
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 4356 22506 4384 24074
rect 4448 23662 4476 24228
rect 4436 23656 4488 23662
rect 4436 23598 4488 23604
rect 4816 23526 4844 25298
rect 4908 24614 4936 25774
rect 5000 25294 5028 26522
rect 5092 26450 5120 26726
rect 5170 26480 5226 26489
rect 5080 26444 5132 26450
rect 5170 26415 5226 26424
rect 5080 26386 5132 26392
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4908 24274 4936 24550
rect 5000 24410 5028 24686
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 4896 24268 4948 24274
rect 4896 24210 4948 24216
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4816 22642 4844 23462
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4264 22030 4292 22374
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4816 22216 4844 22578
rect 4908 22438 4936 24210
rect 4988 23656 5040 23662
rect 4988 23598 5040 23604
rect 5000 23118 5028 23598
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4724 22188 4844 22216
rect 4724 22030 4752 22188
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4804 22024 4856 22030
rect 5000 22012 5028 23054
rect 4856 21984 5028 22012
rect 4804 21966 4856 21972
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3988 20890 4016 21490
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4172 20942 4200 21422
rect 4264 21418 4292 21966
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4356 21554 4384 21626
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4252 21412 4304 21418
rect 4252 21354 4304 21360
rect 4160 20936 4212 20942
rect 4066 20904 4122 20913
rect 3988 20862 4066 20890
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3896 19854 3924 19926
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3896 18766 3924 19314
rect 3988 19174 4016 20862
rect 4160 20878 4212 20884
rect 4066 20839 4122 20848
rect 4172 20534 4200 20878
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 19922 4108 20198
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4172 19378 4200 20470
rect 4264 20330 4292 21354
rect 4356 20602 4384 21490
rect 4724 21332 4752 21966
rect 4816 21554 4844 21966
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4896 21480 4948 21486
rect 4894 21448 4896 21457
rect 4948 21448 4950 21457
rect 4894 21383 4950 21392
rect 4804 21344 4856 21350
rect 4724 21304 4804 21332
rect 4804 21286 4856 21292
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4632 20505 4660 20742
rect 4618 20496 4674 20505
rect 4724 20466 4752 20810
rect 4816 20466 4844 21286
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4618 20431 4674 20440
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4724 20369 4752 20402
rect 4710 20360 4766 20369
rect 4252 20324 4304 20330
rect 4710 20295 4766 20304
rect 4252 20266 4304 20272
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 4172 18902 4200 19314
rect 4264 18970 4292 20266
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 4172 17746 4200 18838
rect 4356 18290 4384 19790
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4436 19372 4488 19378
rect 4724 19360 4752 19722
rect 4816 19718 4844 20402
rect 4908 20398 4936 21082
rect 5000 20602 5028 21830
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4908 19802 4936 20334
rect 5092 19854 5120 26386
rect 5184 23662 5212 26415
rect 5368 26042 5396 27474
rect 5460 27470 5488 28630
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5552 27878 5580 28494
rect 5632 28212 5684 28218
rect 5632 28154 5684 28160
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5540 27328 5592 27334
rect 5644 27316 5672 28154
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5920 27402 5948 27814
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5592 27288 5672 27316
rect 6012 27282 6040 29038
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 6196 28558 6224 28902
rect 6380 28762 6408 29514
rect 6368 28756 6420 28762
rect 6368 28698 6420 28704
rect 6656 28558 6684 29990
rect 6932 29306 6960 30194
rect 7208 29510 7236 30194
rect 7656 29572 7708 29578
rect 7656 29514 7708 29520
rect 8300 29572 8352 29578
rect 8300 29514 8352 29520
rect 7196 29504 7248 29510
rect 7196 29446 7248 29452
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 6932 28558 6960 29242
rect 7208 29102 7236 29446
rect 7196 29096 7248 29102
rect 7196 29038 7248 29044
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6276 28416 6328 28422
rect 6276 28358 6328 28364
rect 6288 28218 6316 28358
rect 6276 28212 6328 28218
rect 6276 28154 6328 28160
rect 6564 27878 6592 28494
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6748 28218 6776 28358
rect 6736 28212 6788 28218
rect 6736 28154 6788 28160
rect 6932 28150 6960 28494
rect 7208 28404 7236 29038
rect 7576 28966 7604 29446
rect 7564 28960 7616 28966
rect 7564 28902 7616 28908
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7288 28416 7340 28422
rect 7208 28376 7288 28404
rect 7340 28376 7420 28404
rect 7288 28358 7340 28364
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6748 27878 6776 28018
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 5540 27270 5592 27276
rect 5552 27062 5580 27270
rect 5920 27254 6040 27282
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5552 26586 5580 26998
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5276 25498 5304 25638
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5368 25158 5396 25434
rect 5552 25294 5580 26522
rect 5920 26382 5948 27254
rect 6092 27056 6144 27062
rect 6012 27004 6092 27010
rect 6012 26998 6144 27004
rect 6012 26982 6132 26998
rect 6012 26858 6040 26982
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 6000 26852 6052 26858
rect 6000 26794 6052 26800
rect 6092 26852 6144 26858
rect 6092 26794 6144 26800
rect 6104 26586 6132 26794
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 6092 26580 6144 26586
rect 6092 26522 6144 26528
rect 6012 26466 6040 26522
rect 6012 26438 6224 26466
rect 6288 26450 6316 26862
rect 6368 26784 6420 26790
rect 6368 26726 6420 26732
rect 6196 26382 6224 26438
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 6380 26382 6408 26726
rect 6564 26382 6592 27814
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6748 26586 6776 27338
rect 6840 27130 6868 28018
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 6736 26580 6788 26586
rect 6736 26522 6788 26528
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6368 26376 6420 26382
rect 6552 26376 6604 26382
rect 6368 26318 6420 26324
rect 6472 26336 6552 26364
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5264 24880 5316 24886
rect 5264 24822 5316 24828
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5276 22250 5304 24822
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5460 24342 5488 24550
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5552 24206 5580 24550
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5368 23730 5396 24142
rect 5644 23798 5672 25230
rect 5736 23798 5764 25298
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5828 24818 5856 25094
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5724 23792 5776 23798
rect 5724 23734 5776 23740
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5368 22409 5396 22578
rect 5354 22400 5410 22409
rect 5354 22335 5410 22344
rect 5184 22222 5304 22250
rect 5184 21332 5212 22222
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 5276 21457 5304 21558
rect 5368 21486 5396 21830
rect 5460 21729 5488 23598
rect 5552 23497 5580 23598
rect 5538 23488 5594 23497
rect 5538 23423 5594 23432
rect 5644 23322 5672 23598
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5552 22778 5580 22918
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5736 22234 5764 23598
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5736 22094 5764 22170
rect 5644 22066 5764 22094
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5446 21720 5502 21729
rect 5446 21655 5448 21664
rect 5500 21655 5502 21664
rect 5448 21626 5500 21632
rect 5552 21593 5580 21966
rect 5538 21584 5594 21593
rect 5448 21548 5500 21554
rect 5538 21519 5540 21528
rect 5448 21490 5500 21496
rect 5592 21519 5594 21528
rect 5540 21490 5592 21496
rect 5356 21480 5408 21486
rect 5262 21448 5318 21457
rect 5356 21422 5408 21428
rect 5262 21383 5318 21392
rect 5184 21304 5396 21332
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5184 20602 5212 20878
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5276 19854 5304 20402
rect 5080 19848 5132 19854
rect 4908 19774 5028 19802
rect 5080 19790 5132 19796
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4908 19360 4936 19654
rect 5000 19496 5028 19774
rect 5276 19514 5304 19790
rect 5264 19508 5316 19514
rect 5000 19468 5212 19496
rect 5080 19372 5132 19378
rect 4488 19332 4844 19360
rect 4908 19332 5080 19360
rect 4436 19314 4488 19320
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4816 18426 4844 19332
rect 5080 19314 5132 19320
rect 5184 19242 5212 19468
rect 5264 19450 5316 19456
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4252 18080 4304 18086
rect 4448 18068 4476 18294
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4252 18022 4304 18028
rect 4356 18040 4476 18068
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4264 17678 4292 18022
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 3896 17338 3924 17614
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3568 16544 3740 16572
rect 3516 16526 3568 16532
rect 3804 16538 3832 17138
rect 4160 16584 4212 16590
rect 3804 16510 3924 16538
rect 4160 16526 4212 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16250 3832 16390
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2148 14822 2176 15846
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2148 14414 2176 14758
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 756 12232 808 12238
rect 756 12174 808 12180
rect 768 12073 796 12174
rect 2056 12102 2084 13466
rect 2148 12918 2176 14350
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2240 12238 2268 15438
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2516 13530 2544 14554
rect 2700 14278 2728 14758
rect 2884 14414 2912 14758
rect 3160 14618 3188 15982
rect 3344 15706 3372 16050
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3804 15502 3832 16050
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2700 14006 2728 14214
rect 2976 14074 3004 14214
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2884 13326 2912 13942
rect 3068 13938 3096 14282
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12238 2636 13126
rect 2884 12986 2912 13262
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3068 12434 3096 13874
rect 2976 12406 3096 12434
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2044 12096 2096 12102
rect 754 12064 810 12073
rect 2044 12038 2096 12044
rect 754 11999 810 12008
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10742 1900 10950
rect 1964 10810 1992 11494
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 756 10668 808 10674
rect 756 10610 808 10616
rect 768 10169 796 10610
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1872 10198 1900 10678
rect 1860 10192 1912 10198
rect 754 10160 810 10169
rect 1860 10134 1912 10140
rect 754 10095 810 10104
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1504 8974 1532 9590
rect 1596 9586 1624 9998
rect 1872 9722 1900 10134
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 9178 1992 9318
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2056 8974 2084 9590
rect 2148 9586 2176 11562
rect 2240 9674 2268 12174
rect 2608 11694 2636 12174
rect 2976 11762 3004 12406
rect 3252 12238 3280 15438
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3344 14618 3372 14962
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3436 14074 3464 14418
rect 3528 14074 3556 14894
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3344 12850 3372 13466
rect 3620 13258 3648 13874
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3344 12442 3372 12786
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11354 2544 11494
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2976 10810 3004 11698
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2240 9646 2544 9674
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2516 9450 2544 9646
rect 2700 9586 2728 10066
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1504 8634 1532 8910
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7274 1716 7686
rect 1780 7342 1808 7822
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 6730 1716 7210
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 754 6352 810 6361
rect 1688 6322 1716 6666
rect 1872 6458 1900 7822
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 754 6287 756 6296
rect 808 6287 810 6296
rect 1676 6316 1728 6322
rect 756 6258 808 6264
rect 1676 6258 1728 6264
rect 2148 4554 2176 9318
rect 2608 9178 2636 9318
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2792 8634 2820 9930
rect 3068 9926 3096 9998
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 9178 2912 9318
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3160 8634 3188 11018
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2332 7546 2360 7822
rect 2792 7546 2820 7822
rect 2884 7546 2912 7822
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 3160 6798 3188 8570
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2240 6458 2268 6734
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 3252 6322 3280 12174
rect 3528 11898 3556 12786
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3620 11830 3648 13194
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 8498 3464 9522
rect 3804 9450 3832 9998
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3608 9376 3660 9382
rect 3660 9336 3740 9364
rect 3608 9318 3660 9324
rect 3712 9042 3740 9336
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3804 8974 3832 9386
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3436 8090 3464 8434
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7546 3464 7822
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3804 7002 3832 7754
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3804 6186 3832 6938
rect 3896 6662 3924 16510
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16046 4016 16390
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3988 15434 4016 15982
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3976 14408 4028 14414
rect 4080 14396 4108 16186
rect 4172 15638 4200 16526
rect 4356 15994 4384 18040
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4816 17882 4844 18090
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4908 17678 4936 19110
rect 5184 18426 5212 19178
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4986 17912 5042 17921
rect 4986 17847 5042 17856
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4908 16590 4936 17070
rect 5000 16590 5028 17847
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4264 15966 4384 15994
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4172 14482 4200 15370
rect 4264 14550 4292 15966
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4356 15706 4384 15846
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4816 15706 4844 16390
rect 4908 16182 4936 16526
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 5000 15994 5028 16526
rect 4908 15966 5028 15994
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4618 15192 4674 15201
rect 4618 15127 4674 15136
rect 4632 15026 4660 15127
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4356 14618 4384 14962
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4028 14368 4108 14396
rect 3976 14350 4028 14356
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13326 4016 13670
rect 4264 13326 4292 14010
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4816 13394 4844 15030
rect 4908 14346 4936 15966
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5000 14550 5028 15438
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 5000 14074 5028 14486
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 3988 11762 4016 13262
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12986 4476 13126
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4172 11898 4200 12786
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4356 12434 4384 12582
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4816 12434 4844 13330
rect 5000 12714 5028 13806
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 4356 12406 4844 12434
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10742 4016 10950
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 4356 10674 4384 12406
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4908 9994 4936 11018
rect 5092 10742 5120 17478
rect 5184 16590 5212 17682
rect 5276 17678 5304 18226
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5368 17490 5396 21304
rect 5460 18358 5488 21490
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5552 21146 5580 21354
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5538 20360 5594 20369
rect 5538 20295 5594 20304
rect 5552 19718 5580 20295
rect 5644 19990 5672 22066
rect 5828 22030 5856 23802
rect 5920 22030 5948 26318
rect 6092 25764 6144 25770
rect 6092 25706 6144 25712
rect 6000 24336 6052 24342
rect 6000 24278 6052 24284
rect 6012 24138 6040 24278
rect 6104 24206 6132 25706
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 6012 23866 6040 24074
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6196 23746 6224 26318
rect 6472 26042 6500 26336
rect 6552 26318 6604 26324
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6472 24886 6500 25978
rect 6564 24954 6592 26182
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6656 25430 6684 25638
rect 6644 25424 6696 25430
rect 6644 25366 6696 25372
rect 6656 24954 6684 25366
rect 6552 24948 6604 24954
rect 6552 24890 6604 24896
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6460 24880 6512 24886
rect 6460 24822 6512 24828
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6288 24188 6316 24754
rect 6368 24200 6420 24206
rect 6288 24160 6368 24188
rect 6368 24142 6420 24148
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6012 23718 6224 23746
rect 6012 22778 6040 23718
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 6092 23044 6144 23050
rect 6092 22986 6144 22992
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5722 21720 5778 21729
rect 5722 21655 5778 21664
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5276 17462 5396 17490
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5276 16096 5304 17462
rect 5354 17368 5410 17377
rect 5552 17338 5580 19314
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 18057 5672 18226
rect 5630 18048 5686 18057
rect 5630 17983 5686 17992
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5354 17303 5356 17312
rect 5408 17303 5410 17312
rect 5540 17332 5592 17338
rect 5356 17274 5408 17280
rect 5540 17274 5592 17280
rect 5368 17218 5396 17274
rect 5368 17190 5580 17218
rect 5276 16068 5488 16096
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 14414 5212 15302
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5170 13696 5226 13705
rect 5170 13631 5226 13640
rect 5184 12986 5212 13631
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5184 10470 5212 11222
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10130 5212 10406
rect 5276 10266 5304 15914
rect 5354 15192 5410 15201
rect 5460 15162 5488 16068
rect 5354 15127 5410 15136
rect 5448 15156 5500 15162
rect 5368 14618 5396 15127
rect 5448 15098 5500 15104
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5460 13530 5488 15098
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 12238 5580 17190
rect 5644 16658 5672 17478
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5644 15162 5672 16594
rect 5736 15570 5764 21655
rect 5828 21434 5856 21966
rect 6012 21894 6040 22578
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5906 21584 5962 21593
rect 5906 21519 5908 21528
rect 5960 21519 5962 21528
rect 5908 21490 5960 21496
rect 5828 21418 5948 21434
rect 5828 21412 5960 21418
rect 5828 21406 5908 21412
rect 5828 20890 5856 21406
rect 5908 21354 5960 21360
rect 5828 20862 5948 20890
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5828 19922 5856 20742
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5920 19786 5948 20862
rect 6104 20602 6132 22986
rect 6196 22098 6224 23598
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6196 21622 6224 21898
rect 6184 21616 6236 21622
rect 6184 21558 6236 21564
rect 6196 20942 6224 21558
rect 6288 21146 6316 24006
rect 6380 23769 6408 24142
rect 6748 24070 6776 25910
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6840 24818 6868 25162
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6840 24274 6868 24754
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6748 23866 6776 24006
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6644 23792 6696 23798
rect 6366 23760 6422 23769
rect 6644 23734 6696 23740
rect 6366 23695 6422 23704
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6380 22166 6408 22714
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6368 22160 6420 22166
rect 6368 22102 6420 22108
rect 6368 22024 6420 22030
rect 6366 21992 6368 22001
rect 6420 21992 6422 22001
rect 6472 21962 6500 22374
rect 6366 21927 6422 21936
rect 6460 21956 6512 21962
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6196 20534 6224 20878
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5828 16250 5856 19654
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5920 17814 5948 18226
rect 6012 18222 6040 19926
rect 6104 19718 6132 20198
rect 6196 19990 6224 20334
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 6104 17270 6132 19654
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6196 18222 6224 18702
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5920 16114 5948 17002
rect 6012 16794 6040 17002
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6196 16454 6224 18158
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 16250 6224 16390
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5736 14414 5764 15302
rect 6012 15162 6040 15506
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6104 15026 6132 15914
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 6288 14006 6316 21082
rect 6380 20618 6408 21927
rect 6460 21898 6512 21904
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6472 21457 6500 21626
rect 6458 21448 6514 21457
rect 6458 21383 6514 21392
rect 6564 20806 6592 23462
rect 6656 23118 6684 23734
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6644 22228 6696 22234
rect 6748 22216 6776 23598
rect 6840 22982 6868 23666
rect 6932 23254 6960 27406
rect 7208 27402 7236 27814
rect 7196 27396 7248 27402
rect 7196 27338 7248 27344
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 7024 26586 7052 26726
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 7116 26489 7144 27066
rect 7392 26994 7420 28376
rect 7484 27656 7512 28494
rect 7576 27962 7604 28902
rect 7668 28762 7696 29514
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7656 28756 7708 28762
rect 7656 28698 7708 28704
rect 7760 28218 7788 28902
rect 8312 28490 8340 29514
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 7748 28212 7800 28218
rect 7748 28154 7800 28160
rect 8404 28150 8432 29038
rect 8484 28960 8536 28966
rect 8484 28902 8536 28908
rect 8852 28960 8904 28966
rect 8852 28902 8904 28908
rect 8496 28558 8524 28902
rect 8864 28558 8892 28902
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8852 28552 8904 28558
rect 8852 28494 8904 28500
rect 8392 28144 8444 28150
rect 8392 28086 8444 28092
rect 7576 27934 7696 27962
rect 7564 27668 7616 27674
rect 7484 27628 7564 27656
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7102 26480 7158 26489
rect 7102 26415 7158 26424
rect 7392 26353 7420 26930
rect 7378 26344 7434 26353
rect 7378 26279 7434 26288
rect 7484 26194 7512 27628
rect 7564 27610 7616 27616
rect 7668 26790 7696 27934
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 8300 26920 8352 26926
rect 8404 26908 8432 28086
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8496 27334 8524 27814
rect 8956 27606 8984 30670
rect 9416 30394 9444 30670
rect 9772 30660 9824 30666
rect 9772 30602 9824 30608
rect 9404 30388 9456 30394
rect 9404 30330 9456 30336
rect 9784 29646 9812 30602
rect 9876 30190 9904 30670
rect 9968 30258 9996 30806
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10060 30394 10088 30534
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 10244 30190 10272 30670
rect 9864 30184 9916 30190
rect 9864 30126 9916 30132
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9876 29578 9904 30126
rect 10336 29850 10364 31282
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10876 31136 10928 31142
rect 10876 31078 10928 31084
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 10428 30870 10456 31078
rect 10416 30864 10468 30870
rect 10416 30806 10468 30812
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10612 30258 10640 30670
rect 10888 30666 10916 31078
rect 11256 30802 11284 31078
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 12072 30864 12124 30870
rect 12072 30806 12124 30812
rect 25870 30832 25926 30841
rect 11244 30796 11296 30802
rect 11244 30738 11296 30744
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10612 29782 10640 30194
rect 10600 29776 10652 29782
rect 10600 29718 10652 29724
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 10704 29510 10732 30330
rect 12084 30190 12112 30806
rect 25870 30767 25926 30776
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 12176 30190 12204 30534
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 10980 29714 11008 30126
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 12084 29850 12112 30126
rect 12176 29850 12204 30126
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12164 29844 12216 29850
rect 12164 29786 12216 29792
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 10968 29708 11020 29714
rect 10968 29650 11020 29656
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 11164 29306 11192 29718
rect 12084 29306 12112 29786
rect 14648 29776 14700 29782
rect 14648 29718 14700 29724
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14372 29572 14424 29578
rect 14372 29514 14424 29520
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 12072 29300 12124 29306
rect 12072 29242 12124 29248
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 9692 28762 9720 29106
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 9048 28218 9076 28426
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9324 28218 9352 28358
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 9784 28150 9812 28494
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9876 28082 9904 28562
rect 10336 28558 10364 29106
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8496 26994 8524 27270
rect 8956 27062 8984 27542
rect 9324 27470 9352 27814
rect 9876 27674 9904 28018
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9312 27464 9364 27470
rect 9312 27406 9364 27412
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8352 26880 8432 26908
rect 8300 26862 8352 26868
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7668 26217 7696 26726
rect 7392 26166 7512 26194
rect 7654 26208 7710 26217
rect 7392 26081 7420 26166
rect 7654 26143 7710 26152
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7378 26072 7434 26081
rect 7896 26075 8204 26084
rect 7378 26007 7434 26016
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7288 25424 7340 25430
rect 7288 25366 7340 25372
rect 7300 25158 7328 25366
rect 7392 25294 7420 25842
rect 7484 25294 7512 25978
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 8024 25900 8076 25906
rect 8024 25842 8076 25848
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7576 25294 7604 25638
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7012 25152 7064 25158
rect 7288 25152 7340 25158
rect 7064 25112 7144 25140
rect 7012 25094 7064 25100
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7024 24206 7052 24754
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7024 23730 7052 24142
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6696 22188 6776 22216
rect 6644 22170 6696 22176
rect 6656 22030 6684 22170
rect 6840 22166 6868 22918
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 7024 22094 7052 22578
rect 6932 22066 7052 22094
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6828 21888 6880 21894
rect 6734 21856 6790 21865
rect 6828 21830 6880 21836
rect 6734 21791 6790 21800
rect 6748 21622 6776 21791
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6644 20936 6696 20942
rect 6696 20884 6776 20890
rect 6644 20878 6776 20884
rect 6656 20862 6776 20878
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6380 20590 6500 20618
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6380 19417 6408 20402
rect 6366 19408 6422 19417
rect 6366 19343 6422 19352
rect 6472 19360 6500 20590
rect 6564 20466 6592 20742
rect 6748 20466 6776 20862
rect 6840 20534 6868 21830
rect 6932 21350 6960 22066
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6748 19446 6776 20402
rect 6840 19514 6868 20470
rect 6932 20058 6960 20946
rect 7024 20777 7052 21898
rect 7116 21146 7144 25112
rect 7208 25112 7288 25140
rect 7208 24818 7236 25112
rect 7288 25094 7340 25100
rect 7392 24954 7420 25230
rect 7380 24948 7432 24954
rect 7380 24890 7432 24896
rect 7288 24880 7340 24886
rect 7288 24822 7340 24828
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24070 7236 24754
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23322 7236 24006
rect 7300 23798 7328 24822
rect 7392 24206 7420 24890
rect 7484 24818 7512 25230
rect 7564 25152 7616 25158
rect 7668 25140 7696 25638
rect 7760 25430 7788 25842
rect 7748 25424 7800 25430
rect 7748 25366 7800 25372
rect 7760 25294 7788 25366
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 8036 25158 8064 25842
rect 8220 25498 8248 25842
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 7616 25112 7696 25140
rect 7748 25152 7800 25158
rect 7564 25094 7616 25100
rect 7748 25094 7800 25100
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7576 24682 7604 25094
rect 7564 24676 7616 24682
rect 7564 24618 7616 24624
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7484 23730 7512 24142
rect 7576 23730 7604 24618
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7208 21486 7236 22578
rect 7300 21554 7328 23462
rect 7484 22778 7512 23530
rect 7576 22982 7604 23666
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21570 7420 21830
rect 7484 21690 7512 22374
rect 7668 22094 7696 24550
rect 7760 23730 7788 25094
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 8312 23848 8340 26862
rect 8496 25838 8524 26930
rect 9140 26926 9168 27270
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9140 26246 9168 26862
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9232 26314 9260 26726
rect 9416 26314 9444 26862
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9508 26314 9536 26726
rect 9968 26586 9996 28018
rect 10336 27538 10364 28494
rect 10612 28218 10640 28494
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10428 26994 10456 27610
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10704 27130 10732 27406
rect 11716 27334 11744 28358
rect 12452 27470 12480 29106
rect 13556 28762 13584 29106
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 14108 28558 14136 29446
rect 14384 28762 14412 29514
rect 14476 29306 14504 29582
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14568 28694 14596 28902
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 12808 28076 12860 28082
rect 12808 28018 12860 28024
rect 12624 27872 12676 27878
rect 12624 27814 12676 27820
rect 12636 27470 12664 27814
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 12452 27062 12480 27406
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 11072 26450 11100 26726
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11992 26586 12020 26930
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9128 26240 9180 26246
rect 9128 26182 9180 26188
rect 8484 25832 8536 25838
rect 8484 25774 8536 25780
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 8404 25226 8432 25366
rect 8496 25294 8524 25774
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9048 25362 9076 25638
rect 9036 25356 9088 25362
rect 9036 25298 9088 25304
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 8496 24732 8524 25230
rect 8588 24886 8616 25230
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 8864 24750 8892 24822
rect 9048 24818 9076 25298
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8576 24744 8628 24750
rect 8496 24704 8576 24732
rect 8576 24686 8628 24692
rect 8852 24744 8904 24750
rect 8852 24686 8904 24692
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8220 23820 8340 23848
rect 7748 23724 7800 23730
rect 7800 23684 7880 23712
rect 7748 23666 7800 23672
rect 7852 23526 7880 23684
rect 8220 23594 8248 23820
rect 8392 23724 8444 23730
rect 8312 23684 8392 23712
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7760 23118 7788 23462
rect 7852 23118 7880 23462
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7760 22710 7788 23054
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7576 22066 7696 22094
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7472 21582 7524 21588
rect 7288 21548 7340 21554
rect 7392 21542 7472 21570
rect 7472 21524 7524 21530
rect 7288 21490 7340 21496
rect 7576 21486 7604 22066
rect 7654 21720 7710 21729
rect 7654 21655 7710 21664
rect 7196 21480 7248 21486
rect 7564 21480 7616 21486
rect 7196 21422 7248 21428
rect 7470 21448 7526 21457
rect 7208 21146 7236 21422
rect 7564 21422 7616 21428
rect 7470 21383 7526 21392
rect 7286 21312 7342 21321
rect 7286 21247 7342 21256
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7010 20768 7066 20777
rect 7010 20703 7066 20712
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6552 19372 6604 19378
rect 6472 19332 6552 19360
rect 6552 19314 6604 19320
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6380 17610 6408 18158
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 12782 6132 13670
rect 6288 13530 6316 13942
rect 6472 13870 6500 19178
rect 6564 18193 6592 19314
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6748 18290 6776 18634
rect 6932 18426 6960 19654
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18766 7052 19110
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6550 18184 6606 18193
rect 6550 18119 6606 18128
rect 6932 17202 6960 18362
rect 7116 17678 7144 20538
rect 7300 18970 7328 21247
rect 7484 20942 7512 21383
rect 7668 21350 7696 21655
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 20466 7420 20742
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7484 18329 7512 20402
rect 7576 20040 7604 21286
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20262 7696 20878
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7656 20052 7708 20058
rect 7576 20012 7656 20040
rect 7656 19994 7708 20000
rect 7668 19310 7696 19994
rect 7760 19854 7788 22170
rect 8036 22166 8064 22578
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 8036 22001 8064 22102
rect 8220 22030 8248 22578
rect 8312 22234 8340 23684
rect 8392 23666 8444 23672
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8404 22778 8432 23190
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8496 22642 8524 23258
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8392 22568 8444 22574
rect 8444 22516 8524 22522
rect 8392 22510 8524 22516
rect 8404 22494 8524 22510
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8208 22024 8260 22030
rect 8022 21992 8078 22001
rect 8208 21966 8260 21972
rect 8022 21927 8078 21936
rect 8220 21876 8248 21966
rect 8220 21848 8340 21876
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 8312 21622 8340 21848
rect 8496 21690 8524 22494
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8482 21584 8538 21593
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 7840 20528 7892 20534
rect 7838 20496 7840 20505
rect 7892 20496 7894 20505
rect 7838 20431 7894 20440
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7852 19700 7880 20431
rect 8312 19990 8340 21558
rect 8482 21519 8484 21528
rect 8536 21519 8538 21528
rect 8484 21490 8536 21496
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8404 20058 8432 21422
rect 8496 20398 8524 21490
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8484 19916 8536 19922
rect 8588 19904 8616 24006
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8680 22982 8708 23462
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 8680 22166 8708 22442
rect 8668 22160 8720 22166
rect 8668 22102 8720 22108
rect 8666 21448 8722 21457
rect 8666 21383 8722 21392
rect 8536 19876 8616 19904
rect 8484 19858 8536 19864
rect 7760 19672 7880 19700
rect 8392 19712 8444 19718
rect 7760 19496 7788 19672
rect 8392 19654 8444 19660
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 8404 19514 8432 19654
rect 8392 19508 8444 19514
rect 7760 19468 7972 19496
rect 7944 19378 7972 19468
rect 8392 19450 8444 19456
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7470 18320 7526 18329
rect 7470 18255 7526 18264
rect 7668 17814 7696 19246
rect 7760 18766 7788 19314
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7760 18290 7788 18702
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17814 8616 18022
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6748 15978 6776 16390
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6104 12434 6132 12718
rect 6196 12646 6224 13262
rect 6288 12850 6316 13466
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6656 12918 6684 13126
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6012 12406 6132 12434
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11354 5672 11698
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5736 11150 5764 11494
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5644 10198 5672 10406
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4158 9616 4214 9625
rect 4158 9551 4214 9560
rect 4172 8566 4200 9551
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 5736 9178 5764 9998
rect 5828 9654 5856 10134
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5920 9586 5948 10542
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5920 9042 5948 9522
rect 6012 9500 6040 12406
rect 6196 12322 6224 12582
rect 6380 12434 6408 12718
rect 6380 12406 6500 12434
rect 6196 12306 6408 12322
rect 6196 12300 6420 12306
rect 6196 12294 6368 12300
rect 6368 12242 6420 12248
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6472 11150 6500 12406
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11354 6868 11494
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10674 6500 11086
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6196 10266 6224 10610
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6092 9512 6144 9518
rect 6012 9472 6092 9500
rect 6092 9454 6144 9460
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6564 8974 6592 9318
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8634 5488 8774
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4816 8090 4844 8366
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 8242 5396 8298
rect 5632 8288 5684 8294
rect 5368 8214 5580 8242
rect 5632 8230 5684 8236
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7546 4476 7686
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4816 7342 4844 8026
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 7546 4936 7754
rect 5552 7546 5580 8214
rect 5644 7818 5672 8230
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4816 6882 4844 7278
rect 4724 6854 4844 6882
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 4724 6458 4752 6854
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4724 6254 4752 6394
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 756 4548 808 4554
rect 756 4490 808 4496
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 768 4457 796 4490
rect 754 4448 810 4457
rect 754 4383 810 4392
rect 4080 3942 4108 6054
rect 4264 5778 4292 6190
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 5370 4200 5646
rect 4816 5370 4844 6258
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4078 4844 4762
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 5276 3602 5304 5170
rect 5552 4622 5580 7482
rect 5736 7478 5764 8230
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5828 7206 5856 8842
rect 6656 8634 6684 9386
rect 6748 8634 6776 9522
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6644 7948 6696 7954
rect 6564 7908 6644 7936
rect 6564 7546 6592 7908
rect 6644 7890 6696 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6458 6132 7142
rect 6656 6730 6684 7754
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7546 6776 7686
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 6458 6592 6598
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5644 5166 5672 5850
rect 6656 5710 6684 6666
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5914 6776 6054
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5302 6684 5646
rect 6840 5302 6868 8230
rect 7024 7002 7052 17138
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16561 7144 16934
rect 7380 16584 7432 16590
rect 7102 16552 7158 16561
rect 7380 16526 7432 16532
rect 7102 16487 7158 16496
rect 7116 16114 7144 16487
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 16250 7236 16390
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7392 15978 7420 16526
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7668 16250 7696 16458
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14414 7144 14894
rect 7392 14414 7420 15302
rect 7760 15162 7788 17206
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 8312 15162 8340 15302
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8128 14482 8156 14894
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7116 13394 7144 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 12986 7696 13194
rect 7760 12986 7788 13670
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8312 12646 8340 13670
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 11830 7420 12242
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10742 7144 10950
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7300 10266 7328 11086
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7392 9994 7420 11766
rect 8496 11642 8524 14214
rect 8588 12434 8616 17614
rect 8680 17202 8708 21383
rect 8772 21146 8800 24142
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8864 21078 8892 24686
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8852 21072 8904 21078
rect 8852 21014 8904 21020
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8772 20058 8800 20810
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8864 17746 8892 20810
rect 8956 19446 8984 23462
rect 9048 23186 9076 24074
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22574 9076 22918
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9048 20058 9076 22510
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 21457 9168 22442
rect 9126 21448 9182 21457
rect 9126 21383 9182 21392
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9140 21146 9168 21286
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9232 20942 9260 26250
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9324 24886 9352 25230
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9324 23798 9352 24210
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9324 22778 9352 23734
rect 9416 23526 9444 26250
rect 10600 26240 10652 26246
rect 10652 26200 10732 26228
rect 10600 26182 10652 26188
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10336 25888 10364 25978
rect 10416 25900 10468 25906
rect 10336 25860 10416 25888
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9508 23322 9536 24754
rect 9600 24410 9628 25230
rect 9784 24614 9812 25774
rect 10336 25294 10364 25860
rect 10416 25842 10468 25848
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10428 25498 10456 25638
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10612 25430 10640 25774
rect 10600 25424 10652 25430
rect 10600 25366 10652 25372
rect 10612 25294 10640 25366
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 10324 25288 10376 25294
rect 10600 25288 10652 25294
rect 10376 25248 10456 25276
rect 10324 25230 10376 25236
rect 9876 24954 9904 25230
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 10324 24880 10376 24886
rect 10324 24822 10376 24828
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9232 19922 9260 20198
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 18290 9076 19314
rect 9232 18766 9260 19858
rect 9324 19514 9352 22034
rect 9404 21684 9456 21690
rect 9456 21644 9536 21672
rect 9404 21626 9456 21632
rect 9508 21078 9536 21644
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9416 20466 9444 20946
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9508 19378 9536 21014
rect 9600 20942 9628 21422
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 19378 9628 20742
rect 9692 19514 9720 22986
rect 9784 21690 9812 24550
rect 9968 24206 9996 24550
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23186 9904 24074
rect 9968 23254 9996 24142
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 10060 23118 10088 23666
rect 10152 23118 10180 23734
rect 10244 23322 10272 24754
rect 10336 24206 10364 24822
rect 10428 24818 10456 25248
rect 10600 25230 10652 25236
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10508 24812 10560 24818
rect 10612 24800 10640 25230
rect 10560 24772 10640 24800
rect 10508 24754 10560 24760
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23866 10364 24142
rect 10428 24070 10456 24754
rect 10416 24064 10468 24070
rect 10416 24006 10468 24012
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10324 23656 10376 23662
rect 10324 23598 10376 23604
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10336 23118 10364 23598
rect 10520 23322 10548 24754
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9876 21418 9904 21558
rect 9968 21554 9996 21898
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9784 20806 9812 21354
rect 9876 21078 9904 21354
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 20800 9824 20806
rect 9824 20760 9904 20788
rect 9772 20742 9824 20748
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9784 19786 9812 20266
rect 9876 20058 9904 20760
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9864 19848 9916 19854
rect 9862 19816 9864 19825
rect 9916 19816 9918 19825
rect 9772 19780 9824 19786
rect 9862 19751 9918 19760
rect 9772 19722 9824 19728
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 18970 9628 19178
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18306 9260 18702
rect 9324 18426 9352 18838
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9508 18426 9536 18702
rect 9692 18426 9720 18702
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9128 18284 9180 18290
rect 9232 18278 9444 18306
rect 9128 18226 9180 18232
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 17082 8708 17138
rect 8680 17054 8800 17082
rect 9140 17066 9168 18226
rect 9416 18222 9444 18278
rect 9496 18284 9548 18290
rect 9548 18244 9812 18272
rect 9496 18226 9548 18232
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17814 9444 18158
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17814 9720 18022
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16182 8708 16934
rect 8772 16522 8800 17054
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9140 16794 9168 17002
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9416 16726 9444 17614
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 8760 16516 8812 16522
rect 8760 16458 8812 16464
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8772 14006 8800 16458
rect 9416 16250 9444 16662
rect 9692 16658 9720 17750
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9508 15706 9536 16390
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9324 15366 9352 15506
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9232 14414 9260 15302
rect 9416 15162 9444 15438
rect 9784 15314 9812 18244
rect 9876 16794 9904 19654
rect 9968 19514 9996 21490
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10060 18834 10088 23054
rect 10704 22094 10732 26200
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10980 25498 11008 25638
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 11256 25294 11284 25978
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10796 24342 10824 24822
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 10784 24336 10836 24342
rect 10784 24278 10836 24284
rect 11808 24274 11836 25230
rect 11900 24954 11928 25230
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10888 23866 10916 24142
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10888 23254 10916 23462
rect 10876 23248 10928 23254
rect 10876 23190 10928 23196
rect 10980 23186 11008 23734
rect 11256 23322 11284 24074
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10612 22066 10732 22094
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10324 20052 10376 20058
rect 10152 20012 10324 20040
rect 10152 19718 10180 20012
rect 10324 19994 10376 20000
rect 10324 19916 10376 19922
rect 10244 19876 10324 19904
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10140 19168 10192 19174
rect 10244 19156 10272 19876
rect 10324 19858 10376 19864
rect 10322 19816 10378 19825
rect 10428 19802 10456 21898
rect 10612 19854 10640 22066
rect 10888 22030 10916 22510
rect 10980 22234 11008 23122
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11532 22778 11560 22918
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11624 22658 11652 22918
rect 11716 22778 11744 24210
rect 11900 24206 11928 24754
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11164 22630 11652 22658
rect 11888 22636 11940 22642
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10980 21690 11008 21966
rect 11072 21894 11100 21966
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 20942 10824 21286
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10378 19774 10456 19802
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10322 19751 10378 19760
rect 10192 19128 10272 19156
rect 10140 19110 10192 19116
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18358 9996 18702
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 10060 18465 10088 18634
rect 10046 18456 10102 18465
rect 10046 18391 10102 18400
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 10046 18320 10102 18329
rect 9968 17542 9996 18294
rect 10046 18255 10048 18264
rect 10100 18255 10102 18264
rect 10048 18226 10100 18232
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9968 16590 9996 16934
rect 10244 16726 10272 19128
rect 10336 17882 10364 19751
rect 10690 19408 10746 19417
rect 10612 19366 10690 19394
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10428 18766 10456 19246
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9876 15706 9904 16050
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9784 15286 9996 15314
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9232 13530 9260 13738
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8588 12406 8800 12434
rect 8496 11626 8708 11642
rect 8496 11620 8720 11626
rect 8496 11614 8668 11620
rect 8668 11562 8720 11568
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11150 7696 11494
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 8680 10674 8708 11562
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7760 10418 7788 10474
rect 7668 10390 7788 10418
rect 7668 10198 7696 10390
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7576 7410 7604 8434
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7668 6882 7696 10134
rect 8772 10062 8800 12406
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10742 8892 11086
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8634 7788 9522
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8974 7972 9318
rect 8772 9178 8800 9590
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 8772 8634 8800 9114
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8496 7886 8524 8366
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 7002 7788 7142
rect 8036 7002 8064 7346
rect 8220 7206 8248 7414
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7668 6854 7788 6882
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7024 5370 7052 5578
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4214 5672 4422
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5828 3738 5856 4558
rect 6840 4282 6868 5238
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4758 7328 5170
rect 7484 5030 7512 5510
rect 7668 5370 7696 5510
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7300 4554 7328 4694
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4282 6960 4422
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7668 4146 7696 4762
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 6564 3534 6592 3878
rect 7668 3738 7696 4082
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 6656 2514 6684 3674
rect 7760 2650 7788 6854
rect 8404 6798 8432 7142
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8496 6458 8524 6734
rect 8588 6730 8616 8366
rect 8864 8090 8892 8502
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8496 5914 8524 6394
rect 8588 6322 8616 6666
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8588 5234 8616 6258
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8956 4826 8984 13262
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12850 9168 13194
rect 9324 12986 9352 14758
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 12986 9444 13670
rect 9692 13462 9720 13874
rect 9784 13802 9812 14350
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9508 12782 9536 13262
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9588 13184 9640 13190
rect 9640 13144 9720 13172
rect 9588 13126 9640 13132
rect 9692 12866 9720 13144
rect 9784 12986 9812 13194
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9692 12838 9904 12866
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9048 11218 9076 11562
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9036 10804 9088 10810
rect 9088 10764 9168 10792
rect 9036 10746 9088 10752
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 8496 4282 8524 4558
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 9048 4146 9076 9930
rect 9140 8906 9168 10764
rect 9232 10266 9260 12582
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9324 10606 9352 11154
rect 9600 11150 9628 12038
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 9772 11348 9824 11354
rect 9692 11286 9720 11319
rect 9772 11290 9824 11296
rect 9680 11280 9732 11286
rect 9784 11257 9812 11290
rect 9680 11222 9732 11228
rect 9770 11248 9826 11257
rect 9876 11218 9904 12838
rect 9770 11183 9826 11192
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 10810 9628 11086
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10266 9352 10406
rect 9508 10266 9536 10678
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 8634 9168 8842
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9232 6866 9260 9998
rect 9600 9994 9628 10746
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9692 9382 9720 10950
rect 9968 10810 9996 15286
rect 10048 14952 10100 14958
rect 10046 14920 10048 14929
rect 10100 14920 10102 14929
rect 10046 14855 10102 14864
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 13938 10364 14214
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10428 13190 10456 18566
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10520 15706 10548 17614
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10060 11898 10088 13126
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9680 9376 9732 9382
rect 9732 9336 9812 9364
rect 9680 9318 9732 9324
rect 9600 9178 9628 9318
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9324 6746 9352 8570
rect 9692 8566 9720 8842
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9232 6730 9352 6746
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9220 6724 9352 6730
rect 9272 6718 9352 6724
rect 9220 6666 9272 6672
rect 9140 5642 9168 6666
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9232 5030 9260 5646
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 7944 3738 7972 4082
rect 9232 3942 9260 4966
rect 9324 4282 9352 6718
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9784 6338 9812 9336
rect 9876 9178 9904 9522
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9862 9072 9918 9081
rect 9862 9007 9864 9016
rect 9916 9007 9918 9016
rect 9956 9036 10008 9042
rect 9864 8978 9916 8984
rect 9956 8978 10008 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8430 9904 8842
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9968 8294 9996 8978
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8022 9996 8230
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 6458 9904 7278
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9784 6322 9904 6338
rect 9784 6316 9916 6322
rect 9784 6310 9864 6316
rect 9864 6258 9916 6264
rect 9876 5914 9904 6258
rect 9968 5914 9996 6734
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 4622 9720 5714
rect 9784 5658 9812 5782
rect 9784 5630 9904 5658
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9784 4690 9812 5102
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9312 4140 9364 4146
rect 9416 4128 9444 4490
rect 9364 4100 9444 4128
rect 9312 4082 9364 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 9600 3466 9628 4490
rect 9784 4214 9812 4490
rect 9876 4214 9904 5630
rect 10060 5234 10088 6666
rect 10152 5846 10180 11290
rect 10612 11218 10640 19366
rect 10690 19343 10746 19352
rect 10796 17882 10824 20878
rect 11072 20806 11100 21490
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10888 20058 10916 20402
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10980 19922 11008 20198
rect 11072 20058 11100 20402
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11072 19514 11100 19994
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10980 19174 11008 19382
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10888 16998 10916 19110
rect 10980 18834 11008 19110
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11164 18698 11192 22630
rect 11888 22578 11940 22584
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11256 21962 11284 22510
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11716 22234 11744 22510
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11624 21894 11652 22102
rect 11808 22030 11836 22510
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 20602 11284 20878
rect 11716 20874 11744 21966
rect 11808 21350 11836 21966
rect 11900 21894 11928 22578
rect 11992 22234 12020 22578
rect 12084 22438 12112 23462
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 21486 11928 21830
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 12084 21010 12112 22374
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 11794 20904 11850 20913
rect 11704 20868 11756 20874
rect 11794 20839 11850 20848
rect 11704 20810 11756 20816
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11716 20058 11744 20810
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11348 19514 11376 19790
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11428 19440 11480 19446
rect 11426 19408 11428 19417
rect 11480 19408 11482 19417
rect 11244 19372 11296 19378
rect 11808 19360 11836 20839
rect 11426 19343 11482 19352
rect 11244 19314 11296 19320
rect 11716 19332 11836 19360
rect 11256 19174 11284 19314
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11256 18426 11284 19110
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11716 17814 11744 19332
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11808 18970 11836 19178
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 12176 18426 12204 26318
rect 12452 25362 12480 26998
rect 12820 26586 12848 28018
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13636 27396 13688 27402
rect 13636 27338 13688 27344
rect 13176 27328 13228 27334
rect 13176 27270 13228 27276
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12912 25906 12940 26862
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 26586 13124 26726
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13188 26518 13216 27270
rect 13648 26518 13676 27338
rect 13924 27130 13952 27814
rect 14568 27470 14596 28630
rect 14660 28098 14688 29718
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14752 28762 14780 29514
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 15488 29170 15516 29446
rect 15672 29306 15700 29990
rect 15856 29850 15884 30194
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15752 29776 15804 29782
rect 15752 29718 15804 29724
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 15304 28558 15332 28902
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 15212 28218 15240 28358
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 14660 28070 15056 28098
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 13912 27124 13964 27130
rect 13912 27066 13964 27072
rect 13176 26512 13228 26518
rect 13176 26454 13228 26460
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 14464 26444 14516 26450
rect 14464 26386 14516 26392
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12360 24818 12388 25230
rect 12452 24818 12480 25298
rect 12820 25294 12848 25638
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12912 25140 12940 25842
rect 12820 25112 12940 25140
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12360 24206 12388 24754
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12820 23730 12848 25112
rect 12992 24812 13044 24818
rect 12992 24754 13044 24760
rect 13004 23866 13032 24754
rect 13096 24138 13124 26250
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 13280 26042 13308 26182
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12820 23633 12848 23666
rect 12806 23624 12862 23633
rect 12806 23559 12862 23568
rect 13004 23050 13032 23802
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12912 22778 12940 22986
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12256 22432 12308 22438
rect 12360 22420 12388 22578
rect 12308 22392 12388 22420
rect 12256 22374 12308 22380
rect 12268 22234 12296 22374
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12544 21962 12572 22578
rect 12728 22409 12756 22578
rect 13096 22438 13124 24074
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13176 22500 13228 22506
rect 13176 22442 13228 22448
rect 13084 22432 13136 22438
rect 12714 22400 12770 22409
rect 13084 22374 13136 22380
rect 12714 22335 12770 22344
rect 13188 22094 13216 22442
rect 13096 22066 13216 22094
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12544 21690 12572 21898
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12820 21554 12848 21966
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12360 18290 12388 19110
rect 12452 18834 12480 19110
rect 12544 18902 12572 21422
rect 12820 21078 12848 21490
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12636 18290 12664 19314
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11716 17270 11744 17750
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14074 10732 14962
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10690 11384 10746 11393
rect 10690 11319 10692 11328
rect 10744 11319 10746 11328
rect 10692 11290 10744 11296
rect 10600 11212 10652 11218
rect 10428 11172 10600 11200
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10674 10272 10950
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 9178 10364 10406
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8634 10272 9046
rect 10428 8634 10456 11172
rect 10600 11154 10652 11160
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10810 10548 10950
rect 10796 10810 10824 16594
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16250 11008 16458
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14414 10916 14758
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10980 12986 11008 15438
rect 11072 13444 11100 15506
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11164 15162 11192 15370
rect 11256 15162 11284 15846
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11164 14006 11192 14894
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11716 14278 11744 14962
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11152 13456 11204 13462
rect 11072 13416 11152 13444
rect 11072 13326 11100 13416
rect 11152 13398 11204 13404
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11624 13326 11652 13359
rect 11716 13326 11744 14214
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 10674 10916 12582
rect 11072 11150 11100 13126
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10612 9625 10640 10610
rect 11060 10600 11112 10606
rect 11058 10568 11060 10577
rect 11112 10568 11114 10577
rect 11058 10503 11114 10512
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 9722 10916 10406
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10598 9616 10654 9625
rect 10598 9551 10600 9560
rect 10652 9551 10654 9560
rect 10600 9522 10652 9528
rect 10980 9382 11008 9930
rect 10692 9376 10744 9382
rect 10968 9376 11020 9382
rect 10692 9318 10744 9324
rect 10796 9336 10968 9364
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10598 9072 10654 9081
rect 10520 8838 10548 9046
rect 10598 9007 10654 9016
rect 10612 8974 10640 9007
rect 10600 8968 10652 8974
rect 10704 8945 10732 9318
rect 10600 8910 10652 8916
rect 10690 8936 10746 8945
rect 10690 8871 10692 8880
rect 10744 8871 10746 8880
rect 10692 8842 10744 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10612 8566 10640 8774
rect 10796 8566 10824 9336
rect 10968 9318 11020 9324
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10232 7948 10284 7954
rect 10284 7908 10456 7936
rect 10232 7890 10284 7896
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 7002 10272 7346
rect 10428 7002 10456 7908
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10520 6798 10548 7686
rect 10612 7410 10640 7686
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 6452 10560 6458
rect 10612 6440 10640 7346
rect 10560 6412 10640 6440
rect 10508 6394 10560 6400
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10140 5840 10192 5846
rect 10428 5794 10456 6054
rect 10140 5782 10192 5788
rect 10244 5766 10456 5794
rect 10520 5778 10548 6394
rect 10244 5710 10272 5766
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 5370 10364 5646
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10428 5302 10456 5766
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 4826 10088 5170
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9692 3534 9720 4014
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6656 1970 6684 2450
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7208 2106 7236 2314
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 8496 2038 8524 2790
rect 9692 2582 9720 3062
rect 9784 2582 9812 4014
rect 9968 3720 9996 4558
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4214 10180 4422
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10520 4146 10548 5714
rect 10888 5166 10916 8570
rect 10966 8528 11022 8537
rect 11072 8498 11100 8774
rect 10966 8463 10968 8472
rect 11020 8463 11022 8472
rect 11060 8492 11112 8498
rect 10968 8434 11020 8440
rect 11060 8434 11112 8440
rect 11164 8362 11192 13262
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11256 12714 11284 13194
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12782 11376 13126
rect 11440 12850 11468 13262
rect 11808 12850 11836 17478
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11808 11830 11836 12786
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11900 11762 11928 18226
rect 11992 16794 12020 18226
rect 12636 17882 12664 18226
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17338 12204 17546
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12084 17241 12112 17274
rect 12070 17232 12126 17241
rect 12070 17167 12126 17176
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12268 17105 12296 17138
rect 12254 17096 12310 17105
rect 12254 17031 12310 17040
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16454 12020 16526
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 14890 12020 16390
rect 12084 16250 12112 16662
rect 12268 16658 12296 16934
rect 12544 16794 12572 17138
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12728 16590 12756 19110
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11992 12986 12020 13874
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12176 12866 12204 16050
rect 12452 15706 12480 16390
rect 12728 16250 12756 16526
rect 12820 16522 12848 18226
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12820 16114 12848 16458
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12438 15192 12494 15201
rect 12438 15127 12440 15136
rect 12492 15127 12494 15136
rect 12440 15098 12492 15104
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12256 13388 12308 13394
rect 12308 13348 12480 13376
rect 12256 13330 12308 13336
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 11992 12838 12204 12866
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 11992 12306 12020 12838
rect 12164 12640 12216 12646
rect 12084 12600 12164 12628
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11348 10742 11376 11222
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11716 10674 11744 11562
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11900 10690 11928 10746
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11808 10662 11928 10690
rect 11256 10266 11284 10610
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11256 8430 11284 9522
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7546 11008 8230
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11072 6866 11100 7958
rect 11716 7834 11744 8434
rect 11808 7970 11836 10662
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 8106 11928 10474
rect 11992 10198 12020 10950
rect 12084 10588 12112 12600
rect 12164 12582 12216 12588
rect 12162 12336 12218 12345
rect 12162 12271 12218 12280
rect 12176 11898 12204 12271
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 10690 12204 11698
rect 12268 10810 12296 12854
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12176 10662 12296 10690
rect 12360 10674 12388 13126
rect 12452 12714 12480 13348
rect 12544 13326 12572 14010
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12452 11370 12480 12650
rect 12452 11354 12572 11370
rect 12452 11348 12584 11354
rect 12452 11342 12532 11348
rect 12532 11290 12584 11296
rect 12084 10560 12204 10588
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 9518 12112 9930
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11992 8838 12020 9386
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8650 12020 8774
rect 11992 8622 12112 8650
rect 12084 8566 12112 8622
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12176 8362 12204 10560
rect 12268 9178 12296 10662
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12452 8974 12480 9862
rect 12544 9586 12572 11290
rect 12728 10690 12756 15642
rect 12912 15570 12940 21286
rect 12990 20904 13046 20913
rect 12990 20839 13046 20848
rect 13004 20806 13032 20839
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 20534 13032 20742
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 13004 19854 13032 20470
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19378 13032 19790
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13004 18426 13032 18566
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13096 17542 13124 22066
rect 13372 22030 13400 22578
rect 13360 22024 13412 22030
rect 13174 21992 13230 22001
rect 13360 21966 13412 21972
rect 13174 21927 13176 21936
rect 13228 21927 13230 21936
rect 13176 21898 13228 21904
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 13188 21146 13216 21490
rect 13648 21350 13676 25094
rect 13924 24342 13952 25094
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23866 13768 24006
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13924 23322 13952 24278
rect 14476 24138 14504 26386
rect 14660 25242 14688 27950
rect 14922 27568 14978 27577
rect 14922 27503 14978 27512
rect 14936 27470 14964 27503
rect 15028 27470 15056 28070
rect 15304 27606 15332 28494
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15212 27470 15240 27542
rect 15304 27470 15332 27542
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 14752 27130 14780 27406
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14832 26784 14884 26790
rect 14752 26732 14832 26738
rect 14752 26726 14884 26732
rect 14752 26710 14872 26726
rect 14752 25430 14780 26710
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14740 25424 14792 25430
rect 14740 25366 14792 25372
rect 14568 25214 14688 25242
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13360 20868 13412 20874
rect 13360 20810 13412 20816
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13280 20466 13308 20538
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13188 18698 13216 20402
rect 13280 19854 13308 20402
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 18766 13308 19790
rect 13372 19174 13400 20810
rect 13556 20777 13584 20878
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14004 20800 14056 20806
rect 13542 20768 13598 20777
rect 14096 20800 14148 20806
rect 14004 20742 14056 20748
rect 14094 20768 14096 20777
rect 14148 20768 14150 20777
rect 13542 20703 13598 20712
rect 14016 20466 14044 20742
rect 14094 20703 14150 20712
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 13452 20392 13504 20398
rect 13636 20392 13688 20398
rect 13504 20352 13636 20380
rect 13452 20334 13504 20340
rect 13636 20334 13688 20340
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18970 13400 19110
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13372 18766 13400 18906
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13542 18728 13598 18737
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13174 18456 13230 18465
rect 13174 18391 13230 18400
rect 13188 18154 13216 18391
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17814 13216 18090
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13280 17746 13308 18702
rect 13542 18663 13598 18672
rect 13556 18630 13584 18663
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 17740 13320 17746
rect 13320 17700 13400 17728
rect 13268 17682 13320 17688
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13188 16114 13216 17546
rect 13266 17232 13322 17241
rect 13372 17202 13400 17700
rect 13266 17167 13268 17176
rect 13320 17167 13322 17176
rect 13360 17196 13412 17202
rect 13268 17138 13320 17144
rect 13360 17138 13412 17144
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15638 13124 15846
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 15162 12940 15302
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14414 12848 14758
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 12850 13032 14282
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12820 12753 12848 12786
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 13096 12442 13124 12786
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 10810 12848 11698
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11150 13032 11494
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12728 10662 12848 10690
rect 13188 10674 13216 14214
rect 13280 13326 13308 16458
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 9110 12572 9318
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 11900 8078 12204 8106
rect 11808 7942 11928 7970
rect 11624 7806 11744 7834
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11624 7546 11652 7806
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11256 6934 11284 7482
rect 11716 7426 11744 7686
rect 11624 7410 11744 7426
rect 11612 7404 11744 7410
rect 11664 7398 11744 7404
rect 11612 7346 11664 7352
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11808 7002 11836 7822
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 5794 11100 6802
rect 11900 6254 11928 7942
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11072 5766 11192 5794
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 11164 4690 11192 5766
rect 11900 5710 11928 6190
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11716 4758 11744 5578
rect 11992 5302 12020 5782
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4486 11100 4558
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11164 4214 11192 4626
rect 11992 4622 12020 4966
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11624 4214 11652 4422
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 9876 3692 9996 3720
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9048 2106 9076 2314
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 4423 1660 4731 1669
rect 4423 1658 4429 1660
rect 4485 1658 4509 1660
rect 4565 1658 4589 1660
rect 4645 1658 4669 1660
rect 4725 1658 4731 1660
rect 4485 1606 4487 1658
rect 4667 1606 4669 1658
rect 4423 1604 4429 1606
rect 4485 1604 4509 1606
rect 4565 1604 4589 1606
rect 4645 1604 4669 1606
rect 4725 1604 4731 1606
rect 4423 1595 4731 1604
rect 7944 1426 7972 1838
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 9508 1358 9536 2246
rect 9692 2038 9720 2518
rect 9784 2106 9812 2518
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9876 1834 9904 3692
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9968 1970 9996 3470
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3126 10088 3334
rect 10244 3194 10272 3402
rect 10336 3194 10364 3878
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10796 3194 10824 3878
rect 11256 3398 11284 3878
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 11256 2514 11284 3334
rect 11624 3058 11652 3674
rect 11716 3534 11744 4422
rect 12084 4196 12112 5646
rect 11900 4168 12112 4196
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 11808 2666 11836 2790
rect 11716 2638 11836 2666
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10060 2106 10088 2382
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10244 2038 10272 2246
rect 11256 2038 11284 2450
rect 11716 2446 11744 2638
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 10232 2032 10284 2038
rect 10232 1974 10284 1980
rect 11244 2032 11296 2038
rect 11244 1974 11296 1980
rect 9956 1964 10008 1970
rect 9956 1906 10008 1912
rect 11900 1834 11928 4168
rect 12176 3738 12204 8078
rect 12268 7818 12296 8298
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12452 6458 12480 7822
rect 12544 7478 12572 7890
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12360 5710 12388 6258
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12348 5364 12400 5370
rect 12452 5352 12480 6258
rect 12636 5914 12664 10542
rect 12820 10146 12848 10662
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13004 10266 13032 10610
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12728 10118 12848 10146
rect 12728 9081 12756 10118
rect 13188 9654 13216 10610
rect 13372 10062 13400 15506
rect 13464 13802 13492 18022
rect 13648 15706 13676 20334
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13832 19854 13860 20266
rect 14108 20058 14136 20402
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19378 13768 19722
rect 13832 19378 13860 19790
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13740 17241 13768 18702
rect 13832 17882 13860 18770
rect 14108 18766 14136 19858
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14200 18766 14228 19790
rect 14292 19174 14320 20266
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14188 18760 14240 18766
rect 14240 18720 14320 18748
rect 14188 18702 14240 18708
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18290 13952 18566
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13726 17232 13782 17241
rect 13726 17167 13728 17176
rect 13780 17167 13782 17176
rect 13728 17138 13780 17144
rect 13818 16144 13874 16153
rect 13818 16079 13874 16088
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13832 15434 13860 16079
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 15094 13860 15370
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13556 13938 13584 14554
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14090 13860 14214
rect 13740 14062 13860 14090
rect 13740 13938 13768 14062
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 13832 12850 13860 13874
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12306 13860 12786
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10674 13676 11154
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13176 9648 13228 9654
rect 13452 9648 13504 9654
rect 13176 9590 13228 9596
rect 13450 9616 13452 9625
rect 13504 9616 13506 9625
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12900 9580 12952 9586
rect 13450 9551 13506 9560
rect 12900 9522 12952 9528
rect 12714 9072 12770 9081
rect 12820 9042 12848 9522
rect 12912 9178 12940 9522
rect 13358 9480 13414 9489
rect 13358 9415 13414 9424
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12714 9007 12770 9016
rect 12808 9036 12860 9042
rect 12728 8838 12756 9007
rect 12808 8978 12860 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8362 12756 8774
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 13096 8090 13124 8842
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12728 7546 12756 7890
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7546 12848 7686
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12716 6384 12768 6390
rect 12768 6344 12848 6372
rect 12716 6326 12768 6332
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5710 12572 5782
rect 12532 5704 12584 5710
rect 12530 5672 12532 5681
rect 12584 5672 12586 5681
rect 12530 5607 12586 5616
rect 12400 5324 12480 5352
rect 12348 5306 12400 5312
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12636 5098 12664 5238
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12728 4758 12756 6054
rect 12820 5681 12848 6344
rect 12912 6118 12940 7822
rect 13004 7546 13032 7822
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13004 6322 13032 7346
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 13188 5914 13216 8978
rect 13280 8945 13308 8978
rect 13372 8974 13400 9415
rect 13360 8968 13412 8974
rect 13266 8936 13322 8945
rect 13360 8910 13412 8916
rect 13266 8871 13322 8880
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8430 13400 8774
rect 13464 8498 13492 9551
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 7886 13400 8366
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13360 7472 13412 7478
rect 13450 7440 13506 7449
rect 13412 7420 13450 7426
rect 13360 7414 13450 7420
rect 13372 7398 13450 7414
rect 13450 7375 13506 7384
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12900 5704 12952 5710
rect 12806 5672 12862 5681
rect 12900 5646 12952 5652
rect 12806 5607 12862 5616
rect 12912 5370 12940 5646
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12268 4214 12296 4490
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 2650 12020 3334
rect 12268 3058 12296 4150
rect 12544 3738 12572 4150
rect 12728 3738 12756 4694
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12820 3534 12848 4422
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3738 12940 4082
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 13280 2650 13308 7142
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5914 13400 6054
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13450 4720 13506 4729
rect 13450 4655 13506 4664
rect 13464 4282 13492 4655
rect 13556 4622 13584 10610
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13648 7410 13676 8298
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 6458 13676 7346
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13648 5030 13676 6394
rect 13740 5914 13768 11222
rect 13832 11082 13860 11562
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13924 8974 13952 18226
rect 14016 17610 14044 18702
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 18193 14228 18226
rect 14186 18184 14242 18193
rect 14186 18119 14242 18128
rect 14292 17814 14320 18720
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 14016 16250 14044 17546
rect 14292 17338 14320 17750
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14108 17105 14136 17206
rect 14188 17128 14240 17134
rect 14094 17096 14150 17105
rect 14188 17070 14240 17076
rect 14094 17031 14150 17040
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13832 6730 13860 7754
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 6798 13952 7142
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 14016 6474 14044 14962
rect 14108 9466 14136 17031
rect 14200 16726 14228 17070
rect 14188 16720 14240 16726
rect 14384 16674 14412 20810
rect 14188 16662 14240 16668
rect 14292 16646 14412 16674
rect 14292 16454 14320 16646
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14200 16250 14228 16390
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14292 15502 14320 16118
rect 14384 15706 14412 16526
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14384 14346 14412 14418
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14200 14006 14228 14282
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14200 13530 14228 13942
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14292 13433 14320 13874
rect 14278 13424 14334 13433
rect 14278 13359 14334 13368
rect 14384 13326 14412 14282
rect 14476 14278 14504 23462
rect 14568 21486 14596 25214
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14660 24886 14688 25094
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14660 23118 14688 24074
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14752 22438 14780 25366
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 15212 23100 15240 27406
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15304 27130 15332 27270
rect 15396 27130 15424 28494
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15488 27010 15516 29106
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 27470 15608 27814
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15396 26982 15516 27010
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15304 23798 15332 24006
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15396 23118 15424 26982
rect 15580 25838 15608 27270
rect 15672 26994 15700 28018
rect 15764 27470 15792 29718
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 17960 29572 18012 29578
rect 17960 29514 18012 29520
rect 16500 29238 16528 29514
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 16120 27464 16172 27470
rect 16172 27412 16252 27418
rect 16120 27406 16252 27412
rect 16132 27390 16252 27406
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 15660 26988 15712 26994
rect 15712 26948 15884 26976
rect 15660 26930 15712 26936
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15488 25294 15516 25638
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15580 25140 15608 25774
rect 15672 25294 15700 26182
rect 15764 26042 15792 26318
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15752 25764 15804 25770
rect 15752 25706 15804 25712
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15580 25112 15700 25140
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24410 15516 24550
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23322 15516 24006
rect 15580 23798 15608 24210
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15292 23112 15344 23118
rect 15212 23072 15292 23100
rect 15292 23054 15344 23060
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 21622 14688 21830
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14568 19718 14596 21422
rect 14752 21146 14780 21966
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14844 21078 14872 21286
rect 15212 21146 15240 22918
rect 15304 22234 15332 23054
rect 15488 22778 15516 23054
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15396 22094 15424 22510
rect 15304 22066 15424 22094
rect 15304 21894 15332 22066
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14844 20942 14872 21014
rect 15488 20942 15516 22578
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20534 14688 20810
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14752 20466 14780 20742
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 15212 20534 15240 20742
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14648 19848 14700 19854
rect 14936 19825 14964 20198
rect 14648 19790 14700 19796
rect 14922 19816 14978 19825
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 17746 14596 19654
rect 14660 19310 14688 19790
rect 14922 19751 14978 19760
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14660 18630 14688 19246
rect 14752 18766 14780 19450
rect 15212 19446 15240 20470
rect 15580 20398 15608 23734
rect 15672 22574 15700 25112
rect 15764 24410 15792 25706
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15764 22030 15792 22646
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15672 20466 15700 21558
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 20058 15424 20198
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15474 19408 15530 19417
rect 15474 19343 15476 19352
rect 15528 19343 15530 19352
rect 15476 19314 15528 19320
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 15120 18714 15148 19110
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14660 18358 14688 18566
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14660 17338 14688 18294
rect 14752 18086 14780 18702
rect 15120 18686 15240 18714
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 15212 18408 15240 18686
rect 15304 18578 15332 19178
rect 15396 18698 15424 19246
rect 15488 18766 15516 19314
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15476 18624 15528 18630
rect 15304 18572 15476 18578
rect 15304 18566 15528 18572
rect 15304 18550 15516 18566
rect 15120 18380 15240 18408
rect 15382 18456 15438 18465
rect 15382 18391 15438 18400
rect 15120 18290 15148 18380
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 15434 14596 16390
rect 14660 16130 14688 16662
rect 14752 16250 14780 17614
rect 14844 17542 14872 18158
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 15212 17338 15240 18226
rect 15396 18154 15424 18391
rect 15488 18222 15516 18550
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14660 16102 14780 16130
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14568 15162 14596 15370
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14464 14272 14516 14278
rect 14660 14226 14688 15982
rect 14752 14521 14780 16102
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15028 15638 15056 15846
rect 15120 15638 15148 16050
rect 15016 15632 15068 15638
rect 14922 15600 14978 15609
rect 15016 15574 15068 15580
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 14922 15535 14978 15544
rect 14936 15502 14964 15535
rect 15304 15518 15332 18022
rect 15580 17954 15608 19722
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15672 18086 15700 18702
rect 15764 18630 15792 21966
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15752 18284 15804 18290
rect 15856 18272 15884 26948
rect 16040 26353 16068 27270
rect 16132 26790 16160 27270
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16026 26344 16082 26353
rect 16026 26279 16082 26288
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15948 25226 15976 25978
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15948 24750 15976 25162
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 16132 24614 16160 26726
rect 16224 25702 16252 27390
rect 16316 25770 16344 28970
rect 16500 28966 16528 29174
rect 17408 29028 17460 29034
rect 17408 28970 17460 28976
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 17132 28960 17184 28966
rect 17132 28902 17184 28908
rect 17224 28960 17276 28966
rect 17224 28902 17276 28908
rect 17144 28762 17172 28902
rect 17132 28756 17184 28762
rect 17132 28698 17184 28704
rect 17236 28558 17264 28902
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17420 27606 17448 28970
rect 17972 28694 18000 29514
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18064 28762 18092 29106
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18052 28756 18104 28762
rect 18052 28698 18104 28704
rect 17960 28688 18012 28694
rect 17960 28630 18012 28636
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 28218 18092 28358
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16500 26994 16528 27270
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 16592 26586 16620 27338
rect 16868 26976 16896 27338
rect 17420 27062 17448 27542
rect 17512 27130 17540 27814
rect 18156 27674 18184 28494
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 17684 27396 17736 27402
rect 17684 27338 17736 27344
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 16948 26988 17000 26994
rect 16868 26948 16948 26976
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16304 25764 16356 25770
rect 16304 25706 16356 25712
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 25226 16252 25638
rect 16776 25498 16804 26454
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 23866 16160 24550
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 23520 16080 23526
rect 15948 23480 16028 23508
rect 15948 18358 15976 23480
rect 16028 23462 16080 23468
rect 16132 23118 16160 23598
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 22574 16160 23054
rect 16396 22976 16448 22982
rect 16394 22944 16396 22953
rect 16448 22944 16450 22953
rect 16394 22879 16450 22888
rect 16120 22568 16172 22574
rect 16040 22528 16120 22556
rect 16040 22098 16068 22528
rect 16120 22510 16172 22516
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 16040 20856 16068 22034
rect 16304 21888 16356 21894
rect 16592 21876 16620 24754
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16684 22137 16712 23598
rect 16776 22778 16804 25434
rect 16868 24818 16896 26948
rect 16948 26930 17000 26936
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24886 16988 25094
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16868 23186 16896 23530
rect 17052 23202 17080 26726
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17144 24818 17172 26318
rect 17236 26042 17264 26318
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17328 25770 17356 26522
rect 17696 25974 17724 27338
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 18064 26382 18092 26862
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18064 25974 18092 26318
rect 17684 25968 17736 25974
rect 17684 25910 17736 25916
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18800 25838 18828 29582
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20824 29306 20852 29446
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 19708 29164 19760 29170
rect 19708 29106 19760 29112
rect 19064 29028 19116 29034
rect 19064 28970 19116 28976
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18892 28558 18920 28902
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 18892 28014 18920 28494
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18892 26926 18920 27950
rect 18984 27674 19012 28018
rect 18972 27668 19024 27674
rect 18972 27610 19024 27616
rect 19076 26976 19104 28970
rect 19156 28484 19208 28490
rect 19156 28426 19208 28432
rect 19168 28218 19196 28426
rect 19720 28218 19748 29106
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 20628 28416 20680 28422
rect 20628 28358 20680 28364
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19892 28076 19944 28082
rect 19892 28018 19944 28024
rect 19904 27674 19932 28018
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 20640 27606 20668 28358
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20732 27674 20760 28086
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 20720 27668 20772 27674
rect 20720 27610 20772 27616
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19156 26988 19208 26994
rect 19076 26948 19156 26976
rect 19156 26930 19208 26936
rect 18880 26920 18932 26926
rect 18880 26862 18932 26868
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18984 26450 19012 26726
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18788 25832 18840 25838
rect 18788 25774 18840 25780
rect 17316 25764 17368 25770
rect 17316 25706 17368 25712
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17144 23662 17172 24550
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16960 23174 17080 23202
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16670 22128 16726 22137
rect 16960 22094 16988 23174
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22438 17080 23054
rect 17236 22964 17264 24550
rect 17328 23202 17356 25706
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18800 25362 18828 25774
rect 18892 25498 18920 25842
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17420 24206 17448 25162
rect 17788 24954 17816 25162
rect 17776 24948 17828 24954
rect 17776 24890 17828 24896
rect 17880 24818 17908 25162
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 17972 24954 18000 25094
rect 17960 24948 18012 24954
rect 17960 24890 18012 24896
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17328 23174 17448 23202
rect 17420 23118 17448 23174
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17144 22936 17264 22964
rect 17408 22976 17460 22982
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16670 22063 16726 22072
rect 16868 22066 16988 22094
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16356 21848 16620 21876
rect 16304 21830 16356 21836
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16120 20868 16172 20874
rect 16040 20828 16120 20856
rect 16120 20810 16172 20816
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 16040 19446 16068 19722
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15804 18244 15884 18272
rect 15752 18226 15804 18232
rect 15660 18080 15712 18086
rect 15764 18057 15792 18226
rect 15948 18086 15976 18294
rect 16040 18222 16068 18566
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15936 18080 15988 18086
rect 15660 18022 15712 18028
rect 15750 18048 15806 18057
rect 15936 18022 15988 18028
rect 15750 17983 15806 17992
rect 15580 17926 15700 17954
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 17338 15424 17546
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15476 16040 15528 16046
rect 15528 15988 15608 15994
rect 15476 15982 15608 15988
rect 15488 15966 15608 15982
rect 15580 15910 15608 15966
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15292 15512 15344 15518
rect 14924 15496 14976 15502
rect 15292 15454 15344 15460
rect 14924 15438 14976 15444
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14738 14512 14794 14521
rect 14738 14447 14794 14456
rect 14464 14214 14516 14220
rect 14568 14198 14688 14226
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13462 14504 13670
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12442 14412 12582
rect 14372 12436 14424 12442
rect 14568 12434 14596 14198
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12986 14688 13126
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14752 12714 14780 13806
rect 14844 13258 14872 13874
rect 15028 13530 15056 13874
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15212 13326 15240 14214
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14568 12406 14780 12434
rect 14372 12378 14424 12384
rect 14370 12336 14426 12345
rect 14370 12271 14426 12280
rect 14384 12238 14412 12271
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11898 14228 12038
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14200 11218 14228 11834
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14200 9586 14228 11154
rect 14384 11082 14412 11630
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14476 11257 14504 11290
rect 14462 11248 14518 11257
rect 14660 11218 14688 12106
rect 14462 11183 14518 11192
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10266 14320 10610
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14476 9722 14504 10134
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14108 9438 14412 9466
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14200 9110 14228 9318
rect 14292 9178 14320 9318
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14096 7880 14148 7886
rect 14148 7840 14320 7868
rect 14096 7822 14148 7828
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 7002 14228 7346
rect 14292 7342 14320 7840
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14292 6882 14320 7278
rect 14384 6916 14412 9438
rect 14476 8974 14504 9522
rect 14568 9382 14596 10950
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14568 8480 14596 9046
rect 14660 8634 14688 9454
rect 14752 9178 14780 12406
rect 15304 12306 15332 15454
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15108 12164 15160 12170
rect 15160 12124 15240 12152
rect 15108 12106 15160 12112
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 15212 10742 15240 12124
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15304 10146 15332 11766
rect 15396 10266 15424 15846
rect 15488 15337 15516 15846
rect 15672 15722 15700 17926
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15580 15694 15700 15722
rect 15580 15473 15608 15694
rect 15566 15464 15622 15473
rect 15566 15399 15622 15408
rect 15568 15360 15620 15366
rect 15474 15328 15530 15337
rect 15568 15302 15620 15308
rect 15474 15263 15530 15272
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15488 13938 15516 14554
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15304 10118 15424 10146
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 15292 9648 15344 9654
rect 15290 9616 15292 9625
rect 15344 9616 15346 9625
rect 15290 9551 15346 9560
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8634 14780 8774
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 8492 14700 8498
rect 14568 8452 14648 8480
rect 14648 8434 14700 8440
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 8090 14504 8230
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 14740 6928 14792 6934
rect 14384 6888 14740 6916
rect 14200 6854 14320 6882
rect 14740 6870 14792 6876
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13924 6446 14044 6474
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3670 13584 3878
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 11992 1970 12020 2586
rect 13464 2378 13492 2790
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 13464 2038 13492 2314
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 13648 1970 13676 3334
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 12164 1964 12216 1970
rect 12164 1906 12216 1912
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 11888 1828 11940 1834
rect 11888 1770 11940 1776
rect 9876 1562 9904 1770
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11369 1660 11677 1669
rect 11369 1658 11375 1660
rect 11431 1658 11455 1660
rect 11511 1658 11535 1660
rect 11591 1658 11615 1660
rect 11671 1658 11677 1660
rect 11431 1606 11433 1658
rect 11613 1606 11615 1658
rect 11369 1604 11375 1606
rect 11431 1604 11455 1606
rect 11511 1604 11535 1606
rect 11591 1604 11615 1606
rect 11671 1604 11677 1606
rect 11369 1595 11677 1604
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 11992 1358 12020 1702
rect 12176 1562 12204 1906
rect 13740 1766 13768 5646
rect 13924 4554 13952 6446
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14016 4690 14044 6326
rect 14108 5710 14136 6734
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14096 5568 14148 5574
rect 14200 5556 14228 6854
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6390 14504 6598
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14292 5914 14320 6190
rect 14568 6186 14780 6202
rect 14568 6180 14792 6186
rect 14568 6174 14740 6180
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14280 5568 14332 5574
rect 14200 5528 14280 5556
rect 14096 5510 14148 5516
rect 14280 5510 14332 5516
rect 14108 5302 14136 5510
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14292 5234 14320 5510
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 5012 14320 5170
rect 14384 5166 14412 5782
rect 14568 5370 14596 6174
rect 14740 6122 14792 6128
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14660 5234 14688 6054
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14752 5370 14780 5578
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14292 4984 14412 5012
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 14016 3602 14044 4626
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14108 4214 14136 4422
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14292 3738 14320 4558
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14384 2774 14412 4984
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 15212 4146 15240 9114
rect 15304 8294 15332 9114
rect 15396 8906 15424 10118
rect 15488 8906 15516 12174
rect 15580 10266 15608 15302
rect 15764 15162 15792 16934
rect 15856 15416 15884 17818
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15948 15706 15976 16186
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15948 15609 15976 15642
rect 15934 15600 15990 15609
rect 15934 15535 15990 15544
rect 15936 15428 15988 15434
rect 15856 15388 15936 15416
rect 15936 15370 15988 15376
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15764 13530 15792 14826
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15842 12880 15898 12889
rect 15948 12850 15976 14010
rect 15842 12815 15898 12824
rect 15936 12844 15988 12850
rect 15856 12442 15884 12815
rect 15936 12786 15988 12792
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 16040 12102 16068 18158
rect 16132 16250 16160 19654
rect 16224 18714 16252 20470
rect 16316 20262 16344 21490
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16304 19236 16356 19242
rect 16304 19178 16356 19184
rect 16316 18970 16344 19178
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16224 18686 16344 18714
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16224 17678 16252 18566
rect 16316 18222 16344 18686
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16316 17746 16344 18158
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15638 16160 16050
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16118 15464 16174 15473
rect 16118 15399 16174 15408
rect 16132 15366 16160 15399
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16132 11830 16160 15302
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16224 11234 16252 17614
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 16114 16344 17478
rect 16408 16114 16436 21848
rect 16684 21690 16712 21898
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16670 21584 16726 21593
rect 16670 21519 16726 21528
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 20942 16620 21286
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16500 20602 16528 20810
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16316 11830 16344 15506
rect 16394 14512 16450 14521
rect 16394 14447 16396 14456
rect 16448 14447 16450 14456
rect 16396 14418 16448 14424
rect 16394 14376 16450 14385
rect 16394 14311 16450 14320
rect 16408 13938 16436 14311
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16500 12850 16528 20198
rect 16592 17882 16620 20878
rect 16684 19310 16712 21519
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 20058 16804 20742
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16684 17762 16712 19246
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18426 16804 18566
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17882 16804 18022
rect 16868 17882 16896 22066
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16960 18290 16988 21966
rect 17052 20346 17080 22374
rect 17144 21298 17172 22936
rect 17408 22918 17460 22924
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17236 21554 17264 22714
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17144 21270 17264 21298
rect 17236 20466 17264 21270
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17316 20392 17368 20398
rect 17052 20318 17264 20346
rect 17316 20334 17368 20340
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17052 18630 17080 20198
rect 17144 19922 17172 20198
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 18358 17172 18566
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16684 17734 17172 17762
rect 16580 17672 16632 17678
rect 16632 17620 16804 17626
rect 16580 17614 16804 17620
rect 16592 17598 16804 17614
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16590 16620 17478
rect 16580 16584 16632 16590
rect 16672 16584 16724 16590
rect 16580 16526 16632 16532
rect 16670 16552 16672 16561
rect 16724 16552 16726 16561
rect 16670 16487 16726 16496
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 13705 16620 14758
rect 16672 13728 16724 13734
rect 16578 13696 16634 13705
rect 16672 13670 16724 13676
rect 16578 13631 16634 13640
rect 16684 13530 16712 13670
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16592 12714 16620 13126
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16500 12374 16528 12650
rect 16684 12646 16712 13262
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16304 11824 16356 11830
rect 16356 11784 16436 11812
rect 16304 11766 16356 11772
rect 16132 11206 16252 11234
rect 15936 11144 15988 11150
rect 15750 11112 15806 11121
rect 15936 11086 15988 11092
rect 15750 11047 15806 11056
rect 15764 11014 15792 11047
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15764 10538 15792 10950
rect 15856 10674 15884 10950
rect 15844 10668 15896 10674
rect 15948 10656 15976 11086
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16040 10810 16068 11018
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15948 10628 16068 10656
rect 15844 10610 15896 10616
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15568 10260 15620 10266
rect 15764 10248 15792 10474
rect 15844 10260 15896 10266
rect 15764 10220 15844 10248
rect 15568 10202 15620 10208
rect 15844 10202 15896 10208
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15476 8900 15528 8906
rect 15528 8860 15608 8888
rect 15476 8842 15528 8848
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7546 15332 8230
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15396 7426 15424 8842
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15304 7398 15424 7426
rect 15304 5681 15332 7398
rect 15488 6866 15516 7686
rect 15580 7478 15608 8860
rect 15856 8838 15884 9998
rect 15948 9178 15976 9998
rect 16040 9382 16068 10628
rect 16132 10062 16160 11206
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10810 16252 11018
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 9722 16160 9998
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15936 8560 15988 8566
rect 15658 8528 15714 8537
rect 16040 8537 16068 9114
rect 16132 9024 16160 9522
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16224 9178 16252 9454
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16132 8996 16252 9024
rect 16118 8936 16174 8945
rect 16118 8871 16174 8880
rect 16132 8838 16160 8871
rect 16120 8832 16172 8838
rect 16224 8809 16252 8996
rect 16120 8774 16172 8780
rect 16210 8800 16266 8809
rect 15936 8502 15988 8508
rect 16026 8528 16082 8537
rect 15658 8463 15714 8472
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15672 5846 15700 8463
rect 15842 8256 15898 8265
rect 15842 8191 15898 8200
rect 15856 8090 15884 8191
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15384 5704 15436 5710
rect 15290 5672 15346 5681
rect 15384 5646 15436 5652
rect 15290 5607 15346 5616
rect 15396 5370 15424 5646
rect 15948 5370 15976 8502
rect 16026 8463 16082 8472
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15488 4214 15516 4422
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14752 2990 14780 4014
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 15212 3194 15240 4082
rect 15672 3738 15700 4558
rect 15856 4214 15884 4966
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15856 3670 15884 4150
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14384 2746 14504 2774
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 12164 1556 12216 1562
rect 12164 1498 12216 1504
rect 14384 1358 14412 2246
rect 14476 1902 14504 2746
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14752 1358 14780 2926
rect 15396 2650 15424 2994
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15856 2446 15884 3334
rect 16040 3126 16068 8230
rect 16132 6390 16160 8774
rect 16210 8735 16266 8744
rect 16224 8430 16252 8735
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 8090 16252 8230
rect 16316 8090 16344 10610
rect 16408 8634 16436 11784
rect 16776 11150 16804 17598
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16868 16697 16896 16730
rect 16854 16688 16910 16697
rect 16854 16623 16910 16632
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16868 10810 16896 16458
rect 16960 15502 16988 17546
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17052 15706 17080 16186
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16960 13802 16988 15302
rect 17144 14929 17172 17734
rect 17236 16454 17264 20318
rect 17328 20058 17356 20334
rect 17420 20262 17448 22918
rect 17512 21894 17540 24754
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17604 23866 17632 24074
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17788 21962 17816 22578
rect 17880 22094 17908 24754
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18156 22574 18184 22918
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 17880 22066 18000 22094
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17972 21894 18000 22066
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17512 21146 17540 21830
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17328 18737 17356 19654
rect 17512 19514 17540 19790
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17420 18766 17448 19110
rect 17408 18760 17460 18766
rect 17314 18728 17370 18737
rect 17408 18702 17460 18708
rect 17314 18663 17370 18672
rect 17328 18358 17356 18663
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17316 18352 17368 18358
rect 17420 18329 17448 18362
rect 17316 18294 17368 18300
rect 17406 18320 17462 18329
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17236 14260 17264 15370
rect 17328 15178 17356 18294
rect 17406 18255 17462 18264
rect 17406 18184 17462 18193
rect 17406 18119 17462 18128
rect 17420 15994 17448 18119
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17512 16153 17540 16458
rect 17498 16144 17554 16153
rect 17498 16079 17554 16088
rect 17420 15966 17540 15994
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15366 17448 15846
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17328 15150 17448 15178
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14618 17356 14962
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17316 14272 17368 14278
rect 17236 14232 17316 14260
rect 17316 14214 17368 14220
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16948 12640 17000 12646
rect 16946 12608 16948 12617
rect 17000 12608 17002 12617
rect 16946 12543 17002 12552
rect 17052 12442 17080 13806
rect 17328 13802 17356 14214
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17132 13184 17184 13190
rect 17236 13161 17264 13738
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17328 13433 17356 13466
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17420 13308 17448 15150
rect 17512 13818 17540 15966
rect 17604 15706 17632 21830
rect 17972 21690 18000 21830
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17696 21185 17724 21490
rect 17682 21176 17738 21185
rect 17682 21111 17738 21120
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17696 15706 17724 20742
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17788 19446 17816 19654
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17788 17202 17816 18022
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16454 17816 17138
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17604 14550 17632 15370
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17788 14890 17816 15098
rect 17880 14958 17908 20402
rect 17972 20058 18000 20538
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17972 19854 18000 19994
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17972 18834 18000 19382
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18290 18000 18770
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17972 16674 18000 17138
rect 18064 16794 18092 22374
rect 18156 21350 18184 22510
rect 18616 22420 18644 22986
rect 18708 22642 18736 23462
rect 18800 23322 18828 24074
rect 18892 23526 18920 25094
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18984 24410 19012 24754
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19168 24154 19196 26930
rect 19444 26314 19472 27338
rect 19628 27062 19656 27406
rect 19800 27396 19852 27402
rect 19800 27338 19852 27344
rect 20444 27396 20496 27402
rect 20444 27338 20496 27344
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19708 26988 19760 26994
rect 19708 26930 19760 26936
rect 19720 26586 19748 26930
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19260 24750 19288 25298
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19260 24274 19288 24686
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19168 24126 19288 24154
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18972 23248 19024 23254
rect 18892 23208 18972 23236
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18800 22438 18828 22918
rect 18892 22556 18920 23208
rect 18972 23190 19024 23196
rect 18972 22976 19024 22982
rect 19260 22930 19288 24126
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 19352 23322 19380 23530
rect 19444 23322 19472 26250
rect 19812 25702 19840 27338
rect 20456 26790 20484 27338
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19340 23112 19392 23118
rect 19392 23072 19472 23100
rect 19340 23054 19392 23060
rect 19444 22982 19472 23072
rect 18972 22918 19024 22924
rect 18984 22710 19012 22918
rect 19076 22902 19288 22930
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 18972 22568 19024 22574
rect 18892 22528 18972 22556
rect 18972 22510 19024 22516
rect 18788 22432 18840 22438
rect 18616 22392 18736 22420
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18708 22250 18736 22392
rect 18788 22374 18840 22380
rect 18708 22222 18828 22250
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18340 21486 18368 21898
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18156 20534 18184 21286
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18708 21146 18736 22102
rect 18800 22012 18828 22222
rect 18880 22024 18932 22030
rect 18800 21984 18880 22012
rect 18880 21966 18932 21972
rect 18892 21350 18920 21966
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18708 20874 18736 21082
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18156 19446 18184 20470
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18708 19854 18736 20402
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18248 19446 18276 19790
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18340 19334 18368 19654
rect 18248 19306 18368 19334
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17972 16646 18092 16674
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17696 14482 17724 14826
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17604 13938 17632 14214
rect 17788 14074 17816 14214
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17880 13818 17908 14418
rect 17972 14074 18000 16458
rect 18064 15638 18092 16646
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18064 14618 18092 15098
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17512 13790 17632 13818
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13394 17540 13670
rect 17604 13530 17632 13790
rect 17788 13790 17908 13818
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17682 13696 17738 13705
rect 17682 13631 17738 13640
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17696 13326 17724 13631
rect 17328 13280 17448 13308
rect 17684 13320 17736 13326
rect 17328 13190 17356 13280
rect 17684 13262 17736 13268
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17316 13184 17368 13190
rect 17132 13126 17184 13132
rect 17222 13152 17278 13161
rect 17144 12850 17172 13126
rect 17316 13126 17368 13132
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17222 13087 17278 13096
rect 17328 12986 17356 13126
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17328 12714 17356 12922
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17144 11694 17172 12650
rect 17420 12306 17448 13126
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16960 10742 16988 10950
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9722 16620 10066
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16592 8566 16620 8842
rect 16488 8560 16540 8566
rect 16486 8528 16488 8537
rect 16580 8560 16632 8566
rect 16540 8528 16542 8537
rect 16580 8502 16632 8508
rect 16486 8463 16542 8472
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7274 16252 7686
rect 16316 7546 16344 7822
rect 16408 7546 16436 8366
rect 16684 8106 16712 9114
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16500 8078 16712 8106
rect 16500 7886 16528 8078
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16394 7304 16450 7313
rect 16212 7268 16264 7274
rect 16394 7239 16450 7248
rect 16212 7210 16264 7216
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16132 6186 16160 6326
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16408 6118 16436 7239
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16120 5704 16172 5710
rect 16500 5658 16528 7414
rect 16592 5914 16620 7822
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16684 5794 16712 7414
rect 16776 6390 16804 8842
rect 16868 7410 16896 9930
rect 16960 9926 16988 10678
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 10062 17172 10542
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9654 17080 9862
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17038 9072 17094 9081
rect 17038 9007 17094 9016
rect 17052 8820 17080 9007
rect 17144 8974 17172 9998
rect 17236 9722 17264 9998
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17132 8832 17184 8838
rect 17052 8792 17132 8820
rect 16948 8560 17000 8566
rect 17052 8548 17080 8792
rect 17132 8774 17184 8780
rect 17000 8520 17080 8548
rect 16948 8502 17000 8508
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16960 7002 16988 8230
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7449 17080 7822
rect 17144 7546 17172 7958
rect 17236 7886 17264 9046
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17236 7546 17264 7822
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17038 7440 17094 7449
rect 17038 7375 17094 7384
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16946 6896 17002 6905
rect 16946 6831 17002 6840
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16172 5652 16528 5658
rect 16120 5646 16528 5652
rect 16132 5630 16528 5646
rect 16500 5574 16528 5630
rect 16592 5766 16712 5794
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16316 2774 16344 5510
rect 16592 5030 16620 5766
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 5370 16712 5646
rect 16776 5624 16804 6326
rect 16960 5914 16988 6831
rect 17224 6724 17276 6730
rect 17328 6712 17356 12174
rect 17512 12102 17540 13194
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 12918 17724 13126
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17604 12442 17632 12786
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17788 12170 17816 13790
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17512 11150 17540 12038
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 8634 17448 10406
rect 17512 8906 17540 11086
rect 17604 11070 17816 11098
rect 17604 10674 17632 11070
rect 17788 11014 17816 11070
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17696 9994 17724 10950
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17696 9625 17724 9930
rect 17788 9654 17816 10066
rect 17776 9648 17828 9654
rect 17682 9616 17738 9625
rect 17776 9590 17828 9596
rect 17682 9551 17738 9560
rect 17500 8900 17552 8906
rect 17776 8900 17828 8906
rect 17552 8860 17724 8888
rect 17500 8842 17552 8848
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17276 6684 17356 6712
rect 17224 6666 17276 6672
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17144 5914 17172 6190
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 16856 5636 16908 5642
rect 16776 5596 16856 5624
rect 16856 5578 16908 5584
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16500 4282 16528 4966
rect 16592 4826 16620 4966
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16868 4622 16896 5306
rect 17236 5234 17264 6190
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 3670 16528 4218
rect 17052 3738 17080 4558
rect 17144 4214 17172 4558
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 17328 3534 17356 5850
rect 17420 5098 17448 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17512 6254 17540 7482
rect 17604 6458 17632 8570
rect 17696 8566 17724 8860
rect 17776 8842 17828 8848
rect 17788 8809 17816 8842
rect 17774 8800 17830 8809
rect 17774 8735 17830 8744
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17696 7274 17724 7346
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17512 5166 17540 5578
rect 17604 5302 17632 6394
rect 17696 5370 17724 7210
rect 17880 5914 17908 13670
rect 17972 13326 18000 13670
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17960 12844 18012 12850
rect 18064 12832 18092 13806
rect 18156 13410 18184 18566
rect 18248 18465 18276 19306
rect 18524 19258 18552 19790
rect 18800 19700 18828 19994
rect 18616 19672 18828 19700
rect 18616 19514 18644 19672
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18602 19408 18658 19417
rect 18708 19394 18736 19450
rect 18658 19366 18736 19394
rect 18602 19343 18658 19352
rect 18524 19242 18828 19258
rect 18524 19236 18840 19242
rect 18524 19230 18788 19236
rect 18788 19178 18840 19184
rect 18512 19168 18564 19174
rect 18564 19128 18736 19156
rect 18512 19110 18564 19116
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18234 18456 18290 18465
rect 18234 18391 18290 18400
rect 18248 18222 18276 18391
rect 18708 18358 18736 19128
rect 18892 18698 18920 21286
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18984 20262 19012 20878
rect 19076 20806 19104 22902
rect 19536 22794 19564 24550
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19720 23338 19748 23734
rect 19812 23526 19840 25638
rect 19800 23520 19852 23526
rect 19984 23520 20036 23526
rect 19800 23462 19852 23468
rect 19982 23488 19984 23497
rect 20036 23488 20038 23497
rect 19982 23423 20038 23432
rect 19720 23310 19840 23338
rect 19614 23216 19670 23225
rect 19614 23151 19670 23160
rect 19352 22766 19564 22794
rect 19628 22778 19656 23151
rect 19812 23050 19840 23310
rect 19812 23044 19868 23050
rect 19812 22992 19816 23044
rect 19812 22986 19868 22992
rect 19616 22772 19668 22778
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19168 22166 19196 22578
rect 19352 22234 19380 22766
rect 19616 22714 19668 22720
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19156 22160 19208 22166
rect 19444 22114 19472 22442
rect 19156 22102 19208 22108
rect 19352 22086 19472 22114
rect 19352 22030 19380 22086
rect 19536 22080 19564 22578
rect 19628 22234 19656 22714
rect 19706 22264 19762 22273
rect 19616 22228 19668 22234
rect 19706 22199 19762 22208
rect 19616 22170 19668 22176
rect 19536 22052 19656 22080
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19352 21570 19380 21966
rect 19444 21690 19472 21966
rect 19628 21962 19656 22052
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19536 21690 19564 21898
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19352 21542 19472 21570
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19168 21146 19196 21422
rect 19444 21350 19472 21542
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19352 21146 19380 21286
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 19168 20618 19196 21082
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 19076 20590 19196 20618
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18248 16590 18276 18022
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18984 17354 19012 19926
rect 19076 19786 19104 20590
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19168 19922 19196 20266
rect 19260 20058 19288 21014
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20602 19380 20878
rect 19536 20874 19564 21626
rect 19524 20868 19576 20874
rect 19524 20810 19576 20816
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 19248 19712 19300 19718
rect 19076 19660 19248 19666
rect 19076 19654 19300 19660
rect 19076 19638 19288 19654
rect 19076 18630 19104 19638
rect 19352 19530 19380 19790
rect 19168 19502 19380 19530
rect 19524 19508 19576 19514
rect 19168 18970 19196 19502
rect 19524 19450 19576 19456
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19260 18970 19288 19382
rect 19340 19304 19392 19310
rect 19430 19272 19486 19281
rect 19392 19252 19430 19258
rect 19340 19246 19430 19252
rect 19352 19230 19430 19246
rect 19430 19207 19486 19216
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18465 19104 18566
rect 19062 18456 19118 18465
rect 19062 18391 19118 18400
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18616 17326 19012 17354
rect 18616 17202 18644 17326
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18340 16182 18368 16662
rect 18708 16590 18736 16934
rect 18800 16794 18828 17138
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18432 16114 18460 16390
rect 18510 16144 18566 16153
rect 18420 16108 18472 16114
rect 18510 16079 18512 16088
rect 18420 16050 18472 16056
rect 18564 16079 18566 16088
rect 18512 16050 18564 16056
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18248 13938 18276 15506
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18340 15162 18368 15370
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 15178 18644 15302
rect 18328 15156 18380 15162
rect 18616 15150 18828 15178
rect 18328 15098 18380 15104
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 14074 18368 14214
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18156 13382 18368 13410
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18012 12804 18092 12832
rect 17960 12786 18012 12792
rect 18064 12434 18092 12804
rect 17972 12406 18092 12434
rect 17972 11218 18000 12406
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17972 9722 18000 10746
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17972 9110 18000 9658
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18064 8634 18092 12174
rect 18156 9178 18184 13262
rect 18340 12866 18368 13382
rect 18248 12838 18368 12866
rect 18248 12442 18276 12838
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11898 18644 12174
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18800 11642 18828 15150
rect 18892 12442 18920 16662
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18984 13734 19012 16594
rect 19076 15502 19104 18158
rect 19168 16658 19196 18634
rect 19260 18290 19288 18906
rect 19444 18834 19472 19207
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19536 18630 19564 19450
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19628 18970 19656 19382
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19628 18630 19656 18906
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19338 17912 19394 17921
rect 19394 17876 19401 17882
rect 19338 17847 19349 17856
rect 19349 17818 19401 17824
rect 19536 17678 19564 18022
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19628 17320 19656 17546
rect 19536 17292 19656 17320
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19444 16590 19472 16934
rect 19536 16658 19564 17292
rect 19720 17218 19748 22199
rect 19812 21486 19840 22986
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19996 22234 20024 22374
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 20088 22094 20116 26726
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20272 25430 20300 25638
rect 20260 25424 20312 25430
rect 20260 25366 20312 25372
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20180 22273 20208 23190
rect 20548 23050 20576 27338
rect 20640 23322 20668 27542
rect 21192 27402 21220 27814
rect 21468 27674 21496 28494
rect 25884 28490 25912 30767
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21652 28218 21680 28358
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21640 28008 21692 28014
rect 21640 27950 21692 27956
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20824 25906 20852 27270
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20824 24886 20852 25842
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20824 24206 20852 24822
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 21100 23526 21128 24278
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20166 22264 20222 22273
rect 20166 22199 20222 22208
rect 20456 22166 20484 22374
rect 20444 22160 20496 22166
rect 20444 22102 20496 22108
rect 20088 22066 20208 22094
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19904 21554 19932 21966
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 18698 19840 21422
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19904 19922 19932 21286
rect 19996 21010 20024 21830
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19984 20800 20036 20806
rect 19982 20768 19984 20777
rect 20076 20800 20128 20806
rect 20036 20768 20038 20777
rect 20076 20742 20128 20748
rect 19982 20703 20038 20712
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19996 20058 20024 20402
rect 20088 20262 20116 20742
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19996 19689 20024 19722
rect 19982 19680 20038 19689
rect 19982 19615 20038 19624
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19996 19281 20024 19450
rect 19982 19272 20038 19281
rect 19892 19236 19944 19242
rect 19982 19207 20038 19216
rect 19892 19178 19944 19184
rect 19904 18834 19932 19178
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19800 18692 19852 18698
rect 20088 18680 20116 20198
rect 20180 18970 20208 22066
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20272 21690 20300 22034
rect 20548 21894 20576 22986
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22710 20760 22918
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20272 19310 20300 21626
rect 20444 21072 20496 21078
rect 20444 21014 20496 21020
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20168 18692 20220 18698
rect 20088 18652 20168 18680
rect 19800 18634 19852 18640
rect 20168 18634 20220 18640
rect 19628 17190 19748 17218
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19432 16448 19484 16454
rect 19430 16416 19432 16425
rect 19524 16448 19576 16454
rect 19484 16416 19486 16425
rect 19524 16390 19576 16396
rect 19430 16351 19486 16360
rect 19536 16046 19564 16390
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19168 14822 19196 15438
rect 19338 15056 19394 15065
rect 19338 14991 19394 15000
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19352 14414 19380 14991
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 18984 13326 19012 13670
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 12850 19196 13194
rect 19260 12889 19288 13670
rect 19246 12880 19302 12889
rect 19156 12844 19208 12850
rect 19246 12815 19302 12824
rect 19156 12786 19208 12792
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18800 11614 18920 11642
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18340 10810 18368 11086
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18248 10266 18276 10610
rect 18328 10600 18380 10606
rect 18326 10568 18328 10577
rect 18380 10568 18382 10577
rect 18326 10503 18382 10512
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17972 8362 18000 8502
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 17972 5914 18000 6831
rect 18064 6730 18092 7482
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 6866 18184 7210
rect 18248 7002 18276 8230
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7546 18736 7754
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18616 7188 18644 7414
rect 18616 7160 18736 7188
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18248 6186 18276 6938
rect 18708 6730 18736 7160
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 6322 18736 6666
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17868 5704 17920 5710
rect 17866 5672 17868 5681
rect 17920 5672 17922 5681
rect 17866 5607 17922 5616
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17408 5092 17460 5098
rect 17408 5034 17460 5040
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4826 17816 4966
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17512 4146 17540 4762
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17512 3534 17540 4082
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16316 2746 16436 2774
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 16408 1834 16436 2746
rect 16488 2372 16540 2378
rect 16488 2314 16540 2320
rect 16500 2106 16528 2314
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 16396 1828 16448 1834
rect 16396 1770 16448 1776
rect 16408 1562 16436 1770
rect 16396 1556 16448 1562
rect 16396 1498 16448 1504
rect 16684 1358 16712 3402
rect 17420 3194 17448 3470
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17512 2446 17540 3470
rect 18064 2922 18092 5850
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18432 5352 18460 5510
rect 18512 5364 18564 5370
rect 18432 5324 18512 5352
rect 18512 5306 18564 5312
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18708 4826 18736 6258
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4146 18644 4558
rect 18708 4214 18736 4762
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18064 2650 18092 2858
rect 18800 2774 18828 11494
rect 18892 5098 18920 11614
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18984 9178 19012 9522
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19076 8566 19104 10678
rect 19168 8820 19196 12174
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19260 11898 19288 12106
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11014 19288 11698
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19352 9994 19380 14350
rect 19536 13870 19564 14418
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13326 19564 13806
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19444 12986 19472 13194
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19628 12306 19656 17190
rect 19812 16522 19840 18634
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 17746 19932 18566
rect 20074 18320 20130 18329
rect 20074 18255 20130 18264
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19904 16590 19932 16934
rect 19996 16794 20024 17614
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19720 16250 19748 16458
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19720 14074 19748 14554
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19996 14006 20024 14758
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 20088 13818 20116 18255
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 17202 20300 17478
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20272 15094 20300 16458
rect 20364 16250 20392 20946
rect 20456 19446 20484 21014
rect 20548 20448 20576 21830
rect 20640 21622 20668 21830
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20720 20460 20772 20466
rect 20548 20420 20720 20448
rect 20720 20402 20772 20408
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20640 19786 20668 20198
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20732 19689 20760 20402
rect 20718 19680 20774 19689
rect 20718 19615 20774 19624
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20456 18902 20484 19382
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20548 18766 20576 19314
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 18834 20668 19178
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20536 18760 20588 18766
rect 20640 18737 20668 18770
rect 20536 18702 20588 18708
rect 20626 18728 20682 18737
rect 20626 18663 20682 18672
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20548 16454 20576 18090
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20536 16448 20588 16454
rect 20534 16416 20536 16425
rect 20588 16416 20590 16425
rect 20534 16351 20590 16360
rect 20640 16250 20668 17546
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20364 15366 20392 16050
rect 20456 15366 20484 16050
rect 20732 15910 20760 19615
rect 20824 18834 20852 22170
rect 21100 22098 21128 23462
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 21192 21146 21220 27338
rect 21560 27130 21588 27474
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21376 25294 21404 26318
rect 21456 26308 21508 26314
rect 21456 26250 21508 26256
rect 21468 26042 21496 26250
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21652 25770 21680 27950
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22204 27674 22232 27814
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 21640 25764 21692 25770
rect 21640 25706 21692 25712
rect 21652 25498 21680 25706
rect 21640 25492 21692 25498
rect 21640 25434 21692 25440
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21284 24954 21312 25162
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21376 23730 21404 25230
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21284 23322 21312 23666
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21284 22094 21312 22986
rect 21284 22066 21404 22094
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 20904 20868 20956 20874
rect 20904 20810 20956 20816
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20180 14414 20208 14554
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 13938 20208 14214
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 19720 13790 20024 13818
rect 20088 13790 20208 13818
rect 19720 13530 19748 13790
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19812 13530 19840 13670
rect 19996 13530 20024 13790
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19720 12442 19748 13194
rect 19996 12986 20024 13330
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 12986 20116 13194
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19984 12368 20036 12374
rect 19982 12336 19984 12345
rect 20036 12336 20038 12345
rect 19616 12300 19668 12306
rect 19982 12271 20038 12280
rect 19616 12242 19668 12248
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19904 11898 19932 12174
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19996 11694 20024 12174
rect 19984 11688 20036 11694
rect 19904 11648 19984 11676
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19628 9994 19656 10678
rect 19904 9994 19932 11648
rect 19984 11630 20036 11636
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19996 10713 20024 10746
rect 19982 10704 20038 10713
rect 19982 10639 20038 10648
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 8974 19288 9862
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19536 9178 19564 9522
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19628 8906 19656 9930
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19340 8832 19392 8838
rect 19168 8792 19288 8820
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19168 7206 19196 7822
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18984 2774 19012 7142
rect 19168 5914 19196 7142
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 3738 19104 4966
rect 19168 4729 19196 5034
rect 19154 4720 19210 4729
rect 19154 4655 19210 4664
rect 19260 4434 19288 8792
rect 19340 8774 19392 8780
rect 19352 7818 19380 8774
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19812 7546 19840 8434
rect 19904 7750 19932 9930
rect 19996 8634 20024 10639
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 7886 20024 8230
rect 20088 8090 20116 12718
rect 20180 12170 20208 13790
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 10810 20208 11698
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 20272 6458 20300 14894
rect 20364 14346 20392 15302
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20364 13870 20392 14282
rect 20456 14074 20484 15302
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20456 12918 20484 13806
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20548 12714 20576 15574
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 14890 20668 15438
rect 20824 14958 20852 18770
rect 20916 18465 20944 20810
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 21008 19786 21036 19994
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 21008 18834 21036 19178
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20902 18456 20958 18465
rect 20902 18391 20958 18400
rect 20916 18358 20944 18391
rect 21008 18358 21036 18566
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20916 15178 20944 18294
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17066 21036 17614
rect 21100 17338 21128 20810
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 21100 16794 21128 17274
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21100 16250 21128 16526
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21008 15473 21036 16050
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15502 21128 15846
rect 21088 15496 21140 15502
rect 20994 15464 21050 15473
rect 21088 15438 21140 15444
rect 20994 15399 20996 15408
rect 21048 15399 21050 15408
rect 20996 15370 21048 15376
rect 20916 15150 21128 15178
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 14074 20668 14214
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20732 13530 20760 14758
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20350 11792 20406 11801
rect 20350 11727 20352 11736
rect 20404 11727 20406 11736
rect 20352 11698 20404 11704
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 11286 20392 11494
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20456 10554 20484 12038
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20548 10742 20576 10950
rect 20536 10736 20588 10742
rect 20536 10678 20588 10684
rect 20456 10526 20576 10554
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20364 9722 20392 10202
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9761 20484 9862
rect 20442 9752 20498 9761
rect 20352 9716 20404 9722
rect 20442 9687 20498 9696
rect 20352 9658 20404 9664
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5710 19380 6054
rect 19444 5914 19472 6326
rect 20456 6118 20484 8298
rect 20548 7993 20576 10526
rect 20640 10266 20668 13262
rect 20718 12880 20774 12889
rect 20718 12815 20774 12824
rect 20732 12646 20760 12815
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20824 12434 20852 14350
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 14074 20944 14282
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20732 12406 20852 12434
rect 20732 11150 20760 12406
rect 20812 12368 20864 12374
rect 20916 12345 20944 13874
rect 21008 13530 21036 14826
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21008 12374 21036 12786
rect 20996 12368 21048 12374
rect 20812 12310 20864 12316
rect 20902 12336 20958 12345
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20732 10062 20760 11086
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9874 20760 9998
rect 20640 9846 20760 9874
rect 20640 9382 20668 9846
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20732 8974 20760 9658
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20732 8022 20760 8434
rect 20720 8016 20772 8022
rect 20534 7984 20590 7993
rect 20720 7958 20772 7964
rect 20534 7919 20590 7928
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20732 6798 20760 7822
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20364 5914 20392 6054
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20272 4826 20300 5170
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19168 4406 19288 4434
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18708 2746 18828 2774
rect 18892 2746 19012 2774
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17512 2106 17540 2382
rect 18708 2310 18736 2746
rect 18892 2650 18920 2746
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 2106 18736 2246
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 17408 1964 17460 1970
rect 17408 1906 17460 1912
rect 17040 1760 17092 1766
rect 17040 1702 17092 1708
rect 17052 1494 17080 1702
rect 17420 1562 17448 1906
rect 18892 1834 18920 2586
rect 18880 1828 18932 1834
rect 18880 1770 18932 1776
rect 18315 1660 18623 1669
rect 18315 1658 18321 1660
rect 18377 1658 18401 1660
rect 18457 1658 18481 1660
rect 18537 1658 18561 1660
rect 18617 1658 18623 1660
rect 18377 1606 18379 1658
rect 18559 1606 18561 1658
rect 18315 1604 18321 1606
rect 18377 1604 18401 1606
rect 18457 1604 18481 1606
rect 18537 1604 18561 1606
rect 18617 1604 18623 1606
rect 18315 1595 18623 1604
rect 19168 1562 19196 4406
rect 19720 4282 19748 4490
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19444 3738 19472 3946
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 20088 3534 20116 4558
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 19260 3126 19288 3402
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19260 1970 19288 3062
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19536 2106 19564 2790
rect 19720 2650 19748 2858
rect 20364 2650 20392 4966
rect 20456 4826 20484 5714
rect 20548 5370 20576 6190
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5574 20760 6054
rect 20824 5914 20852 12310
rect 20996 12310 21048 12316
rect 20902 12271 20958 12280
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20916 11694 20944 12038
rect 21100 11914 21128 15150
rect 21192 12850 21220 20742
rect 21284 15502 21312 21286
rect 21376 20058 21404 22066
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21468 21146 21496 21898
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21376 18086 21404 19994
rect 21652 19496 21680 23462
rect 22204 23118 22232 27610
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22940 26858 22968 27270
rect 24412 26994 24440 27406
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 23940 26988 23992 26994
rect 23940 26930 23992 26936
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 22928 26852 22980 26858
rect 22928 26794 22980 26800
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22388 24750 22416 25094
rect 22480 24954 22508 25162
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22376 24744 22428 24750
rect 22376 24686 22428 24692
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23118 22324 24006
rect 22388 23118 22416 24686
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22112 20262 22140 20470
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 21652 19468 21956 19496
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21376 16658 21404 17478
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 14822 21312 15438
rect 21376 15026 21404 16186
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21376 13938 21404 14962
rect 21468 14890 21496 18090
rect 21546 17912 21602 17921
rect 21546 17847 21602 17856
rect 21560 17338 21588 17847
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21362 13288 21418 13297
rect 21362 13223 21364 13232
rect 21416 13223 21418 13232
rect 21364 13194 21416 13200
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21272 12640 21324 12646
rect 21192 12600 21272 12628
rect 21192 12345 21220 12600
rect 21272 12582 21324 12588
rect 21376 12442 21404 12922
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21178 12336 21234 12345
rect 21468 12306 21496 14010
rect 21178 12271 21234 12280
rect 21456 12300 21508 12306
rect 21192 12238 21220 12271
rect 21456 12242 21508 12248
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21178 12064 21234 12073
rect 21178 11999 21234 12008
rect 21008 11886 21128 11914
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20916 6390 20944 11630
rect 21008 9432 21036 11886
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21100 11014 21128 11698
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10742 21128 10950
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21192 10554 21220 11999
rect 21454 11928 21510 11937
rect 21454 11863 21510 11872
rect 21364 11756 21416 11762
rect 21284 11716 21364 11744
rect 21284 10742 21312 11716
rect 21364 11698 21416 11704
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11150 21404 11494
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21192 10526 21404 10554
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21192 9722 21220 9930
rect 21284 9722 21312 10406
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21088 9444 21140 9450
rect 21008 9404 21088 9432
rect 21088 9386 21140 9392
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 8634 21220 9318
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21008 8430 21036 8502
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 8090 21220 8230
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20904 6248 20956 6254
rect 21008 6236 21036 7958
rect 21376 7750 21404 10526
rect 21468 9382 21496 11863
rect 21560 11558 21588 17138
rect 21652 16250 21680 19246
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21744 18902 21772 19178
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21822 18728 21878 18737
rect 21822 18663 21878 18672
rect 21836 18630 21864 18663
rect 21928 18630 21956 19468
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 21916 18216 21968 18222
rect 21914 18184 21916 18193
rect 21968 18184 21970 18193
rect 21914 18119 21970 18128
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22112 16590 22140 17138
rect 22204 16998 22232 22918
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22296 21622 22324 22646
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22296 21010 22324 21558
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22296 20058 22324 20402
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22388 18970 22416 21286
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22374 18864 22430 18873
rect 22284 18828 22336 18834
rect 22374 18799 22430 18808
rect 22284 18770 22336 18776
rect 22296 18630 22324 18770
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 18329 22324 18566
rect 22388 18358 22416 18799
rect 22376 18352 22428 18358
rect 22282 18320 22338 18329
rect 22376 18294 22428 18300
rect 22282 18255 22338 18264
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22296 17882 22324 18158
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 22388 16266 22416 18158
rect 22480 18086 22508 23462
rect 22572 21486 22600 25842
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22664 23186 22692 23666
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22756 22574 22784 24074
rect 22848 23254 22876 24074
rect 22940 23798 22968 26794
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23032 26586 23060 26726
rect 23020 26580 23072 26586
rect 23020 26522 23072 26528
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 22836 23248 22888 23254
rect 22834 23216 22836 23225
rect 22888 23216 22890 23225
rect 22834 23151 22890 23160
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22756 22234 22784 22510
rect 22848 22234 22876 23054
rect 23032 23050 23060 24006
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 23032 22094 23060 22986
rect 22756 22066 23060 22094
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22664 21350 22692 21830
rect 22756 21554 22784 22066
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 20466 22600 20878
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22572 20058 22600 20402
rect 22756 20262 22784 21490
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 21146 22876 21286
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22848 18834 22876 20946
rect 22940 20942 22968 21966
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22940 20466 22968 20878
rect 23032 20806 23060 21966
rect 23124 21418 23152 26726
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23216 23866 23244 24142
rect 23308 24138 23336 26862
rect 23952 26586 23980 26930
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 24412 25294 24440 26930
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 25870 25936 25926 25945
rect 25870 25871 25926 25880
rect 25780 25764 25832 25770
rect 25780 25706 25832 25712
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25792 25498 25820 25706
rect 25884 25702 25912 25871
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24308 25220 24360 25226
rect 24308 25162 24360 25168
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23676 24954 23704 25094
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23308 22094 23336 24074
rect 23768 23730 23796 25094
rect 24136 24750 24164 25162
rect 24320 24954 24348 25162
rect 24308 24948 24360 24954
rect 24308 24890 24360 24896
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24412 24206 24440 25230
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 24952 24676 25004 24682
rect 24952 24618 25004 24624
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23400 23118 23428 23190
rect 23492 23118 23520 23666
rect 23952 23322 23980 23666
rect 24412 23662 24440 24142
rect 24780 23866 24808 24550
rect 24964 24070 24992 24618
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 24412 23118 24440 23598
rect 24964 23118 24992 24006
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 23940 23044 23992 23050
rect 23940 22986 23992 22992
rect 23952 22778 23980 22986
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 25148 22710 25176 24686
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25792 22778 25820 22918
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23216 22066 23336 22094
rect 23216 21622 23244 22066
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23308 21434 23336 21966
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21690 23520 21830
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23216 21406 23336 21434
rect 23124 21146 23152 21354
rect 23216 21350 23244 21406
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23216 21026 23244 21286
rect 23124 20998 23244 21026
rect 23124 20874 23152 20998
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23124 20618 23152 20810
rect 23032 20590 23152 20618
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22940 19854 22968 20198
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22572 18426 22600 18702
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 16794 22508 17070
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 21640 16244 21692 16250
rect 22388 16238 22508 16266
rect 21640 16186 21692 16192
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21836 15706 21864 15846
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21652 15094 21680 15302
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21640 14952 21692 14958
rect 21744 14929 21772 15098
rect 21640 14894 21692 14900
rect 21730 14920 21786 14929
rect 21652 12918 21680 14894
rect 21730 14855 21786 14864
rect 22204 14618 22232 15370
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22020 13530 22048 13806
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22100 13456 22152 13462
rect 22204 13444 22232 14214
rect 22388 14074 22416 16118
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22152 13416 22232 13444
rect 22100 13398 22152 13404
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21652 11762 21680 12582
rect 22020 12458 22048 12786
rect 22204 12714 22232 13416
rect 22282 13288 22338 13297
rect 22388 13258 22416 13670
rect 22282 13223 22338 13232
rect 22376 13252 22428 13258
rect 22296 12850 22324 13223
rect 22376 13194 22428 13200
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22020 12434 22324 12458
rect 22020 12430 22416 12434
rect 22296 12406 22416 12430
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 21916 11892 21968 11898
rect 21836 11852 21916 11880
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21640 11620 21692 11626
rect 21836 11608 21864 11852
rect 22204 11880 22232 12038
rect 21916 11834 21968 11840
rect 22112 11852 22232 11880
rect 22008 11824 22060 11830
rect 22006 11792 22008 11801
rect 22060 11792 22062 11801
rect 21916 11756 21968 11762
rect 22006 11727 22062 11736
rect 21916 11698 21968 11704
rect 21692 11580 21864 11608
rect 21640 11562 21692 11568
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21928 11082 21956 11698
rect 22112 11626 22140 11852
rect 22192 11756 22244 11762
rect 22244 11716 22324 11744
rect 22192 11698 22244 11704
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22204 10266 22232 10406
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 21652 9382 21680 9862
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 21732 9648 21784 9654
rect 22008 9648 22060 9654
rect 21732 9590 21784 9596
rect 22006 9616 22008 9625
rect 22060 9616 22062 9625
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21744 9194 21772 9590
rect 22006 9551 22062 9560
rect 21652 9166 21772 9194
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 8378 21496 8842
rect 21652 8838 21680 9166
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21560 8566 21588 8774
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21652 8430 21680 8774
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21732 8560 21784 8566
rect 22008 8560 22060 8566
rect 21784 8520 22008 8548
rect 21732 8502 21784 8508
rect 22204 8537 22232 9862
rect 22008 8502 22060 8508
rect 22190 8528 22246 8537
rect 22190 8463 22246 8472
rect 21640 8424 21692 8430
rect 21546 8392 21602 8401
rect 21468 8350 21546 8378
rect 21640 8366 21692 8372
rect 21824 8424 21876 8430
rect 21876 8384 22232 8412
rect 21824 8366 21876 8372
rect 21546 8327 21602 8336
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21192 7546 21220 7686
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6458 21128 6598
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20956 6208 21036 6236
rect 20904 6190 20956 6196
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20824 5234 20852 5850
rect 21008 5624 21036 6208
rect 21088 5636 21140 5642
rect 21008 5596 21088 5624
rect 21008 5234 21036 5596
rect 21088 5578 21140 5584
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20824 4282 20852 4966
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21008 4282 21036 4490
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 21284 3670 21312 6734
rect 21376 6322 21404 7686
rect 21468 7002 21496 7890
rect 21560 7818 21588 8327
rect 22204 7886 22232 8384
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 22112 7274 22140 7482
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22204 7002 22232 7142
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22296 6798 22324 11716
rect 22388 11626 22416 12406
rect 22480 11898 22508 16238
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 15026 22600 15302
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22376 11620 22428 11626
rect 22376 11562 22428 11568
rect 22388 9926 22416 11562
rect 22572 11150 22600 12310
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22664 10810 22692 18702
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18329 22784 18566
rect 22742 18320 22798 18329
rect 22742 18255 22798 18264
rect 22928 18216 22980 18222
rect 22756 18164 22928 18170
rect 22756 18158 22980 18164
rect 22756 18142 22968 18158
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22480 9722 22508 10406
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22388 9110 22416 9590
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21652 6458 21680 6666
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 22388 6390 22416 7142
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21376 5642 21404 6258
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22204 5914 22232 6122
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22112 4570 22140 5102
rect 22112 4542 22232 4570
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 21652 2922 21680 4014
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 21640 2916 21692 2922
rect 21640 2858 21692 2864
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20824 2446 20852 2790
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 19616 2372 19668 2378
rect 19616 2314 19668 2320
rect 19628 2106 19656 2314
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19248 1964 19300 1970
rect 19248 1906 19300 1912
rect 19616 1964 19668 1970
rect 19616 1906 19668 1912
rect 19248 1760 19300 1766
rect 19248 1702 19300 1708
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 19156 1556 19208 1562
rect 19156 1498 19208 1504
rect 17040 1488 17092 1494
rect 17040 1430 17092 1436
rect 19260 1358 19288 1702
rect 19628 1562 19656 1906
rect 19904 1902 19932 2382
rect 21652 1970 21680 2858
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 21640 1964 21692 1970
rect 21640 1906 21692 1912
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 21468 1562 21496 1906
rect 22204 1766 22232 4542
rect 22296 4146 22324 6190
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22480 3194 22508 9114
rect 22572 8090 22600 10406
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22664 9586 22692 9930
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22664 8906 22692 9522
rect 22756 8974 22784 18142
rect 22928 18080 22980 18086
rect 22926 18048 22928 18057
rect 22980 18048 22982 18057
rect 22926 17983 22982 17992
rect 23032 17898 23060 20590
rect 23584 19802 23612 22102
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21146 23704 21286
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 24504 21010 24532 22646
rect 26344 22506 26372 23462
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 24964 22030 24992 22374
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25700 22094 25728 22374
rect 26344 22234 26372 22442
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 25700 22066 25820 22094
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21486 24900 21830
rect 25134 21584 25190 21593
rect 25792 21554 25820 22066
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 26160 21690 26188 21898
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 25134 21519 25190 21528
rect 25780 21548 25832 21554
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 21146 24900 21422
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24492 21004 24544 21010
rect 24492 20946 24544 20952
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23768 20534 23796 20742
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23756 19848 23808 19854
rect 23584 19774 23704 19802
rect 23756 19790 23808 19796
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23584 19514 23612 19654
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23110 18184 23166 18193
rect 23216 18170 23244 18226
rect 23166 18142 23244 18170
rect 23110 18119 23166 18128
rect 22940 17870 23060 17898
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22848 15366 22876 16186
rect 22940 15434 22968 17870
rect 23124 17746 23152 18119
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23216 17338 23244 17614
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23124 16674 23152 17070
rect 23216 16794 23244 17274
rect 23400 16794 23428 17546
rect 23492 17218 23520 18634
rect 23584 17814 23612 18838
rect 23676 18766 23704 19774
rect 23768 18970 23796 19790
rect 24504 19446 24532 20946
rect 25148 20806 25176 21519
rect 25780 21490 25832 21496
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20534 26280 20742
rect 26344 20602 26372 21966
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24964 19854 24992 20402
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 26344 19854 26372 20538
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25424 19514 25452 19722
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 24492 19440 24544 19446
rect 24136 19400 24492 19428
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18970 23980 19110
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 24136 18698 24164 19400
rect 24492 19382 24544 19388
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 23860 18290 23888 18566
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 23584 17338 23612 17750
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23492 17190 23612 17218
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23124 16646 23244 16674
rect 23216 15978 23244 16646
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15706 23152 15846
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 9926 22876 13806
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12918 23060 13126
rect 23020 12912 23072 12918
rect 23020 12854 23072 12860
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23032 11830 23060 12718
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22940 9722 22968 11698
rect 23032 10674 23060 11766
rect 23216 11218 23244 15914
rect 23388 15360 23440 15366
rect 23308 15320 23388 15348
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23308 11150 23336 15320
rect 23492 15337 23520 16526
rect 23584 16522 23612 17190
rect 23676 16697 23704 17614
rect 23768 16794 23796 17614
rect 23952 17338 23980 17750
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24044 17202 24072 18566
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24228 17082 24256 18634
rect 24504 18442 24532 19246
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18970 24624 19110
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25884 18970 25912 19314
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25976 18834 26004 19790
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 24504 18414 24624 18442
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24320 17882 24348 18226
rect 24596 18222 24624 18414
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24596 17542 24624 18158
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25148 17678 25176 17818
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 25504 17604 25556 17610
rect 25504 17546 25556 17552
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24136 17054 24256 17082
rect 24596 17354 24624 17478
rect 24596 17338 24716 17354
rect 24596 17332 24728 17338
rect 24596 17326 24676 17332
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23848 16720 23900 16726
rect 23662 16688 23718 16697
rect 23848 16662 23900 16668
rect 23662 16623 23718 16632
rect 23860 16522 23888 16662
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 24136 15978 24164 17054
rect 24596 16658 24624 17326
rect 24676 17274 24728 17280
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24596 16114 24624 16594
rect 24780 16250 24808 17546
rect 25516 17338 25544 17546
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25608 16794 25636 17138
rect 25700 16969 25728 18770
rect 26252 18766 26280 19110
rect 26240 18760 26292 18766
rect 25778 18728 25834 18737
rect 26240 18702 26292 18708
rect 25778 18663 25834 18672
rect 26700 18692 26752 18698
rect 25686 16960 25742 16969
rect 25686 16895 25742 16904
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24124 15972 24176 15978
rect 24124 15914 24176 15920
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23388 15302 23440 15308
rect 23478 15328 23534 15337
rect 23478 15263 23534 15272
rect 23768 15144 23796 15574
rect 24136 15434 24164 15914
rect 24320 15706 24348 16050
rect 24780 15706 24808 16050
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24768 15496 24820 15502
rect 24766 15464 24768 15473
rect 24820 15464 24822 15473
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 24124 15428 24176 15434
rect 24766 15399 24822 15408
rect 24124 15370 24176 15376
rect 24044 15314 24072 15370
rect 24044 15286 24164 15314
rect 23676 15116 23796 15144
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 14550 23520 14758
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12714 23428 13126
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23400 11762 23428 12650
rect 23492 12238 23520 12718
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23584 11370 23612 12650
rect 23676 11558 23704 15116
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14618 23796 14962
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23768 13530 23796 13874
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23860 13308 23888 14350
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 23768 13280 23888 13308
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23492 11342 23612 11370
rect 23492 11234 23520 11342
rect 23400 11206 23520 11234
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23112 10736 23164 10742
rect 23308 10713 23336 11086
rect 23400 10810 23428 11206
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23112 10678 23164 10684
rect 23294 10704 23350 10713
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23020 10532 23072 10538
rect 23020 10474 23072 10480
rect 23032 10169 23060 10474
rect 23018 10160 23074 10169
rect 23018 10095 23074 10104
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22848 8838 22876 9386
rect 22836 8832 22888 8838
rect 22650 8800 22706 8809
rect 22836 8774 22888 8780
rect 22650 8735 22706 8744
rect 22664 8634 22692 8735
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22572 7002 22600 7346
rect 22650 7304 22706 7313
rect 22650 7239 22706 7248
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22664 5234 22692 7239
rect 22756 6390 22784 7822
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22848 5386 22876 8774
rect 22940 5658 22968 9658
rect 23018 9616 23074 9625
rect 23018 9551 23074 9560
rect 23032 9178 23060 9551
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 23124 6934 23152 10678
rect 23492 10674 23520 11018
rect 23294 10639 23350 10648
rect 23480 10668 23532 10674
rect 23308 10588 23336 10639
rect 23480 10610 23532 10616
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23388 10600 23440 10606
rect 23308 10560 23388 10588
rect 23388 10542 23440 10548
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23020 6656 23072 6662
rect 23124 6610 23152 6870
rect 23072 6604 23152 6610
rect 23020 6598 23152 6604
rect 23032 6582 23152 6598
rect 22940 5630 23060 5658
rect 23032 5574 23060 5630
rect 23020 5568 23072 5574
rect 22926 5536 22982 5545
rect 23020 5510 23072 5516
rect 22926 5471 22982 5480
rect 22756 5358 22876 5386
rect 22756 5302 22784 5358
rect 22744 5296 22796 5302
rect 22744 5238 22796 5244
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4826 22692 4966
rect 22756 4842 22784 5102
rect 22848 4978 22876 5358
rect 22940 5098 22968 5471
rect 23032 5302 23060 5510
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22928 5092 22980 5098
rect 22928 5034 22980 5040
rect 22848 4950 23152 4978
rect 22652 4820 22704 4826
rect 22756 4814 22876 4842
rect 22652 4762 22704 4768
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22572 4282 22600 4626
rect 22848 4554 22876 4814
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 22296 2378 22324 3062
rect 22664 2650 22692 3470
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3194 22876 3334
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 23032 2582 23060 4762
rect 23124 4554 23152 4950
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23216 3602 23244 10202
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23308 8634 23336 8910
rect 23584 8634 23612 10610
rect 23676 10266 23704 11222
rect 23768 10674 23796 13280
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23860 12442 23888 12786
rect 23952 12782 23980 13398
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23860 10810 23888 11154
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23952 10554 23980 11494
rect 23860 10526 23980 10554
rect 24032 10532 24084 10538
rect 23860 10266 23888 10526
rect 24032 10474 24084 10480
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23756 10192 23808 10198
rect 23756 10134 23808 10140
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23676 8809 23704 9998
rect 23768 9178 23796 10134
rect 23952 10062 23980 10406
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 24044 9926 24072 10474
rect 24032 9920 24084 9926
rect 23952 9880 24032 9908
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23662 8800 23718 8809
rect 23662 8735 23718 8744
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23480 8560 23532 8566
rect 23400 8520 23480 8548
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 23308 7546 23336 7754
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23308 6322 23336 6598
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23400 6118 23428 8520
rect 23480 8502 23532 8508
rect 23664 8560 23716 8566
rect 23768 8548 23796 8842
rect 23952 8838 23980 9880
rect 24032 9862 24084 9868
rect 24136 9654 24164 15286
rect 24780 14414 24808 15399
rect 24872 15094 24900 16458
rect 25148 15638 25176 16662
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25700 15706 25728 16118
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25136 15632 25188 15638
rect 25136 15574 25188 15580
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24964 15162 24992 15438
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24872 14906 24900 15030
rect 25596 14952 25648 14958
rect 24872 14878 24992 14906
rect 25596 14894 25648 14900
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24412 12889 24440 13126
rect 24398 12880 24454 12889
rect 24398 12815 24454 12824
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 11234 24440 12582
rect 24412 11206 24716 11234
rect 24872 11218 24900 14758
rect 24964 14482 24992 14878
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 25608 14278 25636 14894
rect 25700 14890 25728 15642
rect 25688 14884 25740 14890
rect 25688 14826 25740 14832
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24964 13326 24992 14010
rect 25608 13870 25636 14214
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 25136 13184 25188 13190
rect 25136 13126 25188 13132
rect 24964 12850 24992 13126
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 25056 12434 25084 12922
rect 25148 12918 25176 13126
rect 25608 12986 25636 13806
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25136 12912 25188 12918
rect 25136 12854 25188 12860
rect 25228 12640 25280 12646
rect 24964 12406 25084 12434
rect 25148 12600 25228 12628
rect 24964 11830 24992 12406
rect 25148 12322 25176 12600
rect 25228 12582 25280 12588
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25056 12294 25176 12322
rect 25056 12238 25084 12294
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24228 10266 24256 11086
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 24044 8634 24072 8910
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23716 8520 23796 8548
rect 23848 8560 23900 8566
rect 23664 8502 23716 8508
rect 23848 8502 23900 8508
rect 23860 8401 23888 8502
rect 23846 8392 23902 8401
rect 23846 8327 23902 8336
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23492 6458 23520 8026
rect 23584 7478 23612 8026
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23400 5370 23428 6054
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 4826 23428 5102
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23492 4622 23520 5170
rect 23480 4616 23532 4622
rect 23676 4570 23704 8230
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7478 23888 7686
rect 24136 7546 24164 8230
rect 24320 7818 24348 10610
rect 24412 8090 24440 11018
rect 24688 10742 24716 11206
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24964 10742 24992 11766
rect 25424 11626 25452 12038
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25608 11150 25636 11494
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24952 10736 25004 10742
rect 24952 10678 25004 10684
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24504 10130 24532 10474
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 24320 7274 24348 7754
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24308 7268 24360 7274
rect 24308 7210 24360 7216
rect 24412 7002 24440 7414
rect 24504 7410 24532 8366
rect 24596 8362 24624 9862
rect 24584 8356 24636 8362
rect 24584 8298 24636 8304
rect 24596 7954 24624 8298
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 23756 6724 23808 6730
rect 23756 6666 23808 6672
rect 23768 6390 23796 6666
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24412 5914 24440 6054
rect 24504 5914 24532 6054
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23768 5234 23796 5510
rect 24688 5370 24716 10678
rect 25700 10538 25728 14214
rect 25792 12345 25820 18663
rect 26700 18634 26752 18640
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18426 26004 18566
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 26712 18290 26740 18634
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 26700 18284 26752 18290
rect 26700 18226 26752 18232
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26528 17814 26556 18022
rect 26516 17808 26568 17814
rect 26516 17750 26568 17756
rect 26712 17610 26740 18226
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26896 17678 26924 18022
rect 26988 17678 27016 18158
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26252 17490 26280 17546
rect 26160 17462 26280 17490
rect 26160 16250 26188 17462
rect 26252 17270 26280 17462
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26436 16250 26464 16458
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26988 16114 27016 17614
rect 27436 17604 27488 17610
rect 27436 17546 27488 17552
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 27080 16590 27108 17478
rect 27448 17338 27476 17546
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 27172 16454 27200 17138
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27540 16250 27568 16390
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25884 15638 25912 15846
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27448 15162 27476 15370
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 26976 14884 27028 14890
rect 26976 14826 27028 14832
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26344 14414 26372 14758
rect 26988 14414 27016 14826
rect 27264 14618 27292 14962
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 27528 14544 27580 14550
rect 27528 14486 27580 14492
rect 26332 14408 26384 14414
rect 26332 14350 26384 14356
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26988 13938 27016 14350
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25976 12434 26004 13194
rect 26160 12986 26188 13670
rect 26988 13530 27016 13874
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26252 12986 26280 13194
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26988 12850 27016 13466
rect 27356 13394 27384 14282
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27448 12442 27476 12786
rect 27436 12436 27488 12442
rect 25976 12406 26280 12434
rect 25778 12336 25834 12345
rect 25778 12271 25834 12280
rect 26252 11694 26280 12406
rect 27436 12378 27488 12384
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 26712 11694 26740 12174
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26252 11150 26280 11630
rect 27356 11354 27384 12174
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27448 11354 27476 11698
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 25688 10532 25740 10538
rect 25688 10474 25740 10480
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24780 9722 24808 9930
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24964 9382 24992 10134
rect 25884 10062 25912 10406
rect 26252 10266 26280 11086
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26896 10742 26924 11018
rect 27448 10810 27476 11086
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 26884 10736 26936 10742
rect 26884 10678 26936 10684
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 26896 9654 26924 10678
rect 27540 10146 27568 14486
rect 28460 14006 28488 15438
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28276 13530 28304 13874
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 27620 13456 27672 13462
rect 27618 13424 27620 13433
rect 27672 13424 27674 13433
rect 27618 13359 27674 13368
rect 27632 12986 27660 13359
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 27618 10160 27674 10169
rect 27540 10118 27618 10146
rect 27618 10095 27674 10104
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27252 9920 27304 9926
rect 27252 9862 27304 9868
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 27264 9450 27292 9862
rect 27540 9722 27568 9930
rect 27528 9716 27580 9722
rect 27528 9658 27580 9664
rect 27252 9444 27304 9450
rect 27252 9386 27304 9392
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 8974 24992 9318
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 27632 9178 27660 10095
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 24872 8634 24900 8842
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25884 8634 25912 8774
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 24872 8514 24900 8570
rect 26344 8566 26372 8842
rect 26620 8634 26648 8910
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 24780 8486 24900 8514
rect 26332 8560 26384 8566
rect 26332 8502 26384 8508
rect 24780 7750 24808 8486
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24780 6458 24808 7686
rect 25792 7546 25820 7890
rect 25884 7857 25912 7890
rect 25870 7848 25926 7857
rect 25870 7783 25926 7792
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 24872 6798 24900 7482
rect 26344 7478 26372 8502
rect 26606 7984 26662 7993
rect 26606 7919 26662 7928
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 26620 7274 26648 7919
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26804 7546 26832 7822
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 26988 7546 27016 7686
rect 28368 7546 28396 7686
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 26608 7268 26660 7274
rect 26660 7228 26740 7256
rect 26608 7210 26660 7216
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 26712 7002 26740 7228
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 25780 6792 25832 6798
rect 25780 6734 25832 6740
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23480 4558 23532 4564
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23308 4282 23336 4490
rect 23492 4282 23520 4558
rect 23584 4542 23704 4570
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23584 3942 23612 4542
rect 24872 4486 24900 6258
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24964 5642 24992 6122
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5914 25084 6054
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25792 5710 25820 6734
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 26160 6458 26188 6666
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 24952 5636 25004 5642
rect 24952 5578 25004 5584
rect 24964 5370 24992 5578
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23584 3738 23612 3878
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23676 3534 23704 4422
rect 23768 4214 23796 4422
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23860 3738 23888 4082
rect 25056 4078 25084 5510
rect 25792 5234 25820 5646
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 5302 26096 5510
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 25056 2990 25084 4014
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25884 3097 25912 3946
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 25870 3088 25926 3097
rect 25870 3023 25926 3032
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 23020 2576 23072 2582
rect 23020 2518 23072 2524
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 19616 1556 19668 1562
rect 19616 1498 19668 1504
rect 21456 1556 21508 1562
rect 21456 1498 21508 1504
rect 22204 1494 22232 1702
rect 22192 1488 22244 1494
rect 22192 1430 22244 1436
rect 22296 1426 22324 2314
rect 23032 2106 23060 2518
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 25261 1660 25569 1669
rect 25261 1658 25267 1660
rect 25323 1658 25347 1660
rect 25403 1658 25427 1660
rect 25483 1658 25507 1660
rect 25563 1658 25569 1660
rect 25323 1606 25325 1658
rect 25505 1606 25507 1658
rect 25261 1604 25267 1606
rect 25323 1604 25347 1606
rect 25403 1604 25427 1606
rect 25483 1604 25507 1606
rect 25563 1604 25569 1606
rect 25261 1595 25569 1604
rect 22284 1420 22336 1426
rect 22284 1362 22336 1368
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 16672 1352 16724 1358
rect 16672 1294 16724 1300
rect 19248 1352 19300 1358
rect 19248 1294 19300 1300
rect 7896 1116 8204 1125
rect 7896 1114 7902 1116
rect 7958 1114 7982 1116
rect 8038 1114 8062 1116
rect 8118 1114 8142 1116
rect 8198 1114 8204 1116
rect 7958 1062 7960 1114
rect 8140 1062 8142 1114
rect 7896 1060 7902 1062
rect 7958 1060 7982 1062
rect 8038 1060 8062 1062
rect 8118 1060 8142 1062
rect 8198 1060 8204 1062
rect 7896 1051 8204 1060
rect 14842 1116 15150 1125
rect 14842 1114 14848 1116
rect 14904 1114 14928 1116
rect 14984 1114 15008 1116
rect 15064 1114 15088 1116
rect 15144 1114 15150 1116
rect 14904 1062 14906 1114
rect 15086 1062 15088 1114
rect 14842 1060 14848 1062
rect 14904 1060 14928 1062
rect 14984 1060 15008 1062
rect 15064 1060 15088 1062
rect 15144 1060 15150 1062
rect 14842 1051 15150 1060
rect 21788 1116 22096 1125
rect 21788 1114 21794 1116
rect 21850 1114 21874 1116
rect 21930 1114 21954 1116
rect 22010 1114 22034 1116
rect 22090 1114 22096 1116
rect 21850 1062 21852 1114
rect 22032 1062 22034 1114
rect 21788 1060 21794 1062
rect 21850 1060 21874 1062
rect 21930 1060 21954 1062
rect 22010 1060 22034 1062
rect 22090 1060 22096 1062
rect 21788 1051 22096 1060
rect 28734 1116 29042 1125
rect 28734 1114 28740 1116
rect 28796 1114 28820 1116
rect 28876 1114 28900 1116
rect 28956 1114 28980 1116
rect 29036 1114 29042 1116
rect 28796 1062 28798 1114
rect 28978 1062 28980 1114
rect 28734 1060 28740 1062
rect 28796 1060 28820 1062
rect 28876 1060 28900 1062
rect 28956 1060 28980 1062
rect 29036 1060 29042 1062
rect 28734 1051 29042 1060
<< via2 >>
rect 7902 32666 7958 32668
rect 7982 32666 8038 32668
rect 8062 32666 8118 32668
rect 8142 32666 8198 32668
rect 7902 32614 7948 32666
rect 7948 32614 7958 32666
rect 7982 32614 8012 32666
rect 8012 32614 8024 32666
rect 8024 32614 8038 32666
rect 8062 32614 8076 32666
rect 8076 32614 8088 32666
rect 8088 32614 8118 32666
rect 8142 32614 8152 32666
rect 8152 32614 8198 32666
rect 7902 32612 7958 32614
rect 7982 32612 8038 32614
rect 8062 32612 8118 32614
rect 8142 32612 8198 32614
rect 14848 32666 14904 32668
rect 14928 32666 14984 32668
rect 15008 32666 15064 32668
rect 15088 32666 15144 32668
rect 14848 32614 14894 32666
rect 14894 32614 14904 32666
rect 14928 32614 14958 32666
rect 14958 32614 14970 32666
rect 14970 32614 14984 32666
rect 15008 32614 15022 32666
rect 15022 32614 15034 32666
rect 15034 32614 15064 32666
rect 15088 32614 15098 32666
rect 15098 32614 15144 32666
rect 14848 32612 14904 32614
rect 14928 32612 14984 32614
rect 15008 32612 15064 32614
rect 15088 32612 15144 32614
rect 21794 32666 21850 32668
rect 21874 32666 21930 32668
rect 21954 32666 22010 32668
rect 22034 32666 22090 32668
rect 21794 32614 21840 32666
rect 21840 32614 21850 32666
rect 21874 32614 21904 32666
rect 21904 32614 21916 32666
rect 21916 32614 21930 32666
rect 21954 32614 21968 32666
rect 21968 32614 21980 32666
rect 21980 32614 22010 32666
rect 22034 32614 22044 32666
rect 22044 32614 22090 32666
rect 21794 32612 21850 32614
rect 21874 32612 21930 32614
rect 21954 32612 22010 32614
rect 22034 32612 22090 32614
rect 28740 32666 28796 32668
rect 28820 32666 28876 32668
rect 28900 32666 28956 32668
rect 28980 32666 29036 32668
rect 28740 32614 28786 32666
rect 28786 32614 28796 32666
rect 28820 32614 28850 32666
rect 28850 32614 28862 32666
rect 28862 32614 28876 32666
rect 28900 32614 28914 32666
rect 28914 32614 28926 32666
rect 28926 32614 28956 32666
rect 28980 32614 28990 32666
rect 28990 32614 29036 32666
rect 28740 32612 28796 32614
rect 28820 32612 28876 32614
rect 28900 32612 28956 32614
rect 28980 32612 29036 32614
rect 4429 32122 4485 32124
rect 4509 32122 4565 32124
rect 4589 32122 4645 32124
rect 4669 32122 4725 32124
rect 4429 32070 4475 32122
rect 4475 32070 4485 32122
rect 4509 32070 4539 32122
rect 4539 32070 4551 32122
rect 4551 32070 4565 32122
rect 4589 32070 4603 32122
rect 4603 32070 4615 32122
rect 4615 32070 4645 32122
rect 4669 32070 4679 32122
rect 4679 32070 4725 32122
rect 4429 32068 4485 32070
rect 4509 32068 4565 32070
rect 4589 32068 4645 32070
rect 4669 32068 4725 32070
rect 11375 32122 11431 32124
rect 11455 32122 11511 32124
rect 11535 32122 11591 32124
rect 11615 32122 11671 32124
rect 11375 32070 11421 32122
rect 11421 32070 11431 32122
rect 11455 32070 11485 32122
rect 11485 32070 11497 32122
rect 11497 32070 11511 32122
rect 11535 32070 11549 32122
rect 11549 32070 11561 32122
rect 11561 32070 11591 32122
rect 11615 32070 11625 32122
rect 11625 32070 11671 32122
rect 11375 32068 11431 32070
rect 11455 32068 11511 32070
rect 11535 32068 11591 32070
rect 11615 32068 11671 32070
rect 18321 32122 18377 32124
rect 18401 32122 18457 32124
rect 18481 32122 18537 32124
rect 18561 32122 18617 32124
rect 18321 32070 18367 32122
rect 18367 32070 18377 32122
rect 18401 32070 18431 32122
rect 18431 32070 18443 32122
rect 18443 32070 18457 32122
rect 18481 32070 18495 32122
rect 18495 32070 18507 32122
rect 18507 32070 18537 32122
rect 18561 32070 18571 32122
rect 18571 32070 18617 32122
rect 18321 32068 18377 32070
rect 18401 32068 18457 32070
rect 18481 32068 18537 32070
rect 18561 32068 18617 32070
rect 25267 32122 25323 32124
rect 25347 32122 25403 32124
rect 25427 32122 25483 32124
rect 25507 32122 25563 32124
rect 25267 32070 25313 32122
rect 25313 32070 25323 32122
rect 25347 32070 25377 32122
rect 25377 32070 25389 32122
rect 25389 32070 25403 32122
rect 25427 32070 25441 32122
rect 25441 32070 25453 32122
rect 25453 32070 25483 32122
rect 25507 32070 25517 32122
rect 25517 32070 25563 32122
rect 25267 32068 25323 32070
rect 25347 32068 25403 32070
rect 25427 32068 25483 32070
rect 25507 32068 25563 32070
rect 1030 31048 1086 31104
rect 1582 29144 1638 29200
rect 1398 24928 1454 24984
rect 1306 21528 1362 21584
rect 754 19624 810 19680
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 2778 27240 2834 27296
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 3514 27648 3570 27704
rect 2778 23432 2834 23488
rect 3146 24656 3202 24712
rect 3514 24928 3570 24984
rect 754 15816 810 15872
rect 754 13932 810 13968
rect 754 13912 756 13932
rect 756 13912 808 13932
rect 808 13912 810 13932
rect 2134 18128 2190 18184
rect 2778 17720 2834 17776
rect 3054 17448 3110 17504
rect 3698 23432 3754 23488
rect 3514 18264 3570 18320
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4802 26424 4858 26480
rect 5262 26968 5318 27024
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 5170 26424 5226 26480
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4066 20848 4122 20904
rect 4894 21428 4896 21448
rect 4896 21428 4948 21448
rect 4948 21428 4950 21448
rect 4894 21392 4950 21428
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4618 20440 4674 20496
rect 4710 20304 4766 20360
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 5354 22344 5410 22400
rect 5538 23432 5594 23488
rect 5446 21684 5502 21720
rect 5446 21664 5448 21684
rect 5448 21664 5500 21684
rect 5500 21664 5502 21684
rect 5538 21548 5594 21584
rect 5538 21528 5540 21548
rect 5540 21528 5592 21548
rect 5592 21528 5594 21548
rect 5262 21392 5318 21448
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 754 12008 810 12064
rect 754 10104 810 10160
rect 1398 8200 1454 8256
rect 754 6316 810 6352
rect 754 6296 756 6316
rect 756 6296 808 6316
rect 808 6296 810 6316
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4986 17856 5042 17912
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4618 15136 4674 15192
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 5538 20304 5594 20360
rect 5722 21664 5778 21720
rect 5354 17332 5410 17368
rect 5630 17992 5686 18048
rect 5354 17312 5356 17332
rect 5356 17312 5408 17332
rect 5408 17312 5410 17332
rect 5170 13640 5226 13696
rect 5354 15136 5410 15192
rect 5906 21548 5962 21584
rect 5906 21528 5908 21548
rect 5908 21528 5960 21548
rect 5960 21528 5962 21548
rect 6366 23704 6422 23760
rect 6366 21972 6368 21992
rect 6368 21972 6420 21992
rect 6420 21972 6422 21992
rect 6366 21936 6422 21972
rect 6458 21392 6514 21448
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 7102 26424 7158 26480
rect 7378 26288 7434 26344
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 25870 30776 25926 30832
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 7654 26152 7710 26208
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7378 26016 7434 26072
rect 6734 21800 6790 21856
rect 6366 19352 6422 19408
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7654 21664 7710 21720
rect 7470 21392 7526 21448
rect 7286 21256 7342 21312
rect 7010 20712 7066 20768
rect 6550 18128 6606 18184
rect 8022 21936 8078 21992
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7838 20476 7840 20496
rect 7840 20476 7892 20496
rect 7892 20476 7894 20496
rect 7838 20440 7894 20476
rect 8482 21548 8538 21584
rect 8482 21528 8484 21548
rect 8484 21528 8536 21548
rect 8536 21528 8538 21548
rect 8666 21392 8722 21448
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7470 18264 7526 18320
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 4158 9560 4214 9616
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 754 4392 810 4448
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7102 16496 7158 16552
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 9126 21392 9182 21448
rect 9862 19796 9864 19816
rect 9864 19796 9916 19816
rect 9916 19796 9918 19816
rect 9862 19760 9918 19796
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 10322 19760 10378 19816
rect 10046 18400 10102 18456
rect 10046 18284 10102 18320
rect 10046 18264 10048 18284
rect 10048 18264 10100 18284
rect 10100 18264 10102 18284
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 9678 11328 9734 11384
rect 9770 11192 9826 11248
rect 10046 14900 10048 14920
rect 10048 14900 10100 14920
rect 10100 14900 10102 14920
rect 10046 14864 10102 14900
rect 9862 9036 9918 9072
rect 9862 9016 9864 9036
rect 9864 9016 9916 9036
rect 9916 9016 9918 9036
rect 10690 19352 10746 19408
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11794 20848 11850 20904
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11426 19388 11428 19408
rect 11428 19388 11480 19408
rect 11480 19388 11482 19408
rect 11426 19352 11482 19388
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 12806 23568 12862 23624
rect 12714 22344 12770 22400
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 10690 11348 10746 11384
rect 10690 11328 10692 11348
rect 10692 11328 10744 11348
rect 10744 11328 10746 11348
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11610 13368 11666 13424
rect 11058 10548 11060 10568
rect 11060 10548 11112 10568
rect 11112 10548 11114 10568
rect 11058 10512 11114 10548
rect 10598 9580 10654 9616
rect 10598 9560 10600 9580
rect 10600 9560 10652 9580
rect 10652 9560 10654 9580
rect 10598 9016 10654 9072
rect 10690 8900 10746 8936
rect 10690 8880 10692 8900
rect 10692 8880 10744 8900
rect 10744 8880 10746 8900
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 10966 8492 11022 8528
rect 10966 8472 10968 8492
rect 10968 8472 11020 8492
rect 11020 8472 11022 8492
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 12070 17176 12126 17232
rect 12254 17040 12310 17096
rect 12438 15156 12494 15192
rect 12438 15136 12440 15156
rect 12440 15136 12492 15156
rect 12492 15136 12494 15156
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 12162 12280 12218 12336
rect 12990 20848 13046 20904
rect 13174 21956 13230 21992
rect 13174 21936 13176 21956
rect 13176 21936 13228 21956
rect 13228 21936 13230 21956
rect 14922 27512 14978 27568
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 13542 20712 13598 20768
rect 14094 20748 14096 20768
rect 14096 20748 14148 20768
rect 14148 20748 14150 20768
rect 14094 20712 14150 20748
rect 13174 18400 13230 18456
rect 13542 18672 13598 18728
rect 13266 17196 13322 17232
rect 13266 17176 13268 17196
rect 13268 17176 13320 17196
rect 13320 17176 13322 17196
rect 12806 12688 12862 12744
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 4429 1658 4485 1660
rect 4509 1658 4565 1660
rect 4589 1658 4645 1660
rect 4669 1658 4725 1660
rect 4429 1606 4475 1658
rect 4475 1606 4485 1658
rect 4509 1606 4539 1658
rect 4539 1606 4551 1658
rect 4551 1606 4565 1658
rect 4589 1606 4603 1658
rect 4603 1606 4615 1658
rect 4615 1606 4645 1658
rect 4669 1606 4679 1658
rect 4679 1606 4725 1658
rect 4429 1604 4485 1606
rect 4509 1604 4565 1606
rect 4589 1604 4645 1606
rect 4669 1604 4725 1606
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 13726 17196 13782 17232
rect 13726 17176 13728 17196
rect 13728 17176 13780 17196
rect 13780 17176 13782 17196
rect 13818 16088 13874 16144
rect 13450 9596 13452 9616
rect 13452 9596 13504 9616
rect 13504 9596 13506 9616
rect 13450 9560 13506 9596
rect 12714 9016 12770 9072
rect 13358 9424 13414 9480
rect 12530 5652 12532 5672
rect 12532 5652 12584 5672
rect 12584 5652 12586 5672
rect 12530 5616 12586 5652
rect 13266 8880 13322 8936
rect 13450 7384 13506 7440
rect 12806 5616 12862 5672
rect 13450 4664 13506 4720
rect 14186 18128 14242 18184
rect 14094 17040 14150 17096
rect 14278 13368 14334 13424
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14922 19760 14978 19816
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 15474 19372 15530 19408
rect 15474 19352 15476 19372
rect 15476 19352 15528 19372
rect 15528 19352 15530 19372
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 15382 18400 15438 18456
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14922 15544 14978 15600
rect 16026 26288 16082 26344
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 16394 22924 16396 22944
rect 16396 22924 16448 22944
rect 16448 22924 16450 22944
rect 16394 22888 16450 22924
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 16670 22072 16726 22128
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 15750 17992 15806 18048
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14738 14456 14794 14512
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 14370 12280 14426 12336
rect 14462 11192 14518 11248
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 15566 15408 15622 15464
rect 15474 15272 15530 15328
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 15290 9596 15292 9616
rect 15292 9596 15344 9616
rect 15344 9596 15346 9616
rect 15290 9560 15346 9596
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 11375 1658 11431 1660
rect 11455 1658 11511 1660
rect 11535 1658 11591 1660
rect 11615 1658 11671 1660
rect 11375 1606 11421 1658
rect 11421 1606 11431 1658
rect 11455 1606 11485 1658
rect 11485 1606 11497 1658
rect 11497 1606 11511 1658
rect 11535 1606 11549 1658
rect 11549 1606 11561 1658
rect 11561 1606 11591 1658
rect 11615 1606 11625 1658
rect 11625 1606 11671 1658
rect 11375 1604 11431 1606
rect 11455 1604 11511 1606
rect 11535 1604 11591 1606
rect 11615 1604 11671 1606
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 15934 15544 15990 15600
rect 15842 12824 15898 12880
rect 16118 15408 16174 15464
rect 16670 21528 16726 21584
rect 16394 14476 16450 14512
rect 16394 14456 16396 14476
rect 16396 14456 16448 14476
rect 16448 14456 16450 14476
rect 16394 14320 16450 14376
rect 16670 16532 16672 16552
rect 16672 16532 16724 16552
rect 16724 16532 16726 16552
rect 16670 16496 16726 16532
rect 16578 13640 16634 13696
rect 15750 11056 15806 11112
rect 15658 8472 15714 8528
rect 16118 8880 16174 8936
rect 15842 8200 15898 8256
rect 15290 5616 15346 5672
rect 16026 8472 16082 8528
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 16210 8744 16266 8800
rect 16854 16632 16910 16688
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 17314 18672 17370 18728
rect 17130 14864 17186 14920
rect 17406 18264 17462 18320
rect 17406 18128 17462 18184
rect 17498 16088 17554 16144
rect 16946 12588 16948 12608
rect 16948 12588 17000 12608
rect 17000 12588 17002 12608
rect 16946 12552 17002 12588
rect 17314 13368 17370 13424
rect 17682 21120 17738 21176
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 17682 13640 17738 13696
rect 17222 13096 17278 13152
rect 16486 8508 16488 8528
rect 16488 8508 16540 8528
rect 16540 8508 16542 8528
rect 16486 8472 16542 8508
rect 16394 7248 16450 7304
rect 17038 9016 17094 9072
rect 17038 7384 17094 7440
rect 16946 6840 17002 6896
rect 17682 9560 17738 9616
rect 17774 8744 17830 8800
rect 18602 19352 18658 19408
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18234 18400 18290 18456
rect 19982 23468 19984 23488
rect 19984 23468 20036 23488
rect 20036 23468 20038 23488
rect 19982 23432 20038 23468
rect 19614 23160 19670 23216
rect 19706 22208 19762 22264
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 19430 19216 19486 19272
rect 19062 18400 19118 18456
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18510 16108 18566 16144
rect 18510 16088 18512 16108
rect 18512 16088 18564 16108
rect 18564 16088 18566 16108
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 19338 17876 19394 17912
rect 19338 17856 19349 17876
rect 19349 17856 19394 17876
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 20166 22208 20222 22264
rect 19982 20748 19984 20768
rect 19984 20748 20036 20768
rect 20036 20748 20038 20768
rect 19982 20712 20038 20748
rect 19982 19624 20038 19680
rect 19982 19216 20038 19272
rect 19430 16396 19432 16416
rect 19432 16396 19484 16416
rect 19484 16396 19486 16416
rect 19430 16360 19486 16396
rect 19338 15000 19394 15056
rect 19246 12824 19302 12880
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18326 10548 18328 10568
rect 18328 10548 18380 10568
rect 18380 10548 18382 10568
rect 18326 10512 18382 10548
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 17958 6840 18014 6896
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 17866 5652 17868 5672
rect 17868 5652 17920 5672
rect 17920 5652 17922 5672
rect 17866 5616 17922 5652
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 20074 18264 20130 18320
rect 20718 19624 20774 19680
rect 20626 18672 20682 18728
rect 20534 16396 20536 16416
rect 20536 16396 20588 16416
rect 20588 16396 20590 16416
rect 20534 16360 20590 16396
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 19982 12316 19984 12336
rect 19984 12316 20036 12336
rect 20036 12316 20038 12336
rect 19982 12280 20038 12316
rect 19982 10648 20038 10704
rect 19154 4664 19210 4720
rect 20902 18400 20958 18456
rect 20994 15428 21050 15464
rect 20994 15408 20996 15428
rect 20996 15408 21048 15428
rect 21048 15408 21050 15428
rect 20350 11756 20406 11792
rect 20350 11736 20352 11756
rect 20352 11736 20404 11756
rect 20404 11736 20406 11756
rect 20442 9696 20498 9752
rect 20718 12824 20774 12880
rect 20534 7928 20590 7984
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 18321 1658 18377 1660
rect 18401 1658 18457 1660
rect 18481 1658 18537 1660
rect 18561 1658 18617 1660
rect 18321 1606 18367 1658
rect 18367 1606 18377 1658
rect 18401 1606 18431 1658
rect 18431 1606 18443 1658
rect 18443 1606 18457 1658
rect 18481 1606 18495 1658
rect 18495 1606 18507 1658
rect 18507 1606 18537 1658
rect 18561 1606 18571 1658
rect 18571 1606 18617 1658
rect 18321 1604 18377 1606
rect 18401 1604 18457 1606
rect 18481 1604 18537 1606
rect 18561 1604 18617 1606
rect 20902 12280 20958 12336
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21546 17856 21602 17912
rect 21362 13252 21418 13288
rect 21362 13232 21364 13252
rect 21364 13232 21416 13252
rect 21416 13232 21418 13252
rect 21178 12280 21234 12336
rect 21178 12008 21234 12064
rect 21454 11872 21510 11928
rect 21822 18672 21878 18728
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21914 18164 21916 18184
rect 21916 18164 21968 18184
rect 21968 18164 21970 18184
rect 21914 18128 21970 18164
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 22374 18808 22430 18864
rect 22282 18264 22338 18320
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 22834 23196 22836 23216
rect 22836 23196 22888 23216
rect 22888 23196 22890 23216
rect 22834 23160 22890 23196
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 25870 25880 25926 25936
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21730 14864 21786 14920
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 22282 13232 22338 13288
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 22006 11772 22008 11792
rect 22008 11772 22060 11792
rect 22060 11772 22062 11792
rect 22006 11736 22062 11772
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 22006 9596 22008 9616
rect 22008 9596 22060 9616
rect 22060 9596 22062 9616
rect 22006 9560 22062 9596
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 22190 8472 22246 8528
rect 21546 8336 21602 8392
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 22742 18264 22798 18320
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 22926 18028 22928 18048
rect 22928 18028 22980 18048
rect 22980 18028 22982 18048
rect 22926 17992 22982 18028
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25134 21528 25190 21584
rect 23110 18128 23166 18184
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 23662 16632 23718 16688
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25778 18672 25834 18728
rect 25686 16904 25742 16960
rect 23478 15272 23534 15328
rect 24766 15444 24768 15464
rect 24768 15444 24820 15464
rect 24820 15444 24822 15464
rect 24766 15408 24822 15444
rect 23018 10104 23074 10160
rect 22650 8744 22706 8800
rect 22650 7248 22706 7304
rect 23018 9560 23074 9616
rect 23294 10648 23350 10704
rect 22926 5480 22982 5536
rect 23662 8744 23718 8800
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 24398 12824 24454 12880
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 23846 8336 23902 8392
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 25778 12280 25834 12336
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 27618 13404 27620 13424
rect 27620 13404 27672 13424
rect 27672 13404 27674 13424
rect 27618 13368 27674 13404
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 27618 10104 27674 10160
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25870 7792 25926 7848
rect 26606 7928 26662 7984
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 25870 3032 25926 3088
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 25267 1658 25323 1660
rect 25347 1658 25403 1660
rect 25427 1658 25483 1660
rect 25507 1658 25563 1660
rect 25267 1606 25313 1658
rect 25313 1606 25323 1658
rect 25347 1606 25377 1658
rect 25377 1606 25389 1658
rect 25389 1606 25403 1658
rect 25427 1606 25441 1658
rect 25441 1606 25453 1658
rect 25453 1606 25483 1658
rect 25507 1606 25517 1658
rect 25517 1606 25563 1658
rect 25267 1604 25323 1606
rect 25347 1604 25403 1606
rect 25427 1604 25483 1606
rect 25507 1604 25563 1606
rect 7902 1114 7958 1116
rect 7982 1114 8038 1116
rect 8062 1114 8118 1116
rect 8142 1114 8198 1116
rect 7902 1062 7948 1114
rect 7948 1062 7958 1114
rect 7982 1062 8012 1114
rect 8012 1062 8024 1114
rect 8024 1062 8038 1114
rect 8062 1062 8076 1114
rect 8076 1062 8088 1114
rect 8088 1062 8118 1114
rect 8142 1062 8152 1114
rect 8152 1062 8198 1114
rect 7902 1060 7958 1062
rect 7982 1060 8038 1062
rect 8062 1060 8118 1062
rect 8142 1060 8198 1062
rect 14848 1114 14904 1116
rect 14928 1114 14984 1116
rect 15008 1114 15064 1116
rect 15088 1114 15144 1116
rect 14848 1062 14894 1114
rect 14894 1062 14904 1114
rect 14928 1062 14958 1114
rect 14958 1062 14970 1114
rect 14970 1062 14984 1114
rect 15008 1062 15022 1114
rect 15022 1062 15034 1114
rect 15034 1062 15064 1114
rect 15088 1062 15098 1114
rect 15098 1062 15144 1114
rect 14848 1060 14904 1062
rect 14928 1060 14984 1062
rect 15008 1060 15064 1062
rect 15088 1060 15144 1062
rect 21794 1114 21850 1116
rect 21874 1114 21930 1116
rect 21954 1114 22010 1116
rect 22034 1114 22090 1116
rect 21794 1062 21840 1114
rect 21840 1062 21850 1114
rect 21874 1062 21904 1114
rect 21904 1062 21916 1114
rect 21916 1062 21930 1114
rect 21954 1062 21968 1114
rect 21968 1062 21980 1114
rect 21980 1062 22010 1114
rect 22034 1062 22044 1114
rect 22044 1062 22090 1114
rect 21794 1060 21850 1062
rect 21874 1060 21930 1062
rect 21954 1060 22010 1062
rect 22034 1060 22090 1062
rect 28740 1114 28796 1116
rect 28820 1114 28876 1116
rect 28900 1114 28956 1116
rect 28980 1114 29036 1116
rect 28740 1062 28786 1114
rect 28786 1062 28796 1114
rect 28820 1062 28850 1114
rect 28850 1062 28862 1114
rect 28862 1062 28876 1114
rect 28900 1062 28914 1114
rect 28914 1062 28926 1114
rect 28926 1062 28956 1114
rect 28980 1062 28990 1114
rect 28990 1062 29036 1114
rect 28740 1060 28796 1062
rect 28820 1060 28876 1062
rect 28900 1060 28956 1062
rect 28980 1060 29036 1062
<< metal3 >>
rect 7892 32672 8208 32673
rect 7892 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8208 32672
rect 7892 32607 8208 32608
rect 14838 32672 15154 32673
rect 14838 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15154 32672
rect 14838 32607 15154 32608
rect 21784 32672 22100 32673
rect 21784 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22100 32672
rect 21784 32607 22100 32608
rect 28730 32672 29046 32673
rect 28730 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29046 32672
rect 28730 32607 29046 32608
rect 4419 32128 4735 32129
rect 4419 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4735 32128
rect 4419 32063 4735 32064
rect 11365 32128 11681 32129
rect 11365 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11681 32128
rect 11365 32063 11681 32064
rect 18311 32128 18627 32129
rect 18311 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18627 32128
rect 18311 32063 18627 32064
rect 25257 32128 25573 32129
rect 25257 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25573 32128
rect 25257 32063 25573 32064
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 0 31106 400 31136
rect 1025 31106 1091 31109
rect 0 31104 1091 31106
rect 0 31048 1030 31104
rect 1086 31048 1091 31104
rect 0 31046 1091 31048
rect 0 31016 400 31046
rect 1025 31043 1091 31046
rect 4419 31040 4735 31041
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 25865 30834 25931 30837
rect 29600 30834 30000 30864
rect 25865 30832 30000 30834
rect 25865 30776 25870 30832
rect 25926 30776 30000 30832
rect 25865 30774 30000 30776
rect 25865 30771 25931 30774
rect 29600 30744 30000 30774
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 28730 30431 29046 30432
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 0 29202 400 29232
rect 1577 29202 1643 29205
rect 0 29200 1643 29202
rect 0 29144 1582 29200
rect 1638 29144 1643 29200
rect 0 29142 1643 29144
rect 0 29112 400 29142
rect 1577 29139 1643 29142
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 7892 28320 8208 28321
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 3509 27706 3575 27709
rect 3734 27706 3740 27708
rect 3509 27704 3740 27706
rect 3509 27648 3514 27704
rect 3570 27648 3740 27704
rect 3509 27646 3740 27648
rect 3509 27643 3575 27646
rect 3734 27644 3740 27646
rect 3804 27644 3810 27708
rect 14917 27570 14983 27573
rect 16430 27570 16436 27572
rect 14917 27568 16436 27570
rect 14917 27512 14922 27568
rect 14978 27512 16436 27568
rect 14917 27510 16436 27512
rect 14917 27507 14983 27510
rect 16430 27508 16436 27510
rect 16500 27508 16506 27572
rect 0 27298 400 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 400 27238
rect 2773 27235 2839 27238
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 5022 26964 5028 27028
rect 5092 27026 5098 27028
rect 5257 27026 5323 27029
rect 5092 27024 5323 27026
rect 5092 26968 5262 27024
rect 5318 26968 5323 27024
rect 5092 26966 5323 26968
rect 5092 26964 5098 26966
rect 5257 26963 5323 26966
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 4797 26482 4863 26485
rect 5165 26482 5231 26485
rect 7097 26482 7163 26485
rect 4797 26480 7163 26482
rect 4797 26424 4802 26480
rect 4858 26424 5170 26480
rect 5226 26424 7102 26480
rect 7158 26424 7163 26480
rect 4797 26422 7163 26424
rect 4797 26419 4863 26422
rect 5165 26419 5231 26422
rect 7097 26419 7163 26422
rect 7230 26284 7236 26348
rect 7300 26346 7306 26348
rect 7373 26346 7439 26349
rect 7300 26344 7439 26346
rect 7300 26288 7378 26344
rect 7434 26288 7439 26344
rect 7300 26286 7439 26288
rect 7300 26284 7306 26286
rect 7373 26283 7439 26286
rect 16021 26346 16087 26349
rect 21214 26346 21220 26348
rect 16021 26344 21220 26346
rect 16021 26288 16026 26344
rect 16082 26288 21220 26344
rect 16021 26286 21220 26288
rect 16021 26283 16087 26286
rect 21214 26284 21220 26286
rect 21284 26284 21290 26348
rect 6678 26148 6684 26212
rect 6748 26210 6754 26212
rect 7649 26210 7715 26213
rect 29600 26210 30000 26240
rect 6748 26208 7715 26210
rect 6748 26152 7654 26208
rect 7710 26152 7715 26208
rect 6748 26150 7715 26152
rect 6748 26148 6754 26150
rect 7649 26147 7715 26150
rect 29134 26150 30000 26210
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 7373 26076 7439 26077
rect 7373 26074 7420 26076
rect 7328 26072 7420 26074
rect 7328 26016 7378 26072
rect 7328 26014 7420 26016
rect 7373 26012 7420 26014
rect 7484 26012 7490 26076
rect 7373 26011 7439 26012
rect 25865 25938 25931 25941
rect 29134 25938 29194 26150
rect 29600 26120 30000 26150
rect 25865 25936 29194 25938
rect 25865 25880 25870 25936
rect 25926 25880 29194 25936
rect 25865 25878 29194 25880
rect 25865 25875 25931 25878
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 0 25394 400 25424
rect 0 25334 858 25394
rect 0 25304 400 25334
rect 798 24986 858 25334
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 1393 24986 1459 24989
rect 798 24984 1459 24986
rect 798 24928 1398 24984
rect 1454 24928 1459 24984
rect 798 24926 1459 24928
rect 1393 24923 1459 24926
rect 3509 24988 3575 24989
rect 3509 24984 3556 24988
rect 3620 24986 3626 24988
rect 3509 24928 3514 24984
rect 3509 24924 3556 24928
rect 3620 24926 3666 24986
rect 3620 24924 3626 24926
rect 3509 24923 3575 24924
rect 3141 24714 3207 24717
rect 4838 24714 4844 24716
rect 3141 24712 4844 24714
rect 3141 24656 3146 24712
rect 3202 24656 4844 24712
rect 3141 24654 4844 24656
rect 3141 24651 3207 24654
rect 4838 24652 4844 24654
rect 4908 24652 4914 24716
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 6361 23764 6427 23765
rect 6310 23700 6316 23764
rect 6380 23762 6427 23764
rect 6380 23760 6472 23762
rect 6422 23704 6472 23760
rect 6380 23702 6472 23704
rect 6380 23700 6427 23702
rect 6361 23699 6427 23700
rect 12801 23628 12867 23629
rect 12750 23564 12756 23628
rect 12820 23626 12867 23628
rect 12820 23624 12912 23626
rect 12862 23568 12912 23624
rect 12820 23566 12912 23568
rect 12820 23564 12867 23566
rect 12801 23563 12867 23564
rect 0 23490 400 23520
rect 2773 23490 2839 23493
rect 3693 23492 3759 23493
rect 3693 23490 3740 23492
rect 0 23488 2839 23490
rect 0 23432 2778 23488
rect 2834 23432 2839 23488
rect 0 23430 2839 23432
rect 3648 23488 3740 23490
rect 3648 23432 3698 23488
rect 3648 23430 3740 23432
rect 0 23400 400 23430
rect 2773 23427 2839 23430
rect 3693 23428 3740 23430
rect 3804 23428 3810 23492
rect 5533 23490 5599 23493
rect 19977 23492 20043 23493
rect 7598 23490 7604 23492
rect 5533 23488 7604 23490
rect 5533 23432 5538 23488
rect 5594 23432 7604 23488
rect 5533 23430 7604 23432
rect 3693 23427 3759 23428
rect 5533 23427 5599 23430
rect 7598 23428 7604 23430
rect 7668 23428 7674 23492
rect 19926 23490 19932 23492
rect 19886 23430 19932 23490
rect 19996 23488 20043 23492
rect 20038 23432 20043 23488
rect 19926 23428 19932 23430
rect 19996 23428 20043 23432
rect 19977 23427 20043 23428
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 19609 23218 19675 23221
rect 22829 23218 22895 23221
rect 19609 23216 22895 23218
rect 19609 23160 19614 23216
rect 19670 23160 22834 23216
rect 22890 23160 22895 23216
rect 19609 23158 22895 23160
rect 19609 23155 19675 23158
rect 22829 23155 22895 23158
rect 16389 22948 16455 22949
rect 16389 22946 16436 22948
rect 16344 22944 16436 22946
rect 16344 22888 16394 22944
rect 16344 22886 16436 22888
rect 16389 22884 16436 22886
rect 16500 22884 16506 22948
rect 16389 22883 16455 22884
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 5349 22404 5415 22405
rect 5349 22400 5396 22404
rect 5460 22402 5466 22404
rect 5349 22344 5354 22400
rect 5349 22340 5396 22344
rect 5460 22342 5506 22402
rect 5460 22340 5466 22342
rect 12566 22340 12572 22404
rect 12636 22402 12642 22404
rect 12709 22402 12775 22405
rect 12636 22400 12775 22402
rect 12636 22344 12714 22400
rect 12770 22344 12775 22400
rect 12636 22342 12775 22344
rect 12636 22340 12642 22342
rect 5349 22339 5415 22340
rect 12709 22339 12775 22342
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 19701 22266 19767 22269
rect 20161 22266 20227 22269
rect 19701 22264 20227 22266
rect 19701 22208 19706 22264
rect 19762 22208 20166 22264
rect 20222 22208 20227 22264
rect 19701 22206 20227 22208
rect 19701 22203 19767 22206
rect 20161 22203 20227 22206
rect 16665 22130 16731 22133
rect 16622 22128 16731 22130
rect 16622 22072 16670 22128
rect 16726 22072 16731 22128
rect 16622 22067 16731 22072
rect 6361 21996 6427 21997
rect 6310 21994 6316 21996
rect 6270 21934 6316 21994
rect 6380 21992 6427 21996
rect 6422 21936 6427 21992
rect 6310 21932 6316 21934
rect 6380 21932 6427 21936
rect 6361 21931 6427 21932
rect 8017 21994 8083 21997
rect 13169 21994 13235 21997
rect 16622 21994 16682 22067
rect 8017 21992 8402 21994
rect 8017 21936 8022 21992
rect 8078 21936 8402 21992
rect 8017 21934 8402 21936
rect 8017 21931 8083 21934
rect 6729 21860 6795 21861
rect 6678 21858 6684 21860
rect 6638 21798 6684 21858
rect 6748 21856 6795 21860
rect 6790 21800 6795 21856
rect 6678 21796 6684 21798
rect 6748 21796 6795 21800
rect 6729 21795 6795 21796
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 5441 21722 5507 21725
rect 5717 21722 5783 21725
rect 7649 21724 7715 21725
rect 5441 21720 5783 21722
rect 5441 21664 5446 21720
rect 5502 21664 5722 21720
rect 5778 21664 5783 21720
rect 5441 21662 5783 21664
rect 5441 21659 5507 21662
rect 5717 21659 5783 21662
rect 7598 21660 7604 21724
rect 7668 21722 7715 21724
rect 7668 21720 7760 21722
rect 7710 21664 7760 21720
rect 7668 21662 7760 21664
rect 7668 21660 7715 21662
rect 7649 21659 7715 21660
rect 0 21586 400 21616
rect 1301 21586 1367 21589
rect 0 21584 1367 21586
rect 0 21528 1306 21584
rect 1362 21528 1367 21584
rect 0 21526 1367 21528
rect 0 21496 400 21526
rect 1301 21523 1367 21526
rect 5533 21586 5599 21589
rect 5901 21586 5967 21589
rect 5533 21584 5967 21586
rect 5533 21528 5538 21584
rect 5594 21528 5906 21584
rect 5962 21528 5967 21584
rect 5533 21526 5967 21528
rect 8342 21586 8402 21934
rect 13169 21992 16682 21994
rect 13169 21936 13174 21992
rect 13230 21936 16682 21992
rect 13169 21934 16682 21936
rect 13169 21931 13235 21934
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 16622 21589 16682 21934
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 8477 21586 8543 21589
rect 8342 21584 8543 21586
rect 8342 21528 8482 21584
rect 8538 21528 8543 21584
rect 8342 21526 8543 21528
rect 16622 21584 16731 21589
rect 16622 21528 16670 21584
rect 16726 21528 16731 21584
rect 16622 21526 16731 21528
rect 5533 21523 5599 21526
rect 5901 21523 5967 21526
rect 8477 21523 8543 21526
rect 16665 21523 16731 21526
rect 25129 21586 25195 21589
rect 29600 21586 30000 21616
rect 25129 21584 30000 21586
rect 25129 21528 25134 21584
rect 25190 21528 30000 21584
rect 25129 21526 30000 21528
rect 25129 21523 25195 21526
rect 29600 21496 30000 21526
rect 4889 21452 4955 21453
rect 4838 21388 4844 21452
rect 4908 21450 4955 21452
rect 5257 21450 5323 21453
rect 6453 21450 6519 21453
rect 4908 21448 5000 21450
rect 4950 21392 5000 21448
rect 4908 21390 5000 21392
rect 5257 21448 6519 21450
rect 5257 21392 5262 21448
rect 5318 21392 6458 21448
rect 6514 21392 6519 21448
rect 5257 21390 6519 21392
rect 4908 21388 4955 21390
rect 4889 21387 4955 21388
rect 5257 21387 5323 21390
rect 6453 21387 6519 21390
rect 7230 21388 7236 21452
rect 7300 21450 7306 21452
rect 7465 21450 7531 21453
rect 7300 21448 7531 21450
rect 7300 21392 7470 21448
rect 7526 21392 7531 21448
rect 7300 21390 7531 21392
rect 7300 21388 7306 21390
rect 7465 21387 7531 21390
rect 8661 21450 8727 21453
rect 9121 21450 9187 21453
rect 8661 21448 9187 21450
rect 8661 21392 8666 21448
rect 8722 21392 9126 21448
rect 9182 21392 9187 21448
rect 8661 21390 9187 21392
rect 8661 21387 8727 21390
rect 9121 21387 9187 21390
rect 7281 21314 7347 21317
rect 7414 21314 7420 21316
rect 7281 21312 7420 21314
rect 7281 21256 7286 21312
rect 7342 21256 7420 21312
rect 7281 21254 7420 21256
rect 7281 21251 7347 21254
rect 7414 21252 7420 21254
rect 7484 21252 7490 21316
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 17534 21116 17540 21180
rect 17604 21178 17610 21180
rect 17677 21178 17743 21181
rect 17604 21176 17743 21178
rect 17604 21120 17682 21176
rect 17738 21120 17743 21176
rect 17604 21118 17743 21120
rect 17604 21116 17610 21118
rect 17677 21115 17743 21118
rect 4061 20906 4127 20909
rect 11789 20906 11855 20909
rect 12985 20906 13051 20909
rect 4061 20904 13051 20906
rect 4061 20848 4066 20904
rect 4122 20848 11794 20904
rect 11850 20848 12990 20904
rect 13046 20848 13051 20904
rect 4061 20846 13051 20848
rect 4061 20843 4127 20846
rect 11789 20843 11855 20846
rect 12985 20843 13051 20846
rect 6862 20708 6868 20772
rect 6932 20770 6938 20772
rect 7005 20770 7071 20773
rect 6932 20768 7071 20770
rect 6932 20712 7010 20768
rect 7066 20712 7071 20768
rect 6932 20710 7071 20712
rect 6932 20708 6938 20710
rect 7005 20707 7071 20710
rect 13537 20770 13603 20773
rect 13670 20770 13676 20772
rect 13537 20768 13676 20770
rect 13537 20712 13542 20768
rect 13598 20712 13676 20768
rect 13537 20710 13676 20712
rect 13537 20707 13603 20710
rect 13670 20708 13676 20710
rect 13740 20708 13746 20772
rect 14089 20770 14155 20773
rect 14222 20770 14228 20772
rect 14089 20768 14228 20770
rect 14089 20712 14094 20768
rect 14150 20712 14228 20768
rect 14089 20710 14228 20712
rect 14089 20707 14155 20710
rect 14222 20708 14228 20710
rect 14292 20708 14298 20772
rect 19977 20770 20043 20773
rect 20110 20770 20116 20772
rect 19977 20768 20116 20770
rect 19977 20712 19982 20768
rect 20038 20712 20116 20768
rect 19977 20710 20116 20712
rect 19977 20707 20043 20710
rect 20110 20708 20116 20710
rect 20180 20708 20186 20772
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 4613 20498 4679 20501
rect 7833 20498 7899 20501
rect 4613 20496 7899 20498
rect 4613 20440 4618 20496
rect 4674 20440 7838 20496
rect 7894 20440 7899 20496
rect 4613 20438 7899 20440
rect 4613 20435 4679 20438
rect 7833 20435 7899 20438
rect 4705 20362 4771 20365
rect 5533 20362 5599 20365
rect 4705 20360 5599 20362
rect 4705 20304 4710 20360
rect 4766 20304 5538 20360
rect 5594 20304 5599 20360
rect 4705 20302 5599 20304
rect 4705 20299 4771 20302
rect 5533 20299 5599 20302
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 9857 19818 9923 19821
rect 10317 19818 10383 19821
rect 9857 19816 10383 19818
rect 9857 19760 9862 19816
rect 9918 19760 10322 19816
rect 10378 19760 10383 19816
rect 9857 19758 10383 19760
rect 9857 19755 9923 19758
rect 10317 19755 10383 19758
rect 14590 19756 14596 19820
rect 14660 19818 14666 19820
rect 14917 19818 14983 19821
rect 14660 19816 14983 19818
rect 14660 19760 14922 19816
rect 14978 19760 14983 19816
rect 14660 19758 14983 19760
rect 14660 19756 14666 19758
rect 14917 19755 14983 19758
rect 0 19682 400 19712
rect 749 19682 815 19685
rect 0 19680 815 19682
rect 0 19624 754 19680
rect 810 19624 815 19680
rect 0 19622 815 19624
rect 0 19592 400 19622
rect 749 19619 815 19622
rect 19977 19682 20043 19685
rect 20713 19682 20779 19685
rect 19977 19680 20779 19682
rect 19977 19624 19982 19680
rect 20038 19624 20718 19680
rect 20774 19624 20779 19680
rect 19977 19622 20779 19624
rect 19977 19619 20043 19622
rect 20713 19619 20779 19622
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 6361 19410 6427 19413
rect 6494 19410 6500 19412
rect 6361 19408 6500 19410
rect 6361 19352 6366 19408
rect 6422 19352 6500 19408
rect 6361 19350 6500 19352
rect 6361 19347 6427 19350
rect 6494 19348 6500 19350
rect 6564 19348 6570 19412
rect 10685 19410 10751 19413
rect 11421 19410 11487 19413
rect 10685 19408 11487 19410
rect 10685 19352 10690 19408
rect 10746 19352 11426 19408
rect 11482 19352 11487 19408
rect 10685 19350 11487 19352
rect 10685 19347 10751 19350
rect 11421 19347 11487 19350
rect 15469 19410 15535 19413
rect 18597 19410 18663 19413
rect 15469 19408 18663 19410
rect 15469 19352 15474 19408
rect 15530 19352 18602 19408
rect 18658 19352 18663 19408
rect 15469 19350 18663 19352
rect 15469 19347 15535 19350
rect 18597 19347 18663 19350
rect 19425 19274 19491 19277
rect 19977 19274 20043 19277
rect 19425 19272 20043 19274
rect 19425 19216 19430 19272
rect 19486 19216 19982 19272
rect 20038 19216 20043 19272
rect 19425 19214 20043 19216
rect 19425 19211 19491 19214
rect 19977 19211 20043 19214
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 21214 18804 21220 18868
rect 21284 18866 21290 18868
rect 22369 18866 22435 18869
rect 21284 18864 22435 18866
rect 21284 18808 22374 18864
rect 22430 18808 22435 18864
rect 21284 18806 22435 18808
rect 21284 18804 21290 18806
rect 22369 18803 22435 18806
rect 13537 18730 13603 18733
rect 17309 18730 17375 18733
rect 13537 18728 17375 18730
rect 13537 18672 13542 18728
rect 13598 18672 17314 18728
rect 17370 18672 17375 18728
rect 13537 18670 17375 18672
rect 13537 18667 13603 18670
rect 17309 18667 17375 18670
rect 20621 18730 20687 18733
rect 21817 18730 21883 18733
rect 25773 18730 25839 18733
rect 20621 18728 25839 18730
rect 20621 18672 20626 18728
rect 20682 18672 21822 18728
rect 21878 18672 25778 18728
rect 25834 18672 25839 18728
rect 20621 18670 25839 18672
rect 20621 18667 20687 18670
rect 21817 18667 21883 18670
rect 25773 18667 25839 18670
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 10041 18458 10107 18461
rect 13169 18458 13235 18461
rect 10041 18456 13235 18458
rect 10041 18400 10046 18456
rect 10102 18400 13174 18456
rect 13230 18400 13235 18456
rect 10041 18398 13235 18400
rect 10041 18395 10107 18398
rect 13169 18395 13235 18398
rect 15377 18458 15443 18461
rect 18229 18458 18295 18461
rect 15377 18456 18295 18458
rect 15377 18400 15382 18456
rect 15438 18400 18234 18456
rect 18290 18400 18295 18456
rect 15377 18398 18295 18400
rect 15377 18395 15443 18398
rect 18229 18395 18295 18398
rect 19057 18458 19123 18461
rect 20897 18458 20963 18461
rect 19057 18456 20963 18458
rect 19057 18400 19062 18456
rect 19118 18400 20902 18456
rect 20958 18400 20963 18456
rect 19057 18398 20963 18400
rect 19057 18395 19123 18398
rect 20897 18395 20963 18398
rect 3509 18322 3575 18325
rect 7465 18322 7531 18325
rect 3509 18320 7531 18322
rect 3509 18264 3514 18320
rect 3570 18264 7470 18320
rect 7526 18264 7531 18320
rect 3509 18262 7531 18264
rect 3509 18259 3575 18262
rect 7465 18259 7531 18262
rect 10041 18322 10107 18325
rect 17401 18322 17467 18325
rect 10041 18320 17467 18322
rect 10041 18264 10046 18320
rect 10102 18264 17406 18320
rect 17462 18264 17467 18320
rect 10041 18262 17467 18264
rect 10041 18259 10107 18262
rect 17401 18259 17467 18262
rect 20069 18322 20135 18325
rect 22277 18322 22343 18325
rect 22737 18324 22803 18325
rect 22686 18322 22692 18324
rect 20069 18320 22343 18322
rect 20069 18264 20074 18320
rect 20130 18264 22282 18320
rect 22338 18264 22343 18320
rect 20069 18262 22343 18264
rect 22646 18262 22692 18322
rect 22756 18320 22803 18324
rect 22798 18264 22803 18320
rect 20069 18259 20135 18262
rect 22277 18259 22343 18262
rect 22686 18260 22692 18262
rect 22756 18260 22803 18264
rect 22737 18259 22803 18260
rect 2129 18186 2195 18189
rect 6545 18186 6611 18189
rect 2129 18184 6611 18186
rect 2129 18128 2134 18184
rect 2190 18128 6550 18184
rect 6606 18128 6611 18184
rect 2129 18126 6611 18128
rect 2129 18123 2195 18126
rect 6545 18123 6611 18126
rect 14181 18186 14247 18189
rect 17401 18186 17467 18189
rect 14181 18184 17467 18186
rect 14181 18128 14186 18184
rect 14242 18128 17406 18184
rect 17462 18128 17467 18184
rect 14181 18126 17467 18128
rect 14181 18123 14247 18126
rect 17401 18123 17467 18126
rect 21909 18186 21975 18189
rect 23105 18186 23171 18189
rect 21909 18184 23171 18186
rect 21909 18128 21914 18184
rect 21970 18128 23110 18184
rect 23166 18128 23171 18184
rect 21909 18126 23171 18128
rect 21909 18123 21975 18126
rect 23105 18123 23171 18126
rect 5625 18052 5691 18053
rect 5574 18050 5580 18052
rect 5534 17990 5580 18050
rect 5644 18048 5691 18052
rect 5686 17992 5691 18048
rect 5574 17988 5580 17990
rect 5644 17988 5691 17992
rect 15510 17988 15516 18052
rect 15580 18050 15586 18052
rect 15745 18050 15811 18053
rect 15580 18048 15811 18050
rect 15580 17992 15750 18048
rect 15806 17992 15811 18048
rect 15580 17990 15811 17992
rect 15580 17988 15586 17990
rect 5625 17987 5691 17988
rect 15745 17987 15811 17990
rect 22921 18050 22987 18053
rect 23054 18050 23060 18052
rect 22921 18048 23060 18050
rect 22921 17992 22926 18048
rect 22982 17992 23060 18048
rect 22921 17990 23060 17992
rect 22921 17987 22987 17990
rect 23054 17988 23060 17990
rect 23124 17988 23130 18052
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 4838 17852 4844 17916
rect 4908 17914 4914 17916
rect 4981 17914 5047 17917
rect 4908 17912 5047 17914
rect 4908 17856 4986 17912
rect 5042 17856 5047 17912
rect 4908 17854 5047 17856
rect 4908 17852 4914 17854
rect 4981 17851 5047 17854
rect 19333 17914 19399 17917
rect 21541 17914 21607 17917
rect 19333 17912 21607 17914
rect 19333 17856 19338 17912
rect 19394 17856 21546 17912
rect 21602 17856 21607 17912
rect 19333 17854 21607 17856
rect 19333 17851 19399 17854
rect 21541 17851 21607 17854
rect 0 17778 400 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 400 17718
rect 2773 17715 2839 17718
rect 3049 17506 3115 17509
rect 6862 17506 6868 17508
rect 3049 17504 6868 17506
rect 3049 17448 3054 17504
rect 3110 17448 6868 17504
rect 3049 17446 6868 17448
rect 3049 17443 3115 17446
rect 6862 17444 6868 17446
rect 6932 17444 6938 17508
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 5349 17372 5415 17373
rect 5349 17370 5396 17372
rect 5304 17368 5396 17370
rect 5304 17312 5354 17368
rect 5304 17310 5396 17312
rect 5349 17308 5396 17310
rect 5460 17308 5466 17372
rect 5349 17307 5415 17308
rect 12065 17234 12131 17237
rect 13261 17234 13327 17237
rect 13721 17234 13787 17237
rect 12065 17232 13787 17234
rect 12065 17176 12070 17232
rect 12126 17176 13266 17232
rect 13322 17176 13726 17232
rect 13782 17176 13787 17232
rect 12065 17174 13787 17176
rect 12065 17171 12131 17174
rect 13261 17171 13327 17174
rect 13721 17171 13787 17174
rect 12249 17098 12315 17101
rect 14089 17098 14155 17101
rect 12249 17096 14155 17098
rect 12249 17040 12254 17096
rect 12310 17040 14094 17096
rect 14150 17040 14155 17096
rect 12249 17038 14155 17040
rect 12249 17035 12315 17038
rect 14089 17035 14155 17038
rect 25681 16962 25747 16965
rect 29600 16962 30000 16992
rect 25681 16960 30000 16962
rect 25681 16904 25686 16960
rect 25742 16904 30000 16960
rect 25681 16902 30000 16904
rect 25681 16899 25747 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 29600 16872 30000 16902
rect 25257 16831 25573 16832
rect 12750 16690 12756 16692
rect 12390 16630 12756 16690
rect 7097 16554 7163 16557
rect 12390 16554 12450 16630
rect 12750 16628 12756 16630
rect 12820 16628 12826 16692
rect 16849 16690 16915 16693
rect 16982 16690 16988 16692
rect 16849 16688 16988 16690
rect 16849 16632 16854 16688
rect 16910 16632 16988 16688
rect 16849 16630 16988 16632
rect 16849 16627 16915 16630
rect 16982 16628 16988 16630
rect 17052 16628 17058 16692
rect 23657 16690 23723 16693
rect 23790 16690 23796 16692
rect 23657 16688 23796 16690
rect 23657 16632 23662 16688
rect 23718 16632 23796 16688
rect 23657 16630 23796 16632
rect 23657 16627 23723 16630
rect 23790 16628 23796 16630
rect 23860 16628 23866 16692
rect 16665 16554 16731 16557
rect 7097 16552 16731 16554
rect 7097 16496 7102 16552
rect 7158 16496 16670 16552
rect 16726 16496 16731 16552
rect 7097 16494 16731 16496
rect 7097 16491 7163 16494
rect 16665 16491 16731 16494
rect 19425 16418 19491 16421
rect 20529 16418 20595 16421
rect 19425 16416 20595 16418
rect 19425 16360 19430 16416
rect 19486 16360 20534 16416
rect 20590 16360 20595 16416
rect 19425 16358 20595 16360
rect 19425 16355 19491 16358
rect 20529 16355 20595 16358
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 13813 16146 13879 16149
rect 17493 16146 17559 16149
rect 18505 16146 18571 16149
rect 13813 16144 18571 16146
rect 13813 16088 13818 16144
rect 13874 16088 17498 16144
rect 17554 16088 18510 16144
rect 18566 16088 18571 16144
rect 13813 16086 18571 16088
rect 13813 16083 13879 16086
rect 17493 16083 17559 16086
rect 18505 16083 18571 16086
rect 0 15874 400 15904
rect 749 15874 815 15877
rect 0 15872 815 15874
rect 0 15816 754 15872
rect 810 15816 815 15872
rect 0 15814 815 15816
rect 0 15784 400 15814
rect 749 15811 815 15814
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 14917 15602 14983 15605
rect 15929 15602 15995 15605
rect 14917 15600 15995 15602
rect 14917 15544 14922 15600
rect 14978 15544 15934 15600
rect 15990 15544 15995 15600
rect 14917 15542 15995 15544
rect 14917 15539 14983 15542
rect 15929 15539 15995 15542
rect 15561 15466 15627 15469
rect 16113 15466 16179 15469
rect 15561 15464 16179 15466
rect 15561 15408 15566 15464
rect 15622 15408 16118 15464
rect 16174 15408 16179 15464
rect 15561 15406 16179 15408
rect 15561 15403 15627 15406
rect 16113 15403 16179 15406
rect 20989 15466 21055 15469
rect 24761 15466 24827 15469
rect 20989 15464 24827 15466
rect 20989 15408 20994 15464
rect 21050 15408 24766 15464
rect 24822 15408 24827 15464
rect 20989 15406 24827 15408
rect 20989 15403 21055 15406
rect 24761 15403 24827 15406
rect 15469 15330 15535 15333
rect 15694 15330 15700 15332
rect 15469 15328 15700 15330
rect 15469 15272 15474 15328
rect 15530 15272 15700 15328
rect 15469 15270 15700 15272
rect 15469 15267 15535 15270
rect 15694 15268 15700 15270
rect 15764 15268 15770 15332
rect 23473 15330 23539 15333
rect 23606 15330 23612 15332
rect 23473 15328 23612 15330
rect 23473 15272 23478 15328
rect 23534 15272 23612 15328
rect 23473 15270 23612 15272
rect 23473 15267 23539 15270
rect 23606 15268 23612 15270
rect 23676 15268 23682 15332
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 4613 15194 4679 15197
rect 5022 15194 5028 15196
rect 4613 15192 5028 15194
rect 4613 15136 4618 15192
rect 4674 15136 5028 15192
rect 4613 15134 5028 15136
rect 4613 15131 4679 15134
rect 5022 15132 5028 15134
rect 5092 15194 5098 15196
rect 5349 15194 5415 15197
rect 5092 15192 5415 15194
rect 5092 15136 5354 15192
rect 5410 15136 5415 15192
rect 5092 15134 5415 15136
rect 5092 15132 5098 15134
rect 5349 15131 5415 15134
rect 12433 15194 12499 15197
rect 12566 15194 12572 15196
rect 12433 15192 12572 15194
rect 12433 15136 12438 15192
rect 12494 15136 12572 15192
rect 12433 15134 12572 15136
rect 12433 15131 12499 15134
rect 12566 15132 12572 15134
rect 12636 15132 12642 15196
rect 14590 15132 14596 15196
rect 14660 15132 14666 15196
rect 14598 15058 14658 15132
rect 19333 15058 19399 15061
rect 14598 15056 19399 15058
rect 14598 15000 19338 15056
rect 19394 15000 19399 15056
rect 14598 14998 19399 15000
rect 19333 14995 19399 14998
rect 10041 14922 10107 14925
rect 17125 14922 17191 14925
rect 21725 14922 21791 14925
rect 10041 14920 21791 14922
rect 10041 14864 10046 14920
rect 10102 14864 17130 14920
rect 17186 14864 21730 14920
rect 21786 14864 21791 14920
rect 10041 14862 21791 14864
rect 10041 14859 10107 14862
rect 17125 14859 17191 14862
rect 21725 14859 21791 14862
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 14733 14514 14799 14517
rect 16062 14514 16068 14516
rect 14733 14512 16068 14514
rect 14733 14456 14738 14512
rect 14794 14456 16068 14512
rect 14733 14454 16068 14456
rect 14733 14451 14799 14454
rect 16062 14452 16068 14454
rect 16132 14514 16138 14516
rect 16389 14514 16455 14517
rect 16132 14512 16455 14514
rect 16132 14456 16394 14512
rect 16450 14456 16455 14512
rect 16132 14454 16455 14456
rect 16132 14452 16138 14454
rect 16389 14451 16455 14454
rect 16389 14380 16455 14381
rect 16389 14378 16436 14380
rect 16344 14376 16436 14378
rect 16344 14320 16394 14376
rect 16344 14318 16436 14320
rect 16389 14316 16436 14318
rect 16500 14316 16506 14380
rect 16389 14315 16455 14316
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 0 13970 400 14000
rect 749 13970 815 13973
rect 0 13968 815 13970
rect 0 13912 754 13968
rect 810 13912 815 13968
rect 0 13910 815 13912
rect 0 13880 400 13910
rect 749 13907 815 13910
rect 5165 13698 5231 13701
rect 5574 13698 5580 13700
rect 5165 13696 5580 13698
rect 5165 13640 5170 13696
rect 5226 13640 5580 13696
rect 5165 13638 5580 13640
rect 5165 13635 5231 13638
rect 5574 13636 5580 13638
rect 5644 13636 5650 13700
rect 16573 13698 16639 13701
rect 17677 13698 17743 13701
rect 16573 13696 17743 13698
rect 16573 13640 16578 13696
rect 16634 13640 17682 13696
rect 17738 13640 17743 13696
rect 16573 13638 17743 13640
rect 16573 13635 16639 13638
rect 17677 13635 17743 13638
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 11605 13426 11671 13429
rect 14273 13426 14339 13429
rect 11605 13424 14339 13426
rect 11605 13368 11610 13424
rect 11666 13368 14278 13424
rect 14334 13368 14339 13424
rect 11605 13366 14339 13368
rect 11605 13363 11671 13366
rect 14273 13363 14339 13366
rect 17309 13426 17375 13429
rect 27613 13426 27679 13429
rect 17309 13424 27679 13426
rect 17309 13368 17314 13424
rect 17370 13368 27618 13424
rect 27674 13368 27679 13424
rect 17309 13366 27679 13368
rect 17309 13363 17375 13366
rect 27613 13363 27679 13366
rect 21357 13290 21423 13293
rect 22277 13290 22343 13293
rect 21357 13288 22343 13290
rect 21357 13232 21362 13288
rect 21418 13232 22282 13288
rect 22338 13232 22343 13288
rect 21357 13230 22343 13232
rect 21357 13227 21423 13230
rect 22277 13227 22343 13230
rect 17217 13156 17283 13157
rect 17166 13154 17172 13156
rect 17126 13094 17172 13154
rect 17236 13152 17283 13156
rect 17278 13096 17283 13152
rect 17166 13092 17172 13094
rect 17236 13092 17283 13096
rect 17217 13091 17283 13092
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 15837 12882 15903 12885
rect 19241 12882 19307 12885
rect 15837 12880 19307 12882
rect 15837 12824 15842 12880
rect 15898 12824 19246 12880
rect 19302 12824 19307 12880
rect 15837 12822 19307 12824
rect 15837 12819 15903 12822
rect 19241 12819 19307 12822
rect 20713 12882 20779 12885
rect 24393 12882 24459 12885
rect 20713 12880 24459 12882
rect 20713 12824 20718 12880
rect 20774 12824 24398 12880
rect 24454 12824 24459 12880
rect 20713 12822 24459 12824
rect 20713 12819 20779 12822
rect 24393 12819 24459 12822
rect 12801 12746 12867 12749
rect 22686 12746 22692 12748
rect 12801 12744 22692 12746
rect 12801 12688 12806 12744
rect 12862 12688 22692 12744
rect 12801 12686 22692 12688
rect 12801 12683 12867 12686
rect 22686 12684 22692 12686
rect 22756 12684 22762 12748
rect 16798 12548 16804 12612
rect 16868 12610 16874 12612
rect 16941 12610 17007 12613
rect 16868 12608 17007 12610
rect 16868 12552 16946 12608
rect 17002 12552 17007 12608
rect 16868 12550 17007 12552
rect 16868 12548 16874 12550
rect 16941 12547 17007 12550
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 12157 12338 12223 12341
rect 13670 12338 13676 12340
rect 12157 12336 13676 12338
rect 12157 12280 12162 12336
rect 12218 12280 13676 12336
rect 12157 12278 13676 12280
rect 12157 12275 12223 12278
rect 13670 12276 13676 12278
rect 13740 12276 13746 12340
rect 14365 12338 14431 12341
rect 19977 12340 20043 12341
rect 17534 12338 17540 12340
rect 14365 12336 17540 12338
rect 14365 12280 14370 12336
rect 14426 12280 17540 12336
rect 14365 12278 17540 12280
rect 14365 12275 14431 12278
rect 17534 12276 17540 12278
rect 17604 12276 17610 12340
rect 19926 12276 19932 12340
rect 19996 12338 20043 12340
rect 20897 12338 20963 12341
rect 21173 12338 21239 12341
rect 25773 12338 25839 12341
rect 29600 12338 30000 12368
rect 19996 12336 20088 12338
rect 20038 12280 20088 12336
rect 19996 12278 20088 12280
rect 20897 12336 21098 12338
rect 20897 12280 20902 12336
rect 20958 12280 21098 12336
rect 20897 12278 21098 12280
rect 19996 12276 20043 12278
rect 19977 12275 20043 12276
rect 20897 12275 20963 12278
rect 0 12066 400 12096
rect 749 12066 815 12069
rect 0 12064 815 12066
rect 0 12008 754 12064
rect 810 12008 815 12064
rect 0 12006 815 12008
rect 21038 12066 21098 12278
rect 21173 12336 21466 12338
rect 21173 12280 21178 12336
rect 21234 12280 21466 12336
rect 21173 12278 21466 12280
rect 21173 12275 21239 12278
rect 21173 12066 21239 12069
rect 21038 12064 21239 12066
rect 21038 12008 21178 12064
rect 21234 12008 21239 12064
rect 21038 12006 21239 12008
rect 0 11976 400 12006
rect 749 12003 815 12006
rect 21173 12003 21239 12006
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21406 11933 21466 12278
rect 25773 12336 30000 12338
rect 25773 12280 25778 12336
rect 25834 12280 30000 12336
rect 25773 12278 30000 12280
rect 25773 12275 25839 12278
rect 29600 12248 30000 12278
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 21406 11928 21515 11933
rect 21406 11872 21454 11928
rect 21510 11872 21515 11928
rect 21406 11870 21515 11872
rect 21449 11867 21515 11870
rect 20345 11794 20411 11797
rect 22001 11794 22067 11797
rect 20345 11792 22067 11794
rect 20345 11736 20350 11792
rect 20406 11736 22006 11792
rect 22062 11736 22067 11792
rect 20345 11734 22067 11736
rect 20345 11731 20411 11734
rect 22001 11731 22067 11734
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 9673 11386 9739 11389
rect 10685 11386 10751 11389
rect 9673 11384 10751 11386
rect 9673 11328 9678 11384
rect 9734 11328 10690 11384
rect 10746 11328 10751 11384
rect 9673 11326 10751 11328
rect 9673 11323 9739 11326
rect 10685 11323 10751 11326
rect 9765 11250 9831 11253
rect 14457 11250 14523 11253
rect 9765 11248 14523 11250
rect 9765 11192 9770 11248
rect 9826 11192 14462 11248
rect 14518 11192 14523 11248
rect 9765 11190 14523 11192
rect 9765 11187 9831 11190
rect 14457 11187 14523 11190
rect 15510 11052 15516 11116
rect 15580 11114 15586 11116
rect 15745 11114 15811 11117
rect 15580 11112 15811 11114
rect 15580 11056 15750 11112
rect 15806 11056 15811 11112
rect 15580 11054 15811 11056
rect 15580 11052 15586 11054
rect 15745 11051 15811 11054
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 19977 10706 20043 10709
rect 23289 10706 23355 10709
rect 19977 10704 23355 10706
rect 19977 10648 19982 10704
rect 20038 10648 23294 10704
rect 23350 10648 23355 10704
rect 19977 10646 23355 10648
rect 19977 10643 20043 10646
rect 23289 10643 23355 10646
rect 11053 10570 11119 10573
rect 18321 10570 18387 10573
rect 11053 10568 18387 10570
rect 11053 10512 11058 10568
rect 11114 10512 18326 10568
rect 18382 10512 18387 10568
rect 11053 10510 18387 10512
rect 11053 10507 11119 10510
rect 18321 10507 18387 10510
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 0 10162 400 10192
rect 749 10162 815 10165
rect 0 10160 815 10162
rect 0 10104 754 10160
rect 810 10104 815 10160
rect 0 10102 815 10104
rect 0 10072 400 10102
rect 749 10099 815 10102
rect 23013 10162 23079 10165
rect 27613 10162 27679 10165
rect 23013 10160 27679 10162
rect 23013 10104 23018 10160
rect 23074 10104 27618 10160
rect 27674 10104 27679 10160
rect 23013 10102 27679 10104
rect 23013 10099 23079 10102
rect 27613 10099 27679 10102
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 20437 9754 20503 9757
rect 20437 9752 20730 9754
rect 20437 9696 20442 9752
rect 20498 9696 20730 9752
rect 20437 9694 20730 9696
rect 20437 9691 20503 9694
rect 3550 9556 3556 9620
rect 3620 9618 3626 9620
rect 4153 9618 4219 9621
rect 3620 9616 4219 9618
rect 3620 9560 4158 9616
rect 4214 9560 4219 9616
rect 3620 9558 4219 9560
rect 3620 9556 3626 9558
rect 4153 9555 4219 9558
rect 10593 9618 10659 9621
rect 13445 9618 13511 9621
rect 10593 9616 13511 9618
rect 10593 9560 10598 9616
rect 10654 9560 13450 9616
rect 13506 9560 13511 9616
rect 10593 9558 13511 9560
rect 10593 9555 10659 9558
rect 13445 9555 13511 9558
rect 15285 9618 15351 9621
rect 17677 9618 17743 9621
rect 15285 9616 17743 9618
rect 15285 9560 15290 9616
rect 15346 9560 17682 9616
rect 17738 9560 17743 9616
rect 15285 9558 17743 9560
rect 20670 9618 20730 9694
rect 22001 9618 22067 9621
rect 23013 9620 23079 9621
rect 23013 9618 23060 9620
rect 20670 9616 22067 9618
rect 20670 9560 22006 9616
rect 22062 9560 22067 9616
rect 20670 9558 22067 9560
rect 22968 9616 23060 9618
rect 22968 9560 23018 9616
rect 22968 9558 23060 9560
rect 15285 9555 15351 9558
rect 17677 9555 17743 9558
rect 22001 9555 22067 9558
rect 23013 9556 23060 9558
rect 23124 9556 23130 9620
rect 23013 9555 23079 9556
rect 13353 9482 13419 9485
rect 20110 9482 20116 9484
rect 13353 9480 20116 9482
rect 13353 9424 13358 9480
rect 13414 9424 20116 9480
rect 13353 9422 20116 9424
rect 13353 9419 13419 9422
rect 20110 9420 20116 9422
rect 20180 9420 20186 9484
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 9857 9074 9923 9077
rect 10593 9074 10659 9077
rect 9857 9072 10659 9074
rect 9857 9016 9862 9072
rect 9918 9016 10598 9072
rect 10654 9016 10659 9072
rect 9857 9014 10659 9016
rect 9857 9011 9923 9014
rect 10593 9011 10659 9014
rect 12709 9074 12775 9077
rect 17033 9074 17099 9077
rect 12709 9072 17099 9074
rect 12709 9016 12714 9072
rect 12770 9016 17038 9072
rect 17094 9016 17099 9072
rect 12709 9014 17099 9016
rect 12709 9011 12775 9014
rect 17033 9011 17099 9014
rect 10685 8938 10751 8941
rect 13261 8938 13327 8941
rect 16113 8940 16179 8941
rect 10685 8936 13327 8938
rect 10685 8880 10690 8936
rect 10746 8880 13266 8936
rect 13322 8880 13327 8936
rect 10685 8878 13327 8880
rect 10685 8875 10751 8878
rect 13261 8875 13327 8878
rect 16062 8876 16068 8940
rect 16132 8938 16179 8940
rect 16132 8936 16224 8938
rect 16174 8880 16224 8936
rect 16132 8878 16224 8880
rect 16132 8876 16179 8878
rect 16113 8875 16179 8876
rect 16205 8802 16271 8805
rect 17769 8802 17835 8805
rect 16205 8800 17835 8802
rect 16205 8744 16210 8800
rect 16266 8744 17774 8800
rect 17830 8744 17835 8800
rect 16205 8742 17835 8744
rect 16205 8739 16271 8742
rect 17769 8739 17835 8742
rect 22645 8802 22711 8805
rect 23657 8802 23723 8805
rect 22645 8800 23723 8802
rect 22645 8744 22650 8800
rect 22706 8744 23662 8800
rect 23718 8744 23723 8800
rect 22645 8742 23723 8744
rect 22645 8739 22711 8742
rect 23657 8739 23723 8742
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 10961 8530 11027 8533
rect 15653 8530 15719 8533
rect 16021 8530 16087 8533
rect 10961 8528 16087 8530
rect 10961 8472 10966 8528
rect 11022 8472 15658 8528
rect 15714 8472 16026 8528
rect 16082 8472 16087 8528
rect 10961 8470 16087 8472
rect 10961 8467 11027 8470
rect 15653 8467 15719 8470
rect 16021 8467 16087 8470
rect 16481 8530 16547 8533
rect 22185 8530 22251 8533
rect 16481 8528 22251 8530
rect 16481 8472 16486 8528
rect 16542 8472 22190 8528
rect 22246 8472 22251 8528
rect 16481 8470 22251 8472
rect 16481 8467 16547 8470
rect 22185 8467 22251 8470
rect 21541 8394 21607 8397
rect 23841 8394 23907 8397
rect 21541 8392 23907 8394
rect 21541 8336 21546 8392
rect 21602 8336 23846 8392
rect 23902 8336 23907 8392
rect 21541 8334 23907 8336
rect 21541 8331 21607 8334
rect 23841 8331 23907 8334
rect 0 8258 400 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 400 8198
rect 1393 8195 1459 8198
rect 15694 8196 15700 8260
rect 15764 8258 15770 8260
rect 15837 8258 15903 8261
rect 15764 8256 15903 8258
rect 15764 8200 15842 8256
rect 15898 8200 15903 8256
rect 15764 8198 15903 8200
rect 15764 8196 15770 8198
rect 15837 8195 15903 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 20529 7986 20595 7989
rect 26601 7986 26667 7989
rect 20529 7984 26667 7986
rect 20529 7928 20534 7984
rect 20590 7928 26606 7984
rect 26662 7928 26667 7984
rect 20529 7926 26667 7928
rect 20529 7923 20595 7926
rect 26601 7923 26667 7926
rect 25865 7850 25931 7853
rect 25865 7848 29194 7850
rect 25865 7792 25870 7848
rect 25926 7792 29194 7848
rect 25865 7790 29194 7792
rect 25865 7787 25931 7790
rect 29134 7714 29194 7790
rect 29600 7714 30000 7744
rect 29134 7654 30000 7714
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 29600 7624 30000 7654
rect 28730 7583 29046 7584
rect 13445 7442 13511 7445
rect 14222 7442 14228 7444
rect 13445 7440 14228 7442
rect 13445 7384 13450 7440
rect 13506 7384 14228 7440
rect 13445 7382 14228 7384
rect 13445 7379 13511 7382
rect 14222 7380 14228 7382
rect 14292 7442 14298 7444
rect 17033 7442 17099 7445
rect 14292 7440 17099 7442
rect 14292 7384 17038 7440
rect 17094 7384 17099 7440
rect 14292 7382 17099 7384
rect 14292 7380 14298 7382
rect 17033 7379 17099 7382
rect 16389 7306 16455 7309
rect 16798 7306 16804 7308
rect 16389 7304 16804 7306
rect 16389 7248 16394 7304
rect 16450 7248 16804 7304
rect 16389 7246 16804 7248
rect 16389 7243 16455 7246
rect 16798 7244 16804 7246
rect 16868 7244 16874 7308
rect 22645 7306 22711 7309
rect 23606 7306 23612 7308
rect 22645 7304 23612 7306
rect 22645 7248 22650 7304
rect 22706 7248 23612 7304
rect 22645 7246 23612 7248
rect 22645 7243 22711 7246
rect 23606 7244 23612 7246
rect 23676 7244 23682 7308
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 16941 6900 17007 6901
rect 16941 6898 16988 6900
rect 16896 6896 16988 6898
rect 16896 6840 16946 6896
rect 16896 6838 16988 6840
rect 16941 6836 16988 6838
rect 17052 6836 17058 6900
rect 17166 6836 17172 6900
rect 17236 6898 17242 6900
rect 17953 6898 18019 6901
rect 17236 6896 18019 6898
rect 17236 6840 17958 6896
rect 18014 6840 18019 6896
rect 17236 6838 18019 6840
rect 17236 6836 17242 6838
rect 16941 6835 17007 6836
rect 17953 6835 18019 6838
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 0 6354 400 6384
rect 749 6354 815 6357
rect 0 6352 815 6354
rect 0 6296 754 6352
rect 810 6296 815 6352
rect 0 6294 815 6296
rect 0 6264 400 6294
rect 749 6291 815 6294
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 12525 5674 12591 5677
rect 12801 5674 12867 5677
rect 15285 5674 15351 5677
rect 17861 5674 17927 5677
rect 12525 5672 17927 5674
rect 12525 5616 12530 5672
rect 12586 5616 12806 5672
rect 12862 5616 15290 5672
rect 15346 5616 17866 5672
rect 17922 5616 17927 5672
rect 12525 5614 17927 5616
rect 12525 5611 12591 5614
rect 12801 5611 12867 5614
rect 15285 5611 15351 5614
rect 17861 5611 17927 5614
rect 22921 5538 22987 5541
rect 23790 5538 23796 5540
rect 22921 5536 23796 5538
rect 22921 5480 22926 5536
rect 22982 5480 23796 5536
rect 22921 5478 23796 5480
rect 22921 5475 22987 5478
rect 23790 5476 23796 5478
rect 23860 5476 23866 5540
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 13445 4722 13511 4725
rect 19149 4722 19215 4725
rect 13445 4720 19215 4722
rect 13445 4664 13450 4720
rect 13506 4664 19154 4720
rect 19210 4664 19215 4720
rect 13445 4662 19215 4664
rect 13445 4659 13511 4662
rect 19149 4659 19215 4662
rect 0 4450 400 4480
rect 749 4450 815 4453
rect 0 4448 815 4450
rect 0 4392 754 4448
rect 810 4392 815 4448
rect 0 4390 815 4392
rect 0 4360 400 4390
rect 749 4387 815 4390
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 25865 3090 25931 3093
rect 29600 3090 30000 3120
rect 25865 3088 30000 3090
rect 25865 3032 25870 3088
rect 25926 3032 30000 3088
rect 25865 3030 30000 3032
rect 25865 3027 25931 3030
rect 29600 3000 30000 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 0 2546 400 2576
rect 6494 2546 6500 2548
rect 0 2486 6500 2546
rect 0 2456 400 2486
rect 6494 2484 6500 2486
rect 6564 2484 6570 2548
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 4419 1664 4735 1665
rect 4419 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4735 1664
rect 4419 1599 4735 1600
rect 11365 1664 11681 1665
rect 11365 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11681 1664
rect 11365 1599 11681 1600
rect 18311 1664 18627 1665
rect 18311 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18627 1664
rect 18311 1599 18627 1600
rect 25257 1664 25573 1665
rect 25257 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25573 1664
rect 25257 1599 25573 1600
rect 7892 1120 8208 1121
rect 7892 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8208 1120
rect 7892 1055 8208 1056
rect 14838 1120 15154 1121
rect 14838 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15154 1120
rect 14838 1055 15154 1056
rect 21784 1120 22100 1121
rect 21784 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22100 1120
rect 21784 1055 22100 1056
rect 28730 1120 29046 1121
rect 28730 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29046 1120
rect 28730 1055 29046 1056
<< via3 >>
rect 7898 32668 7962 32672
rect 7898 32612 7902 32668
rect 7902 32612 7958 32668
rect 7958 32612 7962 32668
rect 7898 32608 7962 32612
rect 7978 32668 8042 32672
rect 7978 32612 7982 32668
rect 7982 32612 8038 32668
rect 8038 32612 8042 32668
rect 7978 32608 8042 32612
rect 8058 32668 8122 32672
rect 8058 32612 8062 32668
rect 8062 32612 8118 32668
rect 8118 32612 8122 32668
rect 8058 32608 8122 32612
rect 8138 32668 8202 32672
rect 8138 32612 8142 32668
rect 8142 32612 8198 32668
rect 8198 32612 8202 32668
rect 8138 32608 8202 32612
rect 14844 32668 14908 32672
rect 14844 32612 14848 32668
rect 14848 32612 14904 32668
rect 14904 32612 14908 32668
rect 14844 32608 14908 32612
rect 14924 32668 14988 32672
rect 14924 32612 14928 32668
rect 14928 32612 14984 32668
rect 14984 32612 14988 32668
rect 14924 32608 14988 32612
rect 15004 32668 15068 32672
rect 15004 32612 15008 32668
rect 15008 32612 15064 32668
rect 15064 32612 15068 32668
rect 15004 32608 15068 32612
rect 15084 32668 15148 32672
rect 15084 32612 15088 32668
rect 15088 32612 15144 32668
rect 15144 32612 15148 32668
rect 15084 32608 15148 32612
rect 21790 32668 21854 32672
rect 21790 32612 21794 32668
rect 21794 32612 21850 32668
rect 21850 32612 21854 32668
rect 21790 32608 21854 32612
rect 21870 32668 21934 32672
rect 21870 32612 21874 32668
rect 21874 32612 21930 32668
rect 21930 32612 21934 32668
rect 21870 32608 21934 32612
rect 21950 32668 22014 32672
rect 21950 32612 21954 32668
rect 21954 32612 22010 32668
rect 22010 32612 22014 32668
rect 21950 32608 22014 32612
rect 22030 32668 22094 32672
rect 22030 32612 22034 32668
rect 22034 32612 22090 32668
rect 22090 32612 22094 32668
rect 22030 32608 22094 32612
rect 28736 32668 28800 32672
rect 28736 32612 28740 32668
rect 28740 32612 28796 32668
rect 28796 32612 28800 32668
rect 28736 32608 28800 32612
rect 28816 32668 28880 32672
rect 28816 32612 28820 32668
rect 28820 32612 28876 32668
rect 28876 32612 28880 32668
rect 28816 32608 28880 32612
rect 28896 32668 28960 32672
rect 28896 32612 28900 32668
rect 28900 32612 28956 32668
rect 28956 32612 28960 32668
rect 28896 32608 28960 32612
rect 28976 32668 29040 32672
rect 28976 32612 28980 32668
rect 28980 32612 29036 32668
rect 29036 32612 29040 32668
rect 28976 32608 29040 32612
rect 4425 32124 4489 32128
rect 4425 32068 4429 32124
rect 4429 32068 4485 32124
rect 4485 32068 4489 32124
rect 4425 32064 4489 32068
rect 4505 32124 4569 32128
rect 4505 32068 4509 32124
rect 4509 32068 4565 32124
rect 4565 32068 4569 32124
rect 4505 32064 4569 32068
rect 4585 32124 4649 32128
rect 4585 32068 4589 32124
rect 4589 32068 4645 32124
rect 4645 32068 4649 32124
rect 4585 32064 4649 32068
rect 4665 32124 4729 32128
rect 4665 32068 4669 32124
rect 4669 32068 4725 32124
rect 4725 32068 4729 32124
rect 4665 32064 4729 32068
rect 11371 32124 11435 32128
rect 11371 32068 11375 32124
rect 11375 32068 11431 32124
rect 11431 32068 11435 32124
rect 11371 32064 11435 32068
rect 11451 32124 11515 32128
rect 11451 32068 11455 32124
rect 11455 32068 11511 32124
rect 11511 32068 11515 32124
rect 11451 32064 11515 32068
rect 11531 32124 11595 32128
rect 11531 32068 11535 32124
rect 11535 32068 11591 32124
rect 11591 32068 11595 32124
rect 11531 32064 11595 32068
rect 11611 32124 11675 32128
rect 11611 32068 11615 32124
rect 11615 32068 11671 32124
rect 11671 32068 11675 32124
rect 11611 32064 11675 32068
rect 18317 32124 18381 32128
rect 18317 32068 18321 32124
rect 18321 32068 18377 32124
rect 18377 32068 18381 32124
rect 18317 32064 18381 32068
rect 18397 32124 18461 32128
rect 18397 32068 18401 32124
rect 18401 32068 18457 32124
rect 18457 32068 18461 32124
rect 18397 32064 18461 32068
rect 18477 32124 18541 32128
rect 18477 32068 18481 32124
rect 18481 32068 18537 32124
rect 18537 32068 18541 32124
rect 18477 32064 18541 32068
rect 18557 32124 18621 32128
rect 18557 32068 18561 32124
rect 18561 32068 18617 32124
rect 18617 32068 18621 32124
rect 18557 32064 18621 32068
rect 25263 32124 25327 32128
rect 25263 32068 25267 32124
rect 25267 32068 25323 32124
rect 25323 32068 25327 32124
rect 25263 32064 25327 32068
rect 25343 32124 25407 32128
rect 25343 32068 25347 32124
rect 25347 32068 25403 32124
rect 25403 32068 25407 32124
rect 25343 32064 25407 32068
rect 25423 32124 25487 32128
rect 25423 32068 25427 32124
rect 25427 32068 25483 32124
rect 25483 32068 25487 32124
rect 25423 32064 25487 32068
rect 25503 32124 25567 32128
rect 25503 32068 25507 32124
rect 25507 32068 25563 32124
rect 25563 32068 25567 32124
rect 25503 32064 25567 32068
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 3740 27644 3804 27708
rect 16436 27508 16500 27572
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 5028 26964 5092 27028
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7236 26284 7300 26348
rect 21220 26284 21284 26348
rect 6684 26148 6748 26212
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 7420 26072 7484 26076
rect 7420 26016 7434 26072
rect 7434 26016 7484 26072
rect 7420 26012 7484 26016
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 3556 24984 3620 24988
rect 3556 24928 3570 24984
rect 3570 24928 3620 24984
rect 3556 24924 3620 24928
rect 4844 24652 4908 24716
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 6316 23760 6380 23764
rect 6316 23704 6366 23760
rect 6366 23704 6380 23760
rect 6316 23700 6380 23704
rect 12756 23624 12820 23628
rect 12756 23568 12806 23624
rect 12806 23568 12820 23624
rect 12756 23564 12820 23568
rect 3740 23488 3804 23492
rect 3740 23432 3754 23488
rect 3754 23432 3804 23488
rect 3740 23428 3804 23432
rect 7604 23428 7668 23492
rect 19932 23488 19996 23492
rect 19932 23432 19982 23488
rect 19982 23432 19996 23488
rect 19932 23428 19996 23432
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 16436 22944 16500 22948
rect 16436 22888 16450 22944
rect 16450 22888 16500 22944
rect 16436 22884 16500 22888
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 5396 22400 5460 22404
rect 5396 22344 5410 22400
rect 5410 22344 5460 22400
rect 5396 22340 5460 22344
rect 12572 22340 12636 22404
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 6316 21992 6380 21996
rect 6316 21936 6366 21992
rect 6366 21936 6380 21992
rect 6316 21932 6380 21936
rect 6684 21856 6748 21860
rect 6684 21800 6734 21856
rect 6734 21800 6748 21856
rect 6684 21796 6748 21800
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 7604 21720 7668 21724
rect 7604 21664 7654 21720
rect 7654 21664 7668 21720
rect 7604 21660 7668 21664
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4844 21448 4908 21452
rect 4844 21392 4894 21448
rect 4894 21392 4908 21448
rect 4844 21388 4908 21392
rect 7236 21388 7300 21452
rect 7420 21252 7484 21316
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 17540 21116 17604 21180
rect 6868 20708 6932 20772
rect 13676 20708 13740 20772
rect 14228 20708 14292 20772
rect 20116 20708 20180 20772
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 14596 19756 14660 19820
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 6500 19348 6564 19412
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 21220 18804 21284 18868
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 22692 18320 22756 18324
rect 22692 18264 22742 18320
rect 22742 18264 22756 18320
rect 22692 18260 22756 18264
rect 5580 18048 5644 18052
rect 5580 17992 5630 18048
rect 5630 17992 5644 18048
rect 5580 17988 5644 17992
rect 15516 17988 15580 18052
rect 23060 17988 23124 18052
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 4844 17852 4908 17916
rect 6868 17444 6932 17508
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 5396 17368 5460 17372
rect 5396 17312 5410 17368
rect 5410 17312 5460 17368
rect 5396 17308 5460 17312
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 12756 16628 12820 16692
rect 16988 16628 17052 16692
rect 23796 16628 23860 16692
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 15700 15268 15764 15332
rect 23612 15268 23676 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 5028 15132 5092 15196
rect 12572 15132 12636 15196
rect 14596 15132 14660 15196
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 16068 14452 16132 14516
rect 16436 14376 16500 14380
rect 16436 14320 16450 14376
rect 16450 14320 16500 14376
rect 16436 14316 16500 14320
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 5580 13636 5644 13700
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 17172 13152 17236 13156
rect 17172 13096 17222 13152
rect 17222 13096 17236 13152
rect 17172 13092 17236 13096
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 22692 12684 22756 12748
rect 16804 12548 16868 12612
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 13676 12276 13740 12340
rect 17540 12276 17604 12340
rect 19932 12336 19996 12340
rect 19932 12280 19982 12336
rect 19982 12280 19996 12336
rect 19932 12276 19996 12280
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 15516 11052 15580 11116
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 3556 9556 3620 9620
rect 23060 9616 23124 9620
rect 23060 9560 23074 9616
rect 23074 9560 23124 9616
rect 23060 9556 23124 9560
rect 20116 9420 20180 9484
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 16068 8936 16132 8940
rect 16068 8880 16118 8936
rect 16118 8880 16132 8936
rect 16068 8876 16132 8880
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 15700 8196 15764 8260
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 14228 7380 14292 7444
rect 16804 7244 16868 7308
rect 23612 7244 23676 7308
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 16988 6896 17052 6900
rect 16988 6840 17002 6896
rect 17002 6840 17052 6896
rect 16988 6836 17052 6840
rect 17172 6836 17236 6900
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 23796 5476 23860 5540
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 6500 2484 6564 2548
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
rect 4425 1660 4489 1664
rect 4425 1604 4429 1660
rect 4429 1604 4485 1660
rect 4485 1604 4489 1660
rect 4425 1600 4489 1604
rect 4505 1660 4569 1664
rect 4505 1604 4509 1660
rect 4509 1604 4565 1660
rect 4565 1604 4569 1660
rect 4505 1600 4569 1604
rect 4585 1660 4649 1664
rect 4585 1604 4589 1660
rect 4589 1604 4645 1660
rect 4645 1604 4649 1660
rect 4585 1600 4649 1604
rect 4665 1660 4729 1664
rect 4665 1604 4669 1660
rect 4669 1604 4725 1660
rect 4725 1604 4729 1660
rect 4665 1600 4729 1604
rect 11371 1660 11435 1664
rect 11371 1604 11375 1660
rect 11375 1604 11431 1660
rect 11431 1604 11435 1660
rect 11371 1600 11435 1604
rect 11451 1660 11515 1664
rect 11451 1604 11455 1660
rect 11455 1604 11511 1660
rect 11511 1604 11515 1660
rect 11451 1600 11515 1604
rect 11531 1660 11595 1664
rect 11531 1604 11535 1660
rect 11535 1604 11591 1660
rect 11591 1604 11595 1660
rect 11531 1600 11595 1604
rect 11611 1660 11675 1664
rect 11611 1604 11615 1660
rect 11615 1604 11671 1660
rect 11671 1604 11675 1660
rect 11611 1600 11675 1604
rect 18317 1660 18381 1664
rect 18317 1604 18321 1660
rect 18321 1604 18377 1660
rect 18377 1604 18381 1660
rect 18317 1600 18381 1604
rect 18397 1660 18461 1664
rect 18397 1604 18401 1660
rect 18401 1604 18457 1660
rect 18457 1604 18461 1660
rect 18397 1600 18461 1604
rect 18477 1660 18541 1664
rect 18477 1604 18481 1660
rect 18481 1604 18537 1660
rect 18537 1604 18541 1660
rect 18477 1600 18541 1604
rect 18557 1660 18621 1664
rect 18557 1604 18561 1660
rect 18561 1604 18617 1660
rect 18617 1604 18621 1660
rect 18557 1600 18621 1604
rect 25263 1660 25327 1664
rect 25263 1604 25267 1660
rect 25267 1604 25323 1660
rect 25323 1604 25327 1660
rect 25263 1600 25327 1604
rect 25343 1660 25407 1664
rect 25343 1604 25347 1660
rect 25347 1604 25403 1660
rect 25403 1604 25407 1660
rect 25343 1600 25407 1604
rect 25423 1660 25487 1664
rect 25423 1604 25427 1660
rect 25427 1604 25483 1660
rect 25483 1604 25487 1660
rect 25423 1600 25487 1604
rect 25503 1660 25567 1664
rect 25503 1604 25507 1660
rect 25507 1604 25563 1660
rect 25563 1604 25567 1660
rect 25503 1600 25567 1604
rect 7898 1116 7962 1120
rect 7898 1060 7902 1116
rect 7902 1060 7958 1116
rect 7958 1060 7962 1116
rect 7898 1056 7962 1060
rect 7978 1116 8042 1120
rect 7978 1060 7982 1116
rect 7982 1060 8038 1116
rect 8038 1060 8042 1116
rect 7978 1056 8042 1060
rect 8058 1116 8122 1120
rect 8058 1060 8062 1116
rect 8062 1060 8118 1116
rect 8118 1060 8122 1116
rect 8058 1056 8122 1060
rect 8138 1116 8202 1120
rect 8138 1060 8142 1116
rect 8142 1060 8198 1116
rect 8198 1060 8202 1116
rect 8138 1056 8202 1060
rect 14844 1116 14908 1120
rect 14844 1060 14848 1116
rect 14848 1060 14904 1116
rect 14904 1060 14908 1116
rect 14844 1056 14908 1060
rect 14924 1116 14988 1120
rect 14924 1060 14928 1116
rect 14928 1060 14984 1116
rect 14984 1060 14988 1116
rect 14924 1056 14988 1060
rect 15004 1116 15068 1120
rect 15004 1060 15008 1116
rect 15008 1060 15064 1116
rect 15064 1060 15068 1116
rect 15004 1056 15068 1060
rect 15084 1116 15148 1120
rect 15084 1060 15088 1116
rect 15088 1060 15144 1116
rect 15144 1060 15148 1116
rect 15084 1056 15148 1060
rect 21790 1116 21854 1120
rect 21790 1060 21794 1116
rect 21794 1060 21850 1116
rect 21850 1060 21854 1116
rect 21790 1056 21854 1060
rect 21870 1116 21934 1120
rect 21870 1060 21874 1116
rect 21874 1060 21930 1116
rect 21930 1060 21934 1116
rect 21870 1056 21934 1060
rect 21950 1116 22014 1120
rect 21950 1060 21954 1116
rect 21954 1060 22010 1116
rect 22010 1060 22014 1116
rect 21950 1056 22014 1060
rect 22030 1116 22094 1120
rect 22030 1060 22034 1116
rect 22034 1060 22090 1116
rect 22090 1060 22094 1116
rect 22030 1056 22094 1060
rect 28736 1116 28800 1120
rect 28736 1060 28740 1116
rect 28740 1060 28796 1116
rect 28796 1060 28800 1116
rect 28736 1056 28800 1060
rect 28816 1116 28880 1120
rect 28816 1060 28820 1116
rect 28820 1060 28876 1116
rect 28876 1060 28880 1116
rect 28816 1056 28880 1060
rect 28896 1116 28960 1120
rect 28896 1060 28900 1116
rect 28900 1060 28956 1116
rect 28956 1060 28960 1116
rect 28896 1056 28960 1060
rect 28976 1116 29040 1120
rect 28976 1060 28980 1116
rect 28980 1060 29036 1116
rect 29036 1060 29040 1116
rect 28976 1056 29040 1060
<< metal4 >>
rect 4417 32128 4737 32688
rect 4417 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4737 32128
rect 4417 31040 4737 32064
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 3739 27708 3805 27709
rect 3739 27644 3740 27708
rect 3804 27644 3805 27708
rect 3739 27643 3805 27644
rect 3555 24988 3621 24989
rect 3555 24924 3556 24988
rect 3620 24924 3621 24988
rect 3555 24923 3621 24924
rect 3558 9621 3618 24923
rect 3742 23493 3802 27643
rect 4417 26688 4737 27712
rect 7890 32672 8210 32688
rect 7890 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8210 32672
rect 7890 31584 8210 32608
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 5027 27028 5093 27029
rect 5027 26964 5028 27028
rect 5092 26964 5093 27028
rect 5027 26963 5093 26964
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4843 24716 4909 24717
rect 4843 24652 4844 24716
rect 4908 24652 4909 24716
rect 4843 24651 4909 24652
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 3739 23492 3805 23493
rect 3739 23428 3740 23492
rect 3804 23428 3805 23492
rect 3739 23427 3805 23428
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4846 21453 4906 24651
rect 4843 21452 4909 21453
rect 4843 21388 4844 21452
rect 4908 21388 4909 21452
rect 4843 21387 4909 21388
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4846 17917 4906 21387
rect 4843 17916 4909 17917
rect 4843 17852 4844 17916
rect 4908 17852 4909 17916
rect 4843 17851 4909 17852
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 5030 15197 5090 26963
rect 7235 26348 7301 26349
rect 7235 26284 7236 26348
rect 7300 26284 7301 26348
rect 7235 26283 7301 26284
rect 6683 26212 6749 26213
rect 6683 26148 6684 26212
rect 6748 26148 6749 26212
rect 6683 26147 6749 26148
rect 6315 23764 6381 23765
rect 6315 23700 6316 23764
rect 6380 23700 6381 23764
rect 6315 23699 6381 23700
rect 5395 22404 5461 22405
rect 5395 22340 5396 22404
rect 5460 22340 5461 22404
rect 5395 22339 5461 22340
rect 5398 17373 5458 22339
rect 6318 21997 6378 23699
rect 6315 21996 6381 21997
rect 6315 21932 6316 21996
rect 6380 21932 6381 21996
rect 6315 21931 6381 21932
rect 6686 21861 6746 26147
rect 6683 21860 6749 21861
rect 6683 21796 6684 21860
rect 6748 21796 6749 21860
rect 6683 21795 6749 21796
rect 7238 21453 7298 26283
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7419 26076 7485 26077
rect 7419 26012 7420 26076
rect 7484 26012 7485 26076
rect 7419 26011 7485 26012
rect 7235 21452 7301 21453
rect 7235 21388 7236 21452
rect 7300 21388 7301 21452
rect 7235 21387 7301 21388
rect 7422 21317 7482 26011
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7603 23492 7669 23493
rect 7603 23428 7604 23492
rect 7668 23428 7669 23492
rect 7603 23427 7669 23428
rect 7606 21725 7666 23427
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7603 21724 7669 21725
rect 7603 21660 7604 21724
rect 7668 21660 7669 21724
rect 7603 21659 7669 21660
rect 7419 21316 7485 21317
rect 7419 21252 7420 21316
rect 7484 21252 7485 21316
rect 7419 21251 7485 21252
rect 6867 20772 6933 20773
rect 6867 20708 6868 20772
rect 6932 20708 6933 20772
rect 6867 20707 6933 20708
rect 6499 19412 6565 19413
rect 6499 19348 6500 19412
rect 6564 19348 6565 19412
rect 6499 19347 6565 19348
rect 5579 18052 5645 18053
rect 5579 17988 5580 18052
rect 5644 17988 5645 18052
rect 5579 17987 5645 17988
rect 5395 17372 5461 17373
rect 5395 17308 5396 17372
rect 5460 17308 5461 17372
rect 5395 17307 5461 17308
rect 5027 15196 5093 15197
rect 5027 15132 5028 15196
rect 5092 15132 5093 15196
rect 5027 15131 5093 15132
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 5582 13701 5642 17987
rect 5579 13700 5645 13701
rect 5579 13636 5580 13700
rect 5644 13636 5645 13700
rect 5579 13635 5645 13636
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 3555 9620 3621 9621
rect 3555 9556 3556 9620
rect 3620 9556 3621 9620
rect 3555 9555 3621 9556
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 1664 4737 2688
rect 6502 2549 6562 19347
rect 6870 17509 6930 20707
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 6867 17508 6933 17509
rect 6867 17444 6868 17508
rect 6932 17444 6933 17508
rect 6867 17443 6933 17444
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 6499 2548 6565 2549
rect 6499 2484 6500 2548
rect 6564 2484 6565 2548
rect 6499 2483 6565 2484
rect 4417 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4737 1664
rect 4417 1040 4737 1600
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 1120 8210 2144
rect 7890 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8210 1120
rect 7890 1040 8210 1056
rect 11363 32128 11683 32688
rect 11363 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11683 32128
rect 11363 31040 11683 32064
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 14836 32672 15156 32688
rect 14836 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15156 32672
rect 14836 31584 15156 32608
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 18309 32128 18629 32688
rect 18309 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18629 32128
rect 18309 31040 18629 32064
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 16435 27572 16501 27573
rect 16435 27508 16436 27572
rect 16500 27508 16501 27572
rect 16435 27507 16501 27508
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 12755 23628 12821 23629
rect 12755 23564 12756 23628
rect 12820 23564 12821 23628
rect 12755 23563 12821 23564
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 12571 22404 12637 22405
rect 12571 22340 12572 22404
rect 12636 22340 12637 22404
rect 12571 22339 12637 22340
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 12574 15197 12634 22339
rect 12758 16693 12818 23563
rect 14836 22880 15156 23904
rect 16438 22949 16498 27507
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 21782 32672 22102 32688
rect 21782 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22102 32672
rect 21782 31584 22102 32608
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21219 26348 21285 26349
rect 21219 26284 21220 26348
rect 21284 26284 21285 26348
rect 21219 26283 21285 26284
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 19931 23492 19997 23493
rect 19931 23428 19932 23492
rect 19996 23428 19997 23492
rect 19931 23427 19997 23428
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 16435 22948 16501 22949
rect 16435 22884 16436 22948
rect 16500 22884 16501 22948
rect 16435 22883 16501 22884
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 13675 20772 13741 20773
rect 13675 20708 13676 20772
rect 13740 20708 13741 20772
rect 13675 20707 13741 20708
rect 14227 20772 14293 20773
rect 14227 20708 14228 20772
rect 14292 20708 14293 20772
rect 14227 20707 14293 20708
rect 12755 16692 12821 16693
rect 12755 16628 12756 16692
rect 12820 16628 12821 16692
rect 12755 16627 12821 16628
rect 12571 15196 12637 15197
rect 12571 15132 12572 15196
rect 12636 15132 12637 15196
rect 12571 15131 12637 15132
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 13678 12341 13738 20707
rect 13675 12340 13741 12341
rect 13675 12276 13676 12340
rect 13740 12276 13741 12340
rect 13675 12275 13741 12276
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 14230 7445 14290 20707
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14595 19820 14661 19821
rect 14595 19756 14596 19820
rect 14660 19756 14661 19820
rect 14595 19755 14661 19756
rect 14598 15197 14658 19755
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14595 15196 14661 15197
rect 14595 15132 14596 15196
rect 14660 15132 14661 15196
rect 14595 15131 14661 15132
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 15518 11117 15578 17987
rect 15699 15332 15765 15333
rect 15699 15268 15700 15332
rect 15764 15268 15765 15332
rect 15699 15267 15765 15268
rect 15515 11116 15581 11117
rect 15515 11052 15516 11116
rect 15580 11052 15581 11116
rect 15515 11051 15581 11052
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 15702 8261 15762 15267
rect 16067 14516 16133 14517
rect 16067 14452 16068 14516
rect 16132 14452 16133 14516
rect 16067 14451 16133 14452
rect 16070 8941 16130 14451
rect 16438 14381 16498 22883
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 17539 21180 17605 21181
rect 17539 21116 17540 21180
rect 17604 21116 17605 21180
rect 17539 21115 17605 21116
rect 16987 16692 17053 16693
rect 16987 16628 16988 16692
rect 17052 16628 17053 16692
rect 16987 16627 17053 16628
rect 16435 14380 16501 14381
rect 16435 14316 16436 14380
rect 16500 14316 16501 14380
rect 16435 14315 16501 14316
rect 16803 12612 16869 12613
rect 16803 12548 16804 12612
rect 16868 12548 16869 12612
rect 16803 12547 16869 12548
rect 16067 8940 16133 8941
rect 16067 8876 16068 8940
rect 16132 8876 16133 8940
rect 16067 8875 16133 8876
rect 15699 8260 15765 8261
rect 15699 8196 15700 8260
rect 15764 8196 15765 8260
rect 15699 8195 15765 8196
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14227 7444 14293 7445
rect 14227 7380 14228 7444
rect 14292 7380 14293 7444
rect 14227 7379 14293 7380
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 1664 11683 2688
rect 11363 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11683 1664
rect 11363 1040 11683 1600
rect 14836 6560 15156 7584
rect 16806 7309 16866 12547
rect 16803 7308 16869 7309
rect 16803 7244 16804 7308
rect 16868 7244 16869 7308
rect 16803 7243 16869 7244
rect 16990 6901 17050 16627
rect 17171 13156 17237 13157
rect 17171 13092 17172 13156
rect 17236 13092 17237 13156
rect 17171 13091 17237 13092
rect 17174 6901 17234 13091
rect 17542 12341 17602 21115
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 17539 12340 17605 12341
rect 17539 12276 17540 12340
rect 17604 12276 17605 12340
rect 17539 12275 17605 12276
rect 18309 11456 18629 12480
rect 19934 12341 19994 23427
rect 20115 20772 20181 20773
rect 20115 20708 20116 20772
rect 20180 20708 20181 20772
rect 20115 20707 20181 20708
rect 19931 12340 19997 12341
rect 19931 12276 19932 12340
rect 19996 12276 19997 12340
rect 19931 12275 19997 12276
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 20118 9485 20178 20707
rect 21222 18869 21282 26283
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21219 18868 21285 18869
rect 21219 18804 21220 18868
rect 21284 18804 21285 18868
rect 21219 18803 21285 18804
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 25255 32128 25575 32688
rect 25255 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25575 32128
rect 25255 31040 25575 32064
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 22691 18324 22757 18325
rect 22691 18260 22692 18324
rect 22756 18260 22757 18324
rect 22691 18259 22757 18260
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 22694 12749 22754 18259
rect 23059 18052 23125 18053
rect 23059 17988 23060 18052
rect 23124 17988 23125 18052
rect 23059 17987 23125 17988
rect 22691 12748 22757 12749
rect 22691 12684 22692 12748
rect 22756 12684 22757 12748
rect 22691 12683 22757 12684
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 20115 9484 20181 9485
rect 20115 9420 20116 9484
rect 20180 9420 20181 9484
rect 20115 9419 20181 9420
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 16987 6900 17053 6901
rect 16987 6836 16988 6900
rect 17052 6836 17053 6900
rect 16987 6835 17053 6836
rect 17171 6900 17237 6901
rect 17171 6836 17172 6900
rect 17236 6836 17237 6900
rect 17171 6835 17237 6836
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 1120 15156 2144
rect 14836 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15156 1120
rect 14836 1040 15156 1056
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 1664 18629 2688
rect 18309 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18629 1664
rect 18309 1040 18629 1600
rect 21782 8736 22102 9760
rect 23062 9621 23122 17987
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 23795 16692 23861 16693
rect 23795 16628 23796 16692
rect 23860 16628 23861 16692
rect 23795 16627 23861 16628
rect 23611 15332 23677 15333
rect 23611 15268 23612 15332
rect 23676 15268 23677 15332
rect 23611 15267 23677 15268
rect 23059 9620 23125 9621
rect 23059 9556 23060 9620
rect 23124 9556 23125 9620
rect 23059 9555 23125 9556
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 23614 7309 23674 15267
rect 23611 7308 23677 7309
rect 23611 7244 23612 7308
rect 23676 7244 23677 7308
rect 23611 7243 23677 7244
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 23798 5541 23858 16627
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 23795 5540 23861 5541
rect 23795 5476 23796 5540
rect 23860 5476 23861 5540
rect 23795 5475 23861 5476
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 1120 22102 2144
rect 21782 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22102 1120
rect 21782 1040 22102 1056
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 1664 25575 2688
rect 25255 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25575 1664
rect 25255 1040 25575 1600
rect 28728 32672 29048 32688
rect 28728 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29048 32672
rect 28728 31584 29048 32608
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 1120 29048 2144
rect 28728 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29048 1120
rect 28728 1040 29048 1056
use sky130_fd_sc_hd__or4_1  _0902_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8096 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _0903_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0904_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2116 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0905_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0906_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0907_
timestamp 1694700623
transform 1 0 2392 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0908_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1840 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0909_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0910_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0911_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3312 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0912_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2300 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0913_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2668 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0914_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0915_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0916_
timestamp 1694700623
transform 1 0 3128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0917_
timestamp 1694700623
transform -1 0 2208 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0918_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0919_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3496 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0920_
timestamp 1694700623
transform -1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0921_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0922_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4416 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_4  _0924_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_1  _0925_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0926_
timestamp 1694700623
transform 1 0 1564 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1694700623
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0928_
timestamp 1694700623
transform -1 0 8832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _0929_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3680 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0930_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0931_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1656 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0932_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0933_
timestamp 1694700623
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1694700623
transform -1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1694700623
transform -1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0936_
timestamp 1694700623
transform -1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0937_
timestamp 1694700623
transform -1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _0938_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 20608 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1694700623
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0940_
timestamp 1694700623
transform -1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0941_
timestamp 1694700623
transform 1 0 12788 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0942_
timestamp 1694700623
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _0943_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1694700623
transform 1 0 17848 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1694700623
transform -1 0 17940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0946_
timestamp 1694700623
transform 1 0 22816 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _0947_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20516 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1694700623
transform 1 0 17480 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1694700623
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_1  _0950_
timestamp 1694700623
transform -1 0 13524 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0951_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19044 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0952_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22540 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0953_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1694700623
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0955_
timestamp 1694700623
transform 1 0 20424 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0956_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19596 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0957_
timestamp 1694700623
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1694700623
transform -1 0 23276 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0959_
timestamp 1694700623
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _0960_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21528 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1694700623
transform 1 0 17940 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0962_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 16284 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1694700623
transform -1 0 18400 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1694700623
transform 1 0 19228 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0965_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 23644 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0966_
timestamp 1694700623
transform -1 0 24012 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _0967_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1694700623
transform 1 0 22816 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0969_
timestamp 1694700623
transform -1 0 13984 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _0970_
timestamp 1694700623
transform 1 0 18308 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0971_
timestamp 1694700623
transform 1 0 23736 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _0972_
timestamp 1694700623
transform -1 0 14444 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1694700623
transform 1 0 22816 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0974_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22908 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0975_
timestamp 1694700623
transform -1 0 23736 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _0976_
timestamp 1694700623
transform -1 0 13248 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _0977_
timestamp 1694700623
transform -1 0 16560 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0978_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0979_
timestamp 1694700623
transform -1 0 16100 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _0980_
timestamp 1694700623
transform 1 0 13248 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0981_
timestamp 1694700623
transform -1 0 19136 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0982_
timestamp 1694700623
transform 1 0 16008 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0983_
timestamp 1694700623
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0984_
timestamp 1694700623
transform 1 0 15364 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0985_
timestamp 1694700623
transform -1 0 22448 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0986_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14628 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0987_
timestamp 1694700623
transform -1 0 16376 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0988_
timestamp 1694700623
transform -1 0 14536 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0989_
timestamp 1694700623
transform -1 0 10672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _0990_
timestamp 1694700623
transform -1 0 14628 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1694700623
transform -1 0 11224 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0992_
timestamp 1694700623
transform -1 0 9752 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0993_
timestamp 1694700623
transform -1 0 17204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0994_
timestamp 1694700623
transform -1 0 10304 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1694700623
transform 1 0 16744 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0996_
timestamp 1694700623
transform -1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0997_
timestamp 1694700623
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0998_
timestamp 1694700623
transform 1 0 9292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0999_
timestamp 1694700623
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1000_
timestamp 1694700623
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1694700623
transform 1 0 20884 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1002_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1003_
timestamp 1694700623
transform -1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1004_
timestamp 1694700623
transform 1 0 23092 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1694700623
transform 1 0 22816 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1006_
timestamp 1694700623
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1007_
timestamp 1694700623
transform -1 0 24288 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 1694700623
transform 1 0 9752 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1694700623
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1010_
timestamp 1694700623
transform -1 0 15272 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1011_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9844 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 1694700623
transform 1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1694700623
transform -1 0 15548 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1014_
timestamp 1694700623
transform -1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1015_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1016_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9108 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 1694700623
transform 1 0 19780 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1018_
timestamp 1694700623
transform 1 0 19596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 1694700623
transform 1 0 19044 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1020_
timestamp 1694700623
transform 1 0 19596 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1694700623
transform -1 0 21160 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1694700623
transform -1 0 21160 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1023_
timestamp 1694700623
transform 1 0 20240 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1024_
timestamp 1694700623
transform 1 0 20332 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1694700623
transform 1 0 15272 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1694700623
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1027_
timestamp 1694700623
transform 1 0 19780 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1028_
timestamp 1694700623
transform -1 0 22356 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1029_
timestamp 1694700623
transform 1 0 19780 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1030_
timestamp 1694700623
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1694700623
transform 1 0 20332 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1032_
timestamp 1694700623
transform -1 0 23368 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1033_
timestamp 1694700623
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _1034_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 20148 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1035_
timestamp 1694700623
transform -1 0 20792 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1036_
timestamp 1694700623
transform -1 0 18768 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 1694700623
transform 1 0 14996 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1038_
timestamp 1694700623
transform 1 0 15640 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1039_
timestamp 1694700623
transform 1 0 15916 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1040_
timestamp 1694700623
transform 1 0 15824 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1041_
timestamp 1694700623
transform 1 0 15824 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1042_
timestamp 1694700623
transform 1 0 15456 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1043_
timestamp 1694700623
transform -1 0 16376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1694700623
transform -1 0 16008 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1045_
timestamp 1694700623
transform 1 0 15456 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 1694700623
transform -1 0 22264 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1047_
timestamp 1694700623
transform 1 0 16928 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1048_
timestamp 1694700623
transform -1 0 18124 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1049_
timestamp 1694700623
transform 1 0 17296 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _1050_
timestamp 1694700623
transform 1 0 15180 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1051_
timestamp 1694700623
transform -1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1052_
timestamp 1694700623
transform -1 0 13064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1053_
timestamp 1694700623
transform 1 0 18952 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1054_
timestamp 1694700623
transform 1 0 18216 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1055_
timestamp 1694700623
transform 1 0 18584 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1056_
timestamp 1694700623
transform -1 0 20056 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1694700623
transform -1 0 15548 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1058_
timestamp 1694700623
transform -1 0 14996 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1059_
timestamp 1694700623
transform 1 0 14260 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1060_
timestamp 1694700623
transform 1 0 14260 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1061_
timestamp 1694700623
transform -1 0 16100 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1062_
timestamp 1694700623
transform -1 0 14536 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1063_
timestamp 1694700623
transform 1 0 12512 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1064_
timestamp 1694700623
transform 1 0 13156 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1694700623
transform -1 0 13524 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1066_
timestamp 1694700623
transform 1 0 12512 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1067_
timestamp 1694700623
transform 1 0 12052 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1068_
timestamp 1694700623
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1694700623
transform 1 0 13064 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1694700623
transform -1 0 14720 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1071_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13432 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1072_
timestamp 1694700623
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1073_
timestamp 1694700623
transform -1 0 17572 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 1694700623
transform -1 0 18860 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1075_
timestamp 1694700623
transform -1 0 17940 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1076_
timestamp 1694700623
transform 1 0 15640 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1077_
timestamp 1694700623
transform 1 0 17112 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1078_
timestamp 1694700623
transform -1 0 20884 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1694700623
transform 1 0 20148 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1080_
timestamp 1694700623
transform -1 0 21160 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1081_
timestamp 1694700623
transform 1 0 20056 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1082_
timestamp 1694700623
transform -1 0 17572 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1694700623
transform 1 0 10764 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1084_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1694700623
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1694700623
transform -1 0 10672 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1694700623
transform 1 0 9292 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1088_
timestamp 1694700623
transform 1 0 16744 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1089_
timestamp 1694700623
transform 1 0 17480 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1090_
timestamp 1694700623
transform 1 0 17204 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1091_
timestamp 1694700623
transform 1 0 17480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 1694700623
transform 1 0 15916 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1093_
timestamp 1694700623
transform -1 0 18400 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1094_
timestamp 1694700623
transform 1 0 16008 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1095_
timestamp 1694700623
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1096_
timestamp 1694700623
transform -1 0 17572 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1097_
timestamp 1694700623
transform 1 0 16100 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1098_
timestamp 1694700623
transform 1 0 16008 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1099_
timestamp 1694700623
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1100_
timestamp 1694700623
transform -1 0 18860 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 1694700623
transform -1 0 19688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1102_
timestamp 1694700623
transform -1 0 18492 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1103_
timestamp 1694700623
transform 1 0 17756 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1104_
timestamp 1694700623
transform -1 0 16928 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1105_
timestamp 1694700623
transform -1 0 19688 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1106_
timestamp 1694700623
transform 1 0 16008 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1107_
timestamp 1694700623
transform -1 0 20424 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1108_
timestamp 1694700623
transform -1 0 17204 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1109_
timestamp 1694700623
transform -1 0 17480 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1110_
timestamp 1694700623
transform -1 0 18860 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1694700623
transform 1 0 16100 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1112_
timestamp 1694700623
transform -1 0 17020 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1113_
timestamp 1694700623
transform 1 0 18584 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 1694700623
transform -1 0 19688 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1115_
timestamp 1694700623
transform -1 0 19136 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1116_
timestamp 1694700623
transform 1 0 18584 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1117_
timestamp 1694700623
transform 1 0 16744 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1118_
timestamp 1694700623
transform -1 0 19044 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1119_
timestamp 1694700623
transform 1 0 17020 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1120_
timestamp 1694700623
transform -1 0 16928 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1121_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11868 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1122_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1123_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11776 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1124_
timestamp 1694700623
transform 1 0 11224 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1125_
timestamp 1694700623
transform -1 0 10488 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _1126_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 11132 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1127_
timestamp 1694700623
transform 1 0 22264 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1128_
timestamp 1694700623
transform 1 0 21804 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1129_
timestamp 1694700623
transform -1 0 22632 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1130_
timestamp 1694700623
transform 1 0 22080 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1694700623
transform -1 0 23276 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 1694700623
transform 1 0 21896 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1133_
timestamp 1694700623
transform -1 0 23736 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1134_
timestamp 1694700623
transform 1 0 22356 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1694700623
transform -1 0 23736 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1136_
timestamp 1694700623
transform 1 0 22632 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1137_
timestamp 1694700623
transform -1 0 24288 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1138_
timestamp 1694700623
transform 1 0 22540 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1139_
timestamp 1694700623
transform 1 0 14996 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1140_
timestamp 1694700623
transform -1 0 15916 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1141_
timestamp 1694700623
transform 1 0 14260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1142_
timestamp 1694700623
transform -1 0 16008 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1143_
timestamp 1694700623
transform 1 0 22356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 1694700623
transform 1 0 10672 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1145_
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1146_
timestamp 1694700623
transform 1 0 10672 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1147_
timestamp 1694700623
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1148_
timestamp 1694700623
transform 1 0 10580 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1149_
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1150_
timestamp 1694700623
transform -1 0 12788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 1694700623
transform -1 0 24196 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1152_
timestamp 1694700623
transform 1 0 20976 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1694700623
transform 1 0 23368 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1154_
timestamp 1694700623
transform 1 0 23276 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1155_
timestamp 1694700623
transform -1 0 12788 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1156_
timestamp 1694700623
transform -1 0 12512 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1157_
timestamp 1694700623
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1158_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 11500 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1159_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 10948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1160_
timestamp 1694700623
transform 1 0 12052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1161_
timestamp 1694700623
transform -1 0 11040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1162_
timestamp 1694700623
transform 1 0 10304 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1163_
timestamp 1694700623
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1164_
timestamp 1694700623
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _1165_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9844 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1166_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1694700623
transform 1 0 10304 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1168_
timestamp 1694700623
transform 1 0 11132 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1694700623
transform 1 0 11500 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1170_
timestamp 1694700623
transform 1 0 10764 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1694700623
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1172_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9568 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1173_
timestamp 1694700623
transform 1 0 10304 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1174_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10948 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__o22ai_2  _1175_
timestamp 1694700623
transform -1 0 9844 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 1694700623
transform 1 0 10304 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1177_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1178_
timestamp 1694700623
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1179_
timestamp 1694700623
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1180_
timestamp 1694700623
transform -1 0 23092 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1181_
timestamp 1694700623
transform 1 0 22264 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1694700623
transform -1 0 22908 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1183_
timestamp 1694700623
transform -1 0 22448 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1694700623
transform -1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1185_
timestamp 1694700623
transform 1 0 14720 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1186_
timestamp 1694700623
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1694700623
transform -1 0 22356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1188_
timestamp 1694700623
transform 1 0 9384 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1189_
timestamp 1694700623
transform 1 0 9936 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1190_
timestamp 1694700623
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1191_
timestamp 1694700623
transform -1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1192_
timestamp 1694700623
transform -1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1193_
timestamp 1694700623
transform 1 0 8924 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1194_
timestamp 1694700623
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1195_
timestamp 1694700623
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1694700623
transform 1 0 9016 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1694700623
transform -1 0 11224 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1198_
timestamp 1694700623
transform -1 0 10212 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1694700623
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1694700623
transform -1 0 9200 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1201_
timestamp 1694700623
transform 1 0 10580 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1694700623
transform -1 0 12604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1203_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10672 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1204_
timestamp 1694700623
transform -1 0 12512 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1205_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1694700623
transform 1 0 10856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _1207_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1694700623
transform -1 0 10672 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1209_
timestamp 1694700623
transform -1 0 11960 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1694700623
transform 1 0 9108 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1211_
timestamp 1694700623
transform -1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1694700623
transform -1 0 11316 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1213_
timestamp 1694700623
transform -1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1694700623
transform -1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1694700623
transform 1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1216_
timestamp 1694700623
transform 1 0 9476 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1217_
timestamp 1694700623
transform 1 0 8188 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1218_
timestamp 1694700623
transform 1 0 8188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1219_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9292 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1220_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8924 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1694700623
transform -1 0 10028 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9752 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1223_
timestamp 1694700623
transform 1 0 8924 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1224_
timestamp 1694700623
transform 1 0 12052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1694700623
transform 1 0 12052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1694700623
transform 1 0 11500 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 1694700623
transform 1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1228_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10120 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_2  _1229_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8832 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_1  _1230_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1231_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6440 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _1232_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1694700623
transform 1 0 5336 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1234_
timestamp 1694700623
transform 1 0 4968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1235_
timestamp 1694700623
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _1236_
timestamp 1694700623
transform -1 0 3220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1694700623
transform -1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1238_
timestamp 1694700623
transform -1 0 2668 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1239_
timestamp 1694700623
transform -1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1240_
timestamp 1694700623
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_4  _1241_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3220 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_2  _1242_
timestamp 1694700623
transform -1 0 3496 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1694700623
transform -1 0 3128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1244_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3680 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _1245_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9844 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o32ai_1  _1246_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10856 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1247_
timestamp 1694700623
transform 1 0 7636 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1248_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7820 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1249_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7360 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1250_
timestamp 1694700623
transform -1 0 7544 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1251_
timestamp 1694700623
transform 1 0 2208 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1694700623
transform 1 0 3864 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1253_
timestamp 1694700623
transform 1 0 5060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1254_
timestamp 1694700623
transform -1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1255_
timestamp 1694700623
transform 1 0 5612 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1256_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3956 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1257_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4232 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1258_
timestamp 1694700623
transform 1 0 4048 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1259_
timestamp 1694700623
transform 1 0 1840 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_4  _1260_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1472 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _1261_
timestamp 1694700623
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1262_
timestamp 1694700623
transform 1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1694700623
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1264_
timestamp 1694700623
transform 1 0 7452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1265_
timestamp 1694700623
transform -1 0 8832 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1266_
timestamp 1694700623
transform -1 0 6256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1267_
timestamp 1694700623
transform -1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1268_
timestamp 1694700623
transform -1 0 5244 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1694700623
transform -1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1270_
timestamp 1694700623
transform 1 0 3128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1271_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1272_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3128 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1273_
timestamp 1694700623
transform -1 0 6164 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1694700623
transform 1 0 4048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1275_
timestamp 1694700623
transform 1 0 7912 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1276_
timestamp 1694700623
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1277_
timestamp 1694700623
transform 1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1278_
timestamp 1694700623
transform 1 0 8280 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1279_
timestamp 1694700623
transform 1 0 7176 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1280_
timestamp 1694700623
transform -1 0 6256 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 1694700623
transform -1 0 7176 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1282_
timestamp 1694700623
transform 1 0 4416 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1283_
timestamp 1694700623
transform -1 0 4416 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1284_
timestamp 1694700623
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1285_
timestamp 1694700623
transform 1 0 2208 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1286_
timestamp 1694700623
transform -1 0 4600 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1694700623
transform 1 0 10028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1694700623
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1289_
timestamp 1694700623
transform 1 0 7636 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1290_
timestamp 1694700623
transform -1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1291_
timestamp 1694700623
transform -1 0 7268 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1694700623
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1694700623
transform 1 0 4232 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1294_
timestamp 1694700623
transform -1 0 4416 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1295_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1694700623
transform 1 0 6992 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1297_
timestamp 1694700623
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 1694700623
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1299_
timestamp 1694700623
transform -1 0 5704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1300_
timestamp 1694700623
transform 1 0 5428 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1301_
timestamp 1694700623
transform 1 0 6164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1302_
timestamp 1694700623
transform -1 0 5520 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1303_
timestamp 1694700623
transform 1 0 4508 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _1304_
timestamp 1694700623
transform -1 0 5152 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1305_
timestamp 1694700623
transform -1 0 3588 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1306_
timestamp 1694700623
transform -1 0 5336 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1307_
timestamp 1694700623
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1694700623
transform 1 0 2300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1309_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3496 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1310_
timestamp 1694700623
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1311_
timestamp 1694700623
transform 1 0 6164 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _1312_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_2  _1313_
timestamp 1694700623
transform 1 0 2668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1314_
timestamp 1694700623
transform -1 0 4876 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1315_
timestamp 1694700623
transform 1 0 4784 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1316_
timestamp 1694700623
transform 1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1317_
timestamp 1694700623
transform -1 0 5612 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1694700623
transform 1 0 5428 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1319_
timestamp 1694700623
transform 1 0 5888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1320_
timestamp 1694700623
transform 1 0 7820 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1321_
timestamp 1694700623
transform -1 0 9660 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1322_
timestamp 1694700623
transform -1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1323_
timestamp 1694700623
transform -1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1324_
timestamp 1694700623
transform 1 0 8740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1325_
timestamp 1694700623
transform 1 0 6164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1326_
timestamp 1694700623
transform 1 0 5336 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1327_
timestamp 1694700623
transform 1 0 4508 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1328_
timestamp 1694700623
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1329_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2484 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1330_
timestamp 1694700623
transform 1 0 1656 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1331_
timestamp 1694700623
transform -1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1694700623
transform 1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1333_
timestamp 1694700623
transform -1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1334_
timestamp 1694700623
transform 1 0 4600 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1335_
timestamp 1694700623
transform 1 0 3956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1694700623
transform 1 0 3772 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1337_
timestamp 1694700623
transform 1 0 2760 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1694700623
transform -1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1694700623
transform -1 0 3588 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1340_
timestamp 1694700623
transform 1 0 2576 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1694700623
transform -1 0 2576 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1694700623
transform -1 0 2300 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1343_
timestamp 1694700623
transform 1 0 2116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1694700623
transform 1 0 2208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1694700623
transform 1 0 2300 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2300 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1694700623
transform 1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1348_
timestamp 1694700623
transform -1 0 4508 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1349_
timestamp 1694700623
transform 1 0 4784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1350_
timestamp 1694700623
transform 1 0 4324 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1694700623
transform -1 0 4692 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1352_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1353_
timestamp 1694700623
transform -1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1354_
timestamp 1694700623
transform 1 0 3128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1694700623
transform -1 0 3128 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1694700623
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1357_
timestamp 1694700623
transform 1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1358_
timestamp 1694700623
transform 1 0 4140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1359_
timestamp 1694700623
transform 1 0 6440 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1694700623
transform -1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1361_
timestamp 1694700623
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1362_
timestamp 1694700623
transform 1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1694700623
transform 1 0 8648 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1364_
timestamp 1694700623
transform 1 0 9016 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1694700623
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1694700623
transform -1 0 11960 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1694700623
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1694700623
transform 1 0 12788 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1694700623
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1694700623
transform -1 0 12880 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1694700623
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1372_
timestamp 1694700623
transform 1 0 12236 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1694700623
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1374_
timestamp 1694700623
transform 1 0 12788 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1694700623
transform 1 0 12880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1376_
timestamp 1694700623
transform 1 0 13156 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1694700623
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1378_
timestamp 1694700623
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1379_
timestamp 1694700623
transform -1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1380_
timestamp 1694700623
transform -1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1694700623
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1382_
timestamp 1694700623
transform 1 0 17664 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1694700623
transform -1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1384_
timestamp 1694700623
transform 1 0 20240 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1385_
timestamp 1694700623
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1386_
timestamp 1694700623
transform 1 0 21528 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1387_
timestamp 1694700623
transform 1 0 22356 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1388_
timestamp 1694700623
transform 1 0 23000 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1694700623
transform -1 0 23920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1390_
timestamp 1694700623
transform 1 0 23552 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1694700623
transform -1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1694700623
transform 1 0 14536 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1694700623
transform -1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1694700623
transform 1 0 17020 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1694700623
transform -1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1694700623
transform -1 0 19688 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1397_
timestamp 1694700623
transform 1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1398_
timestamp 1694700623
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1694700623
transform 1 0 7820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1400_
timestamp 1694700623
transform 1 0 8924 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1694700623
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1402_
timestamp 1694700623
transform -1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1403_
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1404_
timestamp 1694700623
transform -1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1694700623
transform 1 0 14628 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1406_
timestamp 1694700623
transform -1 0 15824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1694700623
transform 1 0 18124 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1694700623
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1694700623
transform 1 0 20332 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1694700623
transform -1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1411_
timestamp 1694700623
transform 1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1412_
timestamp 1694700623
transform -1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1413_
timestamp 1694700623
transform 1 0 23276 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1694700623
transform 1 0 23552 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1415_
timestamp 1694700623
transform 1 0 24656 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1694700623
transform -1 0 25484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1417_
timestamp 1694700623
transform 1 0 18032 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1418_
timestamp 1694700623
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1419_
timestamp 1694700623
transform -1 0 14904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1420_
timestamp 1694700623
transform 1 0 19688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1421_
timestamp 1694700623
transform -1 0 20240 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1694700623
transform 1 0 20792 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1423_
timestamp 1694700623
transform -1 0 21528 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1424_
timestamp 1694700623
transform 1 0 23184 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1425_
timestamp 1694700623
transform -1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1426_
timestamp 1694700623
transform 1 0 24472 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1694700623
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1428_
timestamp 1694700623
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1694700623
transform -1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1694700623
transform -1 0 15824 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1431_
timestamp 1694700623
transform -1 0 14996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1432_
timestamp 1694700623
transform -1 0 15088 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1694700623
transform 1 0 14168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1434_
timestamp 1694700623
transform -1 0 14628 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1435_
timestamp 1694700623
transform 1 0 7452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1436_
timestamp 1694700623
transform -1 0 8648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1694700623
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1438_
timestamp 1694700623
transform 1 0 8740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1694700623
transform -1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1440_
timestamp 1694700623
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1694700623
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1442_
timestamp 1694700623
transform 1 0 14536 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1694700623
transform 1 0 14628 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1444_
timestamp 1694700623
transform 1 0 16008 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1694700623
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1694700623
transform -1 0 17756 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1694700623
transform 1 0 16560 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1448_
timestamp 1694700623
transform 1 0 13432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1449_
timestamp 1694700623
transform -1 0 17756 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1694700623
transform -1 0 17296 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1451_
timestamp 1694700623
transform -1 0 16652 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1452_
timestamp 1694700623
transform 1 0 15640 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1453_
timestamp 1694700623
transform 1 0 15272 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1694700623
transform 1 0 15548 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1455_
timestamp 1694700623
transform 1 0 16836 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1694700623
transform 1 0 17756 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1457_
timestamp 1694700623
transform -1 0 19688 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1694700623
transform -1 0 18768 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1459_
timestamp 1694700623
transform -1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1694700623
transform 1 0 19596 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1694700623
transform 1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1462_
timestamp 1694700623
transform -1 0 14628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1694700623
transform 1 0 13616 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1464_
timestamp 1694700623
transform 1 0 14168 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1694700623
transform -1 0 14996 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1466_
timestamp 1694700623
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1694700623
transform -1 0 17664 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1694700623
transform -1 0 19412 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1694700623
transform -1 0 19780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1694700623
transform 1 0 20240 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1694700623
transform 1 0 20700 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1472_
timestamp 1694700623
transform 1 0 21068 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1694700623
transform -1 0 21712 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1474_
timestamp 1694700623
transform 1 0 21712 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1694700623
transform 1 0 23736 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1476_
timestamp 1694700623
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1694700623
transform -1 0 23644 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1478_
timestamp 1694700623
transform 1 0 23184 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1694700623
transform -1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1694700623
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1694700623
transform -1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1694700623
transform 1 0 19872 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1694700623
transform -1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1694700623
transform 1 0 21068 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1694700623
transform -1 0 21528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1486_
timestamp 1694700623
transform 1 0 23092 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1694700623
transform -1 0 23920 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1488_
timestamp 1694700623
transform 1 0 12696 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1489_
timestamp 1694700623
transform -1 0 25300 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1694700623
transform -1 0 24932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1491_
timestamp 1694700623
transform 1 0 25208 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1694700623
transform -1 0 26036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1694700623
transform -1 0 20148 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1694700623
transform -1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1495_
timestamp 1694700623
transform 1 0 20148 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1694700623
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 1694700623
transform 1 0 21160 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1694700623
transform -1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1499_
timestamp 1694700623
transform 1 0 23092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1694700623
transform -1 0 23920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1501_
timestamp 1694700623
transform -1 0 25484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1694700623
transform 1 0 24748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1503_
timestamp 1694700623
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1694700623
transform -1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1505_
timestamp 1694700623
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1694700623
transform -1 0 26772 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1694700623
transform -1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1694700623
transform 1 0 26680 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1509_
timestamp 1694700623
transform -1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1694700623
transform 1 0 25944 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1511_
timestamp 1694700623
transform 1 0 26404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1512_
timestamp 1694700623
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1513_
timestamp 1694700623
transform 1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1514_
timestamp 1694700623
transform -1 0 24840 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1515_
timestamp 1694700623
transform -1 0 24564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1516_
timestamp 1694700623
transform 1 0 25484 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1694700623
transform -1 0 26312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1518_
timestamp 1694700623
transform 1 0 16928 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1694700623
transform 1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1694700623
transform 1 0 17388 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1521_
timestamp 1694700623
transform 1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 1694700623
transform -1 0 13892 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1694700623
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1524_
timestamp 1694700623
transform -1 0 10120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1694700623
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1526_
timestamp 1694700623
transform -1 0 10856 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1694700623
transform -1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1528_
timestamp 1694700623
transform 1 0 12052 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1529_
timestamp 1694700623
transform -1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1530_
timestamp 1694700623
transform 1 0 16744 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1694700623
transform -1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1532_
timestamp 1694700623
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1533_
timestamp 1694700623
transform -1 0 19688 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1534_
timestamp 1694700623
transform -1 0 19228 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1535_
timestamp 1694700623
transform 1 0 20700 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1694700623
transform 1 0 21252 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1537_
timestamp 1694700623
transform 1 0 21804 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1538_
timestamp 1694700623
transform -1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1539_
timestamp 1694700623
transform -1 0 24196 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1694700623
transform -1 0 24012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1541_
timestamp 1694700623
transform 1 0 21804 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1694700623
transform -1 0 21528 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1543_
timestamp 1694700623
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1544_
timestamp 1694700623
transform 1 0 16928 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1694700623
transform -1 0 17480 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1694700623
transform 1 0 18492 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1694700623
transform -1 0 19228 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1548_
timestamp 1694700623
transform 1 0 17664 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1694700623
transform -1 0 18124 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1694700623
transform -1 0 15824 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1694700623
transform 1 0 15180 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1694700623
transform -1 0 14352 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1694700623
transform -1 0 13524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1554_
timestamp 1694700623
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1694700623
transform 1 0 14628 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1556_
timestamp 1694700623
transform -1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1557_
timestamp 1694700623
transform 1 0 14904 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1558_
timestamp 1694700623
transform -1 0 15916 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1694700623
transform 1 0 15364 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1560_
timestamp 1694700623
transform -1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1694700623
transform 1 0 12788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1562_
timestamp 1694700623
transform -1 0 13340 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1694700623
transform -1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1564_
timestamp 1694700623
transform 1 0 11684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1694700623
transform -1 0 12512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1566_
timestamp 1694700623
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 1694700623
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1568_
timestamp 1694700623
transform 1 0 14168 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 1694700623
transform -1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 1694700623
transform 1 0 15456 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1694700623
transform -1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1572_
timestamp 1694700623
transform 1 0 17848 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 1694700623
transform -1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1694700623
transform 1 0 19964 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1694700623
transform -1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1576_
timestamp 1694700623
transform 1 0 13432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1577_
timestamp 1694700623
transform 1 0 20884 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1694700623
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1579_
timestamp 1694700623
transform -1 0 19688 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1694700623
transform -1 0 19044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 1694700623
transform 1 0 16100 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1694700623
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1583_
timestamp 1694700623
transform 1 0 17664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1694700623
transform -1 0 18768 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 1694700623
transform 1 0 20608 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1694700623
transform -1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1587_
timestamp 1694700623
transform 1 0 23736 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1694700623
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1589_
timestamp 1694700623
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1590_
timestamp 1694700623
transform 1 0 19412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1591_
timestamp 1694700623
transform -1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1592_
timestamp 1694700623
transform -1 0 21620 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1593_
timestamp 1694700623
transform -1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1594_
timestamp 1694700623
transform 1 0 16928 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1595_
timestamp 1694700623
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1596_
timestamp 1694700623
transform 1 0 18308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1694700623
transform -1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 1694700623
transform 1 0 20608 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1694700623
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1694700623
transform 1 0 22172 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1601_
timestamp 1694700623
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1602_
timestamp 1694700623
transform 1 0 23276 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1603_
timestamp 1694700623
transform -1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1604_
timestamp 1694700623
transform 1 0 19136 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1605_
timestamp 1694700623
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1606_
timestamp 1694700623
transform -1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1607_
timestamp 1694700623
transform 1 0 12972 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1608_
timestamp 1694700623
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1609_
timestamp 1694700623
transform 1 0 14444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1694700623
transform 1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1611_
timestamp 1694700623
transform 1 0 7636 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1694700623
transform 1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1613_
timestamp 1694700623
transform 1 0 8096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1615_
timestamp 1694700623
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1694700623
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1617_
timestamp 1694700623
transform 1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1694700623
transform -1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1619_
timestamp 1694700623
transform 1 0 13524 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1620_
timestamp 1694700623
transform -1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1621_
timestamp 1694700623
transform -1 0 14996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1622_
timestamp 1694700623
transform -1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1623_
timestamp 1694700623
transform 1 0 7912 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1694700623
transform 1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1625_
timestamp 1694700623
transform -1 0 10120 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1694700623
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1627_
timestamp 1694700623
transform 1 0 10212 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1628_
timestamp 1694700623
transform -1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1629_
timestamp 1694700623
transform 1 0 11592 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1630_
timestamp 1694700623
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1631_
timestamp 1694700623
transform 1 0 12328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1694700623
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1633_
timestamp 1694700623
transform -1 0 14628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1635_
timestamp 1694700623
transform -1 0 11132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1636_
timestamp 1694700623
transform 1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1637_
timestamp 1694700623
transform -1 0 7360 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1638_
timestamp 1694700623
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1639_
timestamp 1694700623
transform -1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1640_
timestamp 1694700623
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1694700623
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1642_
timestamp 1694700623
transform -1 0 6992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1643_
timestamp 1694700623
transform 1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1644_
timestamp 1694700623
transform -1 0 5796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1694700623
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1646_
timestamp 1694700623
transform -1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1694700623
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1648_
timestamp 1694700623
transform 1 0 5336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1694700623
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1650_
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1694700623
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1652_
timestamp 1694700623
transform -1 0 3680 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1694700623
transform -1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1654_
timestamp 1694700623
transform 1 0 5152 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1655_
timestamp 1694700623
transform 1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1656_
timestamp 1694700623
transform 1 0 3956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1657_
timestamp 1694700623
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1658_
timestamp 1694700623
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1694700623
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1660_
timestamp 1694700623
transform -1 0 7176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1694700623
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1662_
timestamp 1694700623
transform -1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1694700623
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1664_
timestamp 1694700623
transform 1 0 9844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1665_
timestamp 1694700623
transform -1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1666_
timestamp 1694700623
transform -1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1667_
timestamp 1694700623
transform -1 0 12144 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1694700623
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 1694700623
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1694700623
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1671_
timestamp 1694700623
transform -1 0 17204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1694700623
transform -1 0 16560 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1673_
timestamp 1694700623
transform 1 0 18768 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1694700623
transform -1 0 19688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1675_
timestamp 1694700623
transform -1 0 22356 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1694700623
transform -1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1677_
timestamp 1694700623
transform 1 0 22264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1694700623
transform -1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1679_
timestamp 1694700623
transform -1 0 22448 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1694700623
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1681_
timestamp 1694700623
transform -1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1694700623
transform -1 0 19688 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1683_
timestamp 1694700623
transform -1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1694700623
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1685_
timestamp 1694700623
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1694700623
transform -1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1694700623
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1688_
timestamp 1694700623
transform 1 0 20608 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1694700623
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1690_
timestamp 1694700623
transform -1 0 23184 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1694700623
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1692_
timestamp 1694700623
transform 1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1693_
timestamp 1694700623
transform -1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1694_
timestamp 1694700623
transform 1 0 24564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1694700623
transform -1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1696_
timestamp 1694700623
transform 1 0 25576 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1697_
timestamp 1694700623
transform 1 0 26128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1698_
timestamp 1694700623
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1694700623
transform -1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1700_
timestamp 1694700623
transform 1 0 23828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1694700623
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1702_
timestamp 1694700623
transform -1 0 24932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1703_
timestamp 1694700623
transform -1 0 24288 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1704_
timestamp 1694700623
transform -1 0 26404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1705_
timestamp 1694700623
transform -1 0 25392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1706_
timestamp 1694700623
transform -1 0 27508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1694700623
transform -1 0 26864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1708_
timestamp 1694700623
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1709_
timestamp 1694700623
transform 1 0 27140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1694700623
transform -1 0 27508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1711_
timestamp 1694700623
transform 1 0 25576 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1694700623
transform -1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1713_
timestamp 1694700623
transform 1 0 25300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1694700623
transform 1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1715_
timestamp 1694700623
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1716_
timestamp 1694700623
transform 1 0 27508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1717_
timestamp 1694700623
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1694700623
transform 1 0 27416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1719_
timestamp 1694700623
transform 1 0 26864 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1694700623
transform -1 0 27600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1721_
timestamp 1694700623
transform 1 0 27324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1694700623
transform -1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1723_
timestamp 1694700623
transform 1 0 25668 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1694700623
transform -1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1725_
timestamp 1694700623
transform -1 0 25760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1694700623
transform -1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1727_
timestamp 1694700623
transform 1 0 24840 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1694700623
transform -1 0 25668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1729_
timestamp 1694700623
transform -1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1730_
timestamp 1694700623
transform 1 0 16652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1694700623
transform -1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1732_
timestamp 1694700623
transform 1 0 15272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1733_
timestamp 1694700623
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1734_
timestamp 1694700623
transform -1 0 16376 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1735_
timestamp 1694700623
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1736_
timestamp 1694700623
transform -1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1694700623
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1738_
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1739_
timestamp 1694700623
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1740_
timestamp 1694700623
transform 1 0 9384 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1741_
timestamp 1694700623
transform -1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1742_
timestamp 1694700623
transform 1 0 11500 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1743_
timestamp 1694700623
transform -1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1744_
timestamp 1694700623
transform 1 0 13616 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1745_
timestamp 1694700623
transform -1 0 14628 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1746_
timestamp 1694700623
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1694700623
transform -1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1748_
timestamp 1694700623
transform -1 0 11316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1694700623
transform 1 0 7176 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1750_
timestamp 1694700623
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1694700623
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1752_
timestamp 1694700623
transform 1 0 5244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1694700623
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1754_
timestamp 1694700623
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1694700623
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1756_
timestamp 1694700623
transform -1 0 6900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1757_
timestamp 1694700623
transform -1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1758_
timestamp 1694700623
transform 1 0 12144 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1759_
timestamp 1694700623
transform -1 0 13064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1760_
timestamp 1694700623
transform -1 0 4324 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1761_
timestamp 1694700623
transform 1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1762_
timestamp 1694700623
transform 1 0 5612 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1763_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6256 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1764_
timestamp 1694700623
transform -1 0 6808 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1765_
timestamp 1694700623
transform -1 0 5612 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _1766_
timestamp 1694700623
transform 1 0 6900 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1767_
timestamp 1694700623
transform 1 0 6624 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1768_
timestamp 1694700623
transform 1 0 4784 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1769_
timestamp 1694700623
transform -1 0 6256 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _1770_
timestamp 1694700623
transform -1 0 10396 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1771_
timestamp 1694700623
transform 1 0 10396 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1772_
timestamp 1694700623
transform -1 0 10120 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1773_
timestamp 1694700623
transform 1 0 9752 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1774_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4324 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _1775_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1776_
timestamp 1694700623
transform -1 0 2300 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1777_
timestamp 1694700623
transform 1 0 1564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1778_
timestamp 1694700623
transform -1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1779_
timestamp 1694700623
transform 1 0 2392 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1780_
timestamp 1694700623
transform 1 0 1840 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1781_
timestamp 1694700623
transform 1 0 2024 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1782_
timestamp 1694700623
transform 1 0 3220 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1694700623
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1784_
timestamp 1694700623
transform -1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1785_
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1786_
timestamp 1694700623
transform 1 0 2852 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1787_
timestamp 1694700623
transform 1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1788_
timestamp 1694700623
transform -1 0 4232 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1789_
timestamp 1694700623
transform 1 0 3036 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1790_
timestamp 1694700623
transform -1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1791_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4784 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1792_
timestamp 1694700623
transform 1 0 4784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1793_
timestamp 1694700623
transform 1 0 4140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1794_
timestamp 1694700623
transform 1 0 6900 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1795_
timestamp 1694700623
transform 1 0 5796 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1796_
timestamp 1694700623
transform -1 0 6900 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1797_
timestamp 1694700623
transform -1 0 5980 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1798_
timestamp 1694700623
transform 1 0 4600 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1799_
timestamp 1694700623
transform 1 0 5244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1800_
timestamp 1694700623
transform 1 0 4876 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1801_
timestamp 1694700623
transform 1 0 7268 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1802_
timestamp 1694700623
transform -1 0 7084 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1694700623
transform 1 0 6348 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1804_
timestamp 1694700623
transform -1 0 7452 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1805_
timestamp 1694700623
transform 1 0 7452 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1806_
timestamp 1694700623
transform -1 0 9936 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1807_
timestamp 1694700623
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1808_
timestamp 1694700623
transform -1 0 9476 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1809_
timestamp 1694700623
transform -1 0 9200 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1810_
timestamp 1694700623
transform -1 0 7268 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1811_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1694700623
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1694700623
transform 1 0 7912 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1694700623
transform 1 0 9568 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1694700623
transform 1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1694700623
transform 1 0 11868 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1694700623
transform 1 0 11684 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1694700623
transform 1 0 12328 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1694700623
transform 1 0 12512 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1694700623
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1694700623
transform 1 0 14720 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1694700623
transform 1 0 18308 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1694700623
transform 1 0 20792 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1694700623
transform 1 0 22080 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1694700623
transform -1 0 25116 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1694700623
transform -1 0 25852 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1694700623
transform 1 0 15088 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1694700623
transform 1 0 17848 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1694700623
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1694700623
transform 1 0 9660 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1694700623
transform 1 0 12236 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1694700623
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1694700623
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1694700623
transform 1 0 21344 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1694700623
transform -1 0 24932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1694700623
transform 1 0 23184 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1694700623
transform -1 0 25852 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1694700623
transform 1 0 18492 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1694700623
transform 1 0 19964 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1694700623
transform 1 0 21344 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1694700623
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1694700623
transform -1 0 26312 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1694700623
transform -1 0 26772 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1694700623
transform 1 0 14996 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1694700623
transform 1 0 13616 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1694700623
transform 1 0 7084 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1694700623
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1694700623
transform 1 0 9660 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1694700623
transform 1 0 12880 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1694700623
transform 1 0 14536 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1694700623
transform 1 0 16100 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1694700623
transform 1 0 16100 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1694700623
transform -1 0 18308 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1694700623
transform 1 0 14904 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1694700623
transform 1 0 15364 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1694700623
transform 1 0 17296 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1694700623
transform 1 0 18768 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1694700623
transform 1 0 19412 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1694700623
transform 1 0 13248 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1694700623
transform 1 0 14628 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1694700623
transform 1 0 17756 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1694700623
transform 1 0 19412 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1694700623
transform 1 0 20240 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1694700623
transform 1 0 21804 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1694700623
transform -1 0 23736 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1694700623
transform -1 0 24564 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1694700623
transform -1 0 24840 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1694700623
transform -1 0 23276 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1694700623
transform 1 0 20332 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1694700623
transform 1 0 21804 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1694700623
transform 1 0 24380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1694700623
transform 1 0 24932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1694700623
transform 1 0 26312 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1694700623
transform 1 0 19780 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1694700623
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1694700623
transform 1 0 21896 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1694700623
transform 1 0 23460 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1694700623
transform 1 0 24472 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1694700623
transform 1 0 25208 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1694700623
transform 1 0 26956 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1694700623
transform 1 0 27140 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1694700623
transform 1 0 25852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1694700623
transform 1 0 27140 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1694700623
transform 1 0 24564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1694700623
transform 1 0 25944 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1694700623
transform 1 0 16836 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1694700623
transform -1 0 18492 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1694700623
transform 1 0 8096 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1694700623
transform 1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1694700623
transform 1 0 12512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1694700623
transform 1 0 17296 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1694700623
transform 1 0 19228 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1694700623
transform 1 0 20700 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1694700623
transform 1 0 22172 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1694700623
transform 1 0 24380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1694700623
transform -1 0 22172 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1694700623
transform 1 0 17480 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1694700623
transform 1 0 19228 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1694700623
transform -1 0 18952 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1694700623
transform 1 0 14628 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1694700623
transform 1 0 13524 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1694700623
transform 1 0 13984 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1694700623
transform 1 0 14628 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1694700623
transform 1 0 14904 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1694700623
transform 1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1694700623
transform -1 0 13708 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1694700623
transform -1 0 12604 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1694700623
transform 1 0 12788 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1694700623
transform 1 0 14536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1694700623
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1694700623
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1694700623
transform 1 0 20700 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1694700623
transform 1 0 20700 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1694700623
transform -1 0 19688 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1694700623
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1694700623
transform 1 0 19688 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1694700623
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1694700623
transform 1 0 22816 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1694700623
transform 1 0 19688 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1694700623
transform -1 0 19136 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1694700623
transform 1 0 17112 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1694700623
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1694700623
transform 1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1694700623
transform 1 0 22172 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1694700623
transform -1 0 25116 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1694700623
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1694700623
transform 1 0 13248 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1694700623
transform 1 0 14352 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1694700623
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1694700623
transform 1 0 8556 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1694700623
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1694700623
transform 1 0 14444 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1694700623
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1694700623
transform 1 0 9016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1694700623
transform 1 0 10580 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1694700623
transform 1 0 11408 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1694700623
transform 1 0 12144 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1694700623
transform 1 0 13616 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1694700623
transform 1 0 7636 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1694700623
transform 1 0 6256 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1694700623
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1694700623
transform 1 0 6072 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1694700623
transform 1 0 4232 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1694700623
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1694700623
transform 1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1694700623
transform -1 0 4876 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1694700623
transform 1 0 4508 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1694700623
transform 1 0 6716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1694700623
transform 1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1694700623
transform 1 0 9936 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1694700623
transform 1 0 11960 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1694700623
transform 1 0 14076 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1694700623
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1694700623
transform 1 0 19872 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1694700623
transform 1 0 21804 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1694700623
transform -1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1694700623
transform 1 0 20700 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1694700623
transform -1 0 20700 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1694700623
transform 1 0 17664 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1694700623
transform 1 0 20056 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1694700623
transform 1 0 21160 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1694700623
transform 1 0 22264 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1694700623
transform -1 0 25852 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1694700623
transform -1 0 26404 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1694700623
transform 1 0 25760 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1694700623
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1694700623
transform 1 0 24380 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1694700623
transform 1 0 24380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1694700623
transform 1 0 25392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1694700623
transform 1 0 26864 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1694700623
transform -1 0 28520 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1694700623
transform -1 0 27140 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1694700623
transform 1 0 25576 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1981_
timestamp 1694700623
transform 1 0 27140 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1982_
timestamp 1694700623
transform 1 0 27140 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1983_
timestamp 1694700623
transform 1 0 27140 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1694700623
transform -1 0 28612 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1694700623
transform -1 0 27324 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1986_
timestamp 1694700623
transform -1 0 26772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1987_
timestamp 1694700623
transform -1 0 26220 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1988_
timestamp 1694700623
transform -1 0 18124 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1989_
timestamp 1694700623
transform 1 0 15088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1990_
timestamp 1694700623
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1694700623
transform 1 0 7912 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1694700623
transform 1 0 8924 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1694700623
transform 1 0 9936 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1994_
timestamp 1694700623
transform 1 0 12052 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1995_
timestamp 1694700623
transform 1 0 14720 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1996_
timestamp 1694700623
transform 1 0 17296 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1997_
timestamp 1694700623
transform 1 0 6716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1998_
timestamp 1694700623
transform 1 0 6716 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1999_
timestamp 1694700623
transform -1 0 5980 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2000_
timestamp 1694700623
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2001_
timestamp 1694700623
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2002_
timestamp 1694700623
transform 1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _2003_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2004_
timestamp 1694700623
transform 1 0 5612 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2005_
timestamp 1694700623
transform 1 0 7084 0 1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2006_
timestamp 1694700623
transform 1 0 6348 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2007_
timestamp 1694700623
transform 1 0 10396 0 1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2008_
timestamp 1694700623
transform 1 0 10304 0 1 28288
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _2009_
timestamp 1694700623
transform 1 0 1932 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2010_
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2011_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2012_
timestamp 1694700623
transform -1 0 4416 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2013_
timestamp 1694700623
transform 1 0 2116 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2014_
timestamp 1694700623
transform 1 0 3588 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2015_
timestamp 1694700623
transform 1 0 4784 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2016_
timestamp 1694700623
transform 1 0 4692 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2017_
timestamp 1694700623
transform -1 0 6900 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2018_
timestamp 1694700623
transform 1 0 4140 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2019_
timestamp 1694700623
transform 1 0 4416 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2020_
timestamp 1694700623
transform 1 0 5888 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1694700623
transform 1 0 7360 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1694700623
transform -1 0 10488 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2023_
timestamp 1694700623
transform 1 0 6900 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0380_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6992 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_in[0]
timestamp 1694700623
transform 1 0 6348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net67
timestamp 1694700623
transform 1 0 3772 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.dcdel_capnode_notouch_
timestamp 1694700623
transform -1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1694700623
transform 1 0 2668 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0380_
timestamp 1694700623
transform -1 0 8280 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_io_in[0]
timestamp 1694700623
transform -1 0 7084 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net67
timestamp 1694700623
transform -1 0 5612 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.dcdel_capnode_notouch_
timestamp 1694700623
transform -1 0 3680 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1694700623
transform 1 0 3772 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0380_
timestamp 1694700623
transform 1 0 8280 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_io_in[0]
timestamp 1694700623
transform 1 0 6072 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net67
timestamp 1694700623
transform -1 0 5428 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.dcdel_capnode_notouch_
timestamp 1694700623
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1694700623
transform -1 0 3496 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1694700623
transform -1 0 11132 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout9
timestamp 1694700623
transform 1 0 9660 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1694700623
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1694700623
transform -1 0 8832 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1694700623
transform -1 0 11408 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1694700623
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1694700623
transform -1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout24
timestamp 1694700623
transform -1 0 5152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1694700623
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1694700623
transform -1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1694700623
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout28
timestamp 1694700623
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1694700623
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1694700623
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1694700623
transform -1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout32
timestamp 1694700623
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1694700623
transform 1 0 23184 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 1694700623
transform 1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1694700623
transform -1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 1694700623
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1694700623
transform -1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1694700623
transform -1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1694700623
transform 1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 1694700623
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1694700623
transform -1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1694700623
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1694700623
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1694700623
transform 1 0 17848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1694700623
transform -1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1694700623
transform -1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1694700623
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1694700623
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1694700623
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1694700623
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1694700623
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1694700623
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1694700623
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1694700623
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_101 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10396 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1694700623
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1694700623
transform 1 0 11868 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121
timestamp 1694700623
transform 1 0 12236 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13340 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1694700623
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_157
timestamp 1694700623
transform 1 0 15548 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1694700623
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_178
timestamp 1694700623
transform 1 0 17480 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_190
timestamp 1694700623
transform 1 0 18584 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19228 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_202
timestamp 1694700623
transform 1 0 19688 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_214
timestamp 1694700623
transform 1 0 20792 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1694700623
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_231
timestamp 1694700623
transform 1 0 22356 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_243
timestamp 1694700623
transform 1 0 23460 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1694700623
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1694700623
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1694700623
transform 1 0 25484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1694700623
transform 1 0 26588 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1694700623
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1694700623
transform 1 0 28060 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1694700623
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1694700623
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1694700623
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1694700623
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1694700623
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1694700623
transform 1 0 6348 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_65
timestamp 1694700623
transform 1 0 7084 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_69
timestamp 1694700623
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 1694700623
transform 1 0 7820 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_135
timestamp 1694700623
transform 1 0 13524 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_142
timestamp 1694700623
transform 1 0 14168 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_147
timestamp 1694700623
transform 1 0 14628 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_164
timestamp 1694700623
transform 1 0 16192 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_175
timestamp 1694700623
transform 1 0 17204 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_198
timestamp 1694700623
transform 1 0 19320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_202
timestamp 1694700623
transform 1 0 19688 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_220
timestamp 1694700623
transform 1 0 21344 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_241
timestamp 1694700623
transform 1 0 23276 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_253
timestamp 1694700623
transform 1 0 24380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_265
timestamp 1694700623
transform 1 0 25484 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1694700623
transform 1 0 26588 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1694700623
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_293
timestamp 1694700623
transform 1 0 28060 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1694700623
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1694700623
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1694700623
transform 1 0 5980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1694700623
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1694700623
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_94
timestamp 1694700623
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_100
timestamp 1694700623
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_104
timestamp 1694700623
transform 1 0 10672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_111
timestamp 1694700623
transform 1 0 11316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_144
timestamp 1694700623
transform 1 0 14352 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_152
timestamp 1694700623
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_158
timestamp 1694700623
transform 1 0 15640 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_170
timestamp 1694700623
transform 1 0 16744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_187
timestamp 1694700623
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1694700623
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_229
timestamp 1694700623
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_236
timestamp 1694700623
transform 1 0 22816 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_248
timestamp 1694700623
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1694700623
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1694700623
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1694700623
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_289
timestamp 1694700623
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_297
timestamp 1694700623
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1694700623
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1694700623
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1694700623
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1694700623
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_77
timestamp 1694700623
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_83
timestamp 1694700623
transform 1 0 8740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_95
timestamp 1694700623
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_99
timestamp 1694700623
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1694700623
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1694700623
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_124
timestamp 1694700623
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_136
timestamp 1694700623
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_148
timestamp 1694700623
transform 1 0 14720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_165
timestamp 1694700623
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_169
timestamp 1694700623
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_177
timestamp 1694700623
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_186
timestamp 1694700623
transform 1 0 18216 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_198
timestamp 1694700623
transform 1 0 19320 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_206
timestamp 1694700623
transform 1 0 20056 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1694700623
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1694700623
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_225
timestamp 1694700623
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_248
timestamp 1694700623
transform 1 0 23920 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_260
timestamp 1694700623
transform 1 0 25024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_272
timestamp 1694700623
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1694700623
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_293
timestamp 1694700623
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1694700623
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_41
timestamp 1694700623
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_51
timestamp 1694700623
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_55
timestamp 1694700623
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_72
timestamp 1694700623
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1694700623
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1694700623
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1694700623
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_131
timestamp 1694700623
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1694700623
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_147
timestamp 1694700623
transform 1 0 14628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 1694700623
transform 1 0 15180 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_166
timestamp 1694700623
transform 1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_175
timestamp 1694700623
transform 1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_222
timestamp 1694700623
transform 1 0 21528 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_237
timestamp 1694700623
transform 1 0 22908 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_248
timestamp 1694700623
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1694700623
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1694700623
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1694700623
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_289
timestamp 1694700623
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_297
timestamp 1694700623
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1694700623
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_39
timestamp 1694700623
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_64
timestamp 1694700623
transform 1 0 6992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_70
timestamp 1694700623
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_101
timestamp 1694700623
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1694700623
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_117
timestamp 1694700623
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_185
timestamp 1694700623
transform 1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_193
timestamp 1694700623
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_205
timestamp 1694700623
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_216
timestamp 1694700623
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1694700623
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1694700623
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1694700623
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1694700623
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1694700623
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_293
timestamp 1694700623
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_7
timestamp 1694700623
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 1694700623
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_52
timestamp 1694700623
transform 1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_60
timestamp 1694700623
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_72
timestamp 1694700623
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_101
timestamp 1694700623
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_110
timestamp 1694700623
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_114
timestamp 1694700623
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_118
timestamp 1694700623
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_128
timestamp 1694700623
transform 1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1694700623
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_144
timestamp 1694700623
transform 1 0 14352 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_159
timestamp 1694700623
transform 1 0 15732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_167
timestamp 1694700623
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_175
timestamp 1694700623
transform 1 0 17204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_181
timestamp 1694700623
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1694700623
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1694700623
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_234
timestamp 1694700623
transform 1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1694700623
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1694700623
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1694700623
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1694700623
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_289
timestamp 1694700623
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_297
timestamp 1694700623
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1694700623
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1694700623
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1694700623
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_67
timestamp 1694700623
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_89
timestamp 1694700623
transform 1 0 9292 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_97
timestamp 1694700623
transform 1 0 10028 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_104
timestamp 1694700623
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_119
timestamp 1694700623
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_123
timestamp 1694700623
transform 1 0 12420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_129
timestamp 1694700623
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_151
timestamp 1694700623
transform 1 0 14996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1694700623
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp 1694700623
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_177
timestamp 1694700623
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_186
timestamp 1694700623
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_192
timestamp 1694700623
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_204
timestamp 1694700623
transform 1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1694700623
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1694700623
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_244
timestamp 1694700623
transform 1 0 23552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_252
timestamp 1694700623
transform 1 0 24288 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_258
timestamp 1694700623
transform 1 0 24840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_275
timestamp 1694700623
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1694700623
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1694700623
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_293
timestamp 1694700623
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1694700623
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_50
timestamp 1694700623
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_70
timestamp 1694700623
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1694700623
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1694700623
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1694700623
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_127
timestamp 1694700623
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_160
timestamp 1694700623
transform 1 0 15824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1694700623
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_218
timestamp 1694700623
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_230
timestamp 1694700623
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_242
timestamp 1694700623
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_250
timestamp 1694700623
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_272
timestamp 1694700623
transform 1 0 26128 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_284
timestamp 1694700623
transform 1 0 27232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_296
timestamp 1694700623
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_9
timestamp 1694700623
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_15
timestamp 1694700623
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_21
timestamp 1694700623
transform 1 0 3036 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_25
timestamp 1694700623
transform 1 0 3404 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_33
timestamp 1694700623
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1694700623
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_77
timestamp 1694700623
transform 1 0 8188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 1694700623
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1694700623
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_121
timestamp 1694700623
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_134
timestamp 1694700623
transform 1 0 13432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_142
timestamp 1694700623
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_151
timestamp 1694700623
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_159
timestamp 1694700623
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1694700623
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1694700623
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_177
timestamp 1694700623
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_183
timestamp 1694700623
transform 1 0 17940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_196
timestamp 1694700623
transform 1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_204
timestamp 1694700623
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_220
timestamp 1694700623
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_228
timestamp 1694700623
transform 1 0 22080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_265
timestamp 1694700623
transform 1 0 25484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_275
timestamp 1694700623
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1694700623
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1694700623
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_293
timestamp 1694700623
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_32
timestamp 1694700623
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_44
timestamp 1694700623
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_56
timestamp 1694700623
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_66
timestamp 1694700623
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_98
timestamp 1694700623
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_103
timestamp 1694700623
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_107
timestamp 1694700623
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_114
timestamp 1694700623
transform 1 0 11592 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_126
timestamp 1694700623
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_130
timestamp 1694700623
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1694700623
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_151
timestamp 1694700623
transform 1 0 14996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_163
timestamp 1694700623
transform 1 0 16100 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_171
timestamp 1694700623
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1694700623
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1694700623
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_209
timestamp 1694700623
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_244
timestamp 1694700623
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_253
timestamp 1694700623
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_259
timestamp 1694700623
transform 1 0 24932 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_267
timestamp 1694700623
transform 1 0 25668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_284
timestamp 1694700623
transform 1 0 27232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_296
timestamp 1694700623
transform 1 0 28336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_23
timestamp 1694700623
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 1694700623
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_73
timestamp 1694700623
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_82
timestamp 1694700623
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_94
timestamp 1694700623
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1694700623
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_140
timestamp 1694700623
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1694700623
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1694700623
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_187
timestamp 1694700623
transform 1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_192
timestamp 1694700623
transform 1 0 18768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_198
timestamp 1694700623
transform 1 0 19320 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1694700623
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1694700623
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1694700623
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_225
timestamp 1694700623
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_234
timestamp 1694700623
transform 1 0 22632 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_240
timestamp 1694700623
transform 1 0 23184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_244
timestamp 1694700623
transform 1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_269
timestamp 1694700623
transform 1 0 25852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_273
timestamp 1694700623
transform 1 0 26220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_297
timestamp 1694700623
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_11
timestamp 1694700623
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1694700623
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_62
timestamp 1694700623
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_74
timestamp 1694700623
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1694700623
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_88
timestamp 1694700623
transform 1 0 9200 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_96
timestamp 1694700623
transform 1 0 9936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_107
timestamp 1694700623
transform 1 0 10948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_116
timestamp 1694700623
transform 1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1694700623
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1694700623
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_157
timestamp 1694700623
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_175
timestamp 1694700623
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_223
timestamp 1694700623
transform 1 0 21620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_229
timestamp 1694700623
transform 1 0 22172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_235
timestamp 1694700623
transform 1 0 22724 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1694700623
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1694700623
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_277
timestamp 1694700623
transform 1 0 26588 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_282
timestamp 1694700623
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_294
timestamp 1694700623
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_298
timestamp 1694700623
transform 1 0 28520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_12
timestamp 1694700623
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1694700623
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_63
timestamp 1694700623
transform 1 0 6900 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_97
timestamp 1694700623
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_103
timestamp 1694700623
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1694700623
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_121
timestamp 1694700623
transform 1 0 12236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_133
timestamp 1694700623
transform 1 0 13340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_141
timestamp 1694700623
transform 1 0 14076 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_148
timestamp 1694700623
transform 1 0 14720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1694700623
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1694700623
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_175
timestamp 1694700623
transform 1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_183
timestamp 1694700623
transform 1 0 17940 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_189
timestamp 1694700623
transform 1 0 18492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_201
timestamp 1694700623
transform 1 0 19596 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_206
timestamp 1694700623
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_215
timestamp 1694700623
transform 1 0 20884 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1694700623
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_251
timestamp 1694700623
transform 1 0 24196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_259
timestamp 1694700623
transform 1 0 24932 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_287
timestamp 1694700623
transform 1 0 27508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1694700623
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_45
timestamp 1694700623
transform 1 0 5244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_51
timestamp 1694700623
transform 1 0 5796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1694700623
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_95
timestamp 1694700623
transform 1 0 9844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_125
timestamp 1694700623
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_129
timestamp 1694700623
transform 1 0 12972 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp 1694700623
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_146
timestamp 1694700623
transform 1 0 14536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_150
timestamp 1694700623
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_166
timestamp 1694700623
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_175
timestamp 1694700623
transform 1 0 17204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_179
timestamp 1694700623
transform 1 0 17572 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_186
timestamp 1694700623
transform 1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1694700623
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1694700623
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_209
timestamp 1694700623
transform 1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_217
timestamp 1694700623
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_223
timestamp 1694700623
transform 1 0 21620 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_231
timestamp 1694700623
transform 1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_239
timestamp 1694700623
transform 1 0 23092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_247
timestamp 1694700623
transform 1 0 23828 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_275
timestamp 1694700623
transform 1 0 26404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_296
timestamp 1694700623
transform 1 0 28336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_22
timestamp 1694700623
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_32
timestamp 1694700623
transform 1 0 4048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_62
timestamp 1694700623
transform 1 0 6808 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_77
timestamp 1694700623
transform 1 0 8188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_89
timestamp 1694700623
transform 1 0 9292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_95
timestamp 1694700623
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_104
timestamp 1694700623
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_117
timestamp 1694700623
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_125
timestamp 1694700623
transform 1 0 12604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_157
timestamp 1694700623
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1694700623
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1694700623
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_230
timestamp 1694700623
transform 1 0 22264 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_242
timestamp 1694700623
transform 1 0 23368 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_258
timestamp 1694700623
transform 1 0 24840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_270
timestamp 1694700623
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1694700623
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_290
timestamp 1694700623
transform 1 0 27784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_298
timestamp 1694700623
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1694700623
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_54
timestamp 1694700623
transform 1 0 6072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_62
timestamp 1694700623
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_71
timestamp 1694700623
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1694700623
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_92
timestamp 1694700623
transform 1 0 9568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_100
timestamp 1694700623
transform 1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_108
timestamp 1694700623
transform 1 0 11040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_114
timestamp 1694700623
transform 1 0 11592 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_124
timestamp 1694700623
transform 1 0 12512 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1694700623
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_148
timestamp 1694700623
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_165
timestamp 1694700623
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_176
timestamp 1694700623
transform 1 0 17296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_188
timestamp 1694700623
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_202
timestamp 1694700623
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_234
timestamp 1694700623
transform 1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1694700623
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_261
timestamp 1694700623
transform 1 0 25116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_265
timestamp 1694700623
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_282
timestamp 1694700623
transform 1 0 27048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_7
timestamp 1694700623
transform 1 0 1748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_13
timestamp 1694700623
transform 1 0 2300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_17
timestamp 1694700623
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_36
timestamp 1694700623
transform 1 0 4416 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_77
timestamp 1694700623
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_81
timestamp 1694700623
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_90
timestamp 1694700623
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_94
timestamp 1694700623
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1694700623
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_127
timestamp 1694700623
transform 1 0 12788 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_137
timestamp 1694700623
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1694700623
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_169
timestamp 1694700623
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_188
timestamp 1694700623
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_195
timestamp 1694700623
transform 1 0 19044 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_203
timestamp 1694700623
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_210
timestamp 1694700623
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_214
timestamp 1694700623
transform 1 0 20792 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1694700623
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_225
timestamp 1694700623
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_237
timestamp 1694700623
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_257
timestamp 1694700623
transform 1 0 24748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1694700623
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_287
timestamp 1694700623
transform 1 0 27508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_32
timestamp 1694700623
transform 1 0 4048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_40
timestamp 1694700623
transform 1 0 4784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_63
timestamp 1694700623
transform 1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_100
timestamp 1694700623
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_104
timestamp 1694700623
transform 1 0 10672 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_110
timestamp 1694700623
transform 1 0 11224 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_118
timestamp 1694700623
transform 1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1694700623
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_151
timestamp 1694700623
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_155
timestamp 1694700623
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_177
timestamp 1694700623
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_181
timestamp 1694700623
transform 1 0 17756 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_190
timestamp 1694700623
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_229
timestamp 1694700623
transform 1 0 22172 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_237
timestamp 1694700623
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1694700623
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_273
timestamp 1694700623
transform 1 0 26220 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_279
timestamp 1694700623
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_289
timestamp 1694700623
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_297
timestamp 1694700623
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_20
timestamp 1694700623
transform 1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_28
timestamp 1694700623
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_37
timestamp 1694700623
transform 1 0 4508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1694700623
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1694700623
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_63
timestamp 1694700623
transform 1 0 6900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_71
timestamp 1694700623
transform 1 0 7636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_82
timestamp 1694700623
transform 1 0 8648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_89
timestamp 1694700623
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1694700623
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_121
timestamp 1694700623
transform 1 0 12236 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_130
timestamp 1694700623
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_142
timestamp 1694700623
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_154
timestamp 1694700623
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1694700623
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1694700623
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1694700623
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_193
timestamp 1694700623
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_200
timestamp 1694700623
transform 1 0 19504 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_206
timestamp 1694700623
transform 1 0 20056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_210
timestamp 1694700623
transform 1 0 20424 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_241
timestamp 1694700623
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_253
timestamp 1694700623
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_257
timestamp 1694700623
transform 1 0 24748 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_267
timestamp 1694700623
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1694700623
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_281
timestamp 1694700623
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_6
timestamp 1694700623
transform 1 0 1656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_20
timestamp 1694700623
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_49
timestamp 1694700623
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_53
timestamp 1694700623
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_73
timestamp 1694700623
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1694700623
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1694700623
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_109
timestamp 1694700623
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_117
timestamp 1694700623
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_126
timestamp 1694700623
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 1694700623
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1694700623
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_145
timestamp 1694700623
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_159
timestamp 1694700623
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_166
timestamp 1694700623
transform 1 0 16376 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_172
timestamp 1694700623
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_178
timestamp 1694700623
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1694700623
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_210
timestamp 1694700623
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_214
timestamp 1694700623
transform 1 0 20792 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_220
timestamp 1694700623
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_232
timestamp 1694700623
transform 1 0 22448 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_244
timestamp 1694700623
transform 1 0 23552 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_248
timestamp 1694700623
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_253
timestamp 1694700623
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_259
timestamp 1694700623
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_279
timestamp 1694700623
transform 1 0 26772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_288
timestamp 1694700623
transform 1 0 27600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_296
timestamp 1694700623
transform 1 0 28336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_20
timestamp 1694700623
transform 1 0 2944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_52
timestamp 1694700623
transform 1 0 5888 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_76
timestamp 1694700623
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_84
timestamp 1694700623
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 1694700623
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1694700623
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1694700623
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_124
timestamp 1694700623
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_128
timestamp 1694700623
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_145
timestamp 1694700623
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_178
timestamp 1694700623
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_198
timestamp 1694700623
transform 1 0 19320 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_206
timestamp 1694700623
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1694700623
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_233
timestamp 1694700623
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_237
timestamp 1694700623
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_244
timestamp 1694700623
transform 1 0 23552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_261
timestamp 1694700623
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_268
timestamp 1694700623
transform 1 0 25760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_274
timestamp 1694700623
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1694700623
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_19
timestamp 1694700623
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1694700623
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_56
timestamp 1694700623
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_63
timestamp 1694700623
transform 1 0 6900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_67
timestamp 1694700623
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_109
timestamp 1694700623
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_119
timestamp 1694700623
transform 1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1694700623
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1694700623
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1694700623
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_154
timestamp 1694700623
transform 1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_162
timestamp 1694700623
transform 1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_172
timestamp 1694700623
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_179
timestamp 1694700623
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_187
timestamp 1694700623
transform 1 0 18308 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1694700623
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_207
timestamp 1694700623
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_218
timestamp 1694700623
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1694700623
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_294
timestamp 1694700623
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_298
timestamp 1694700623
transform 1 0 28520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_6
timestamp 1694700623
transform 1 0 1656 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_14
timestamp 1694700623
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_28
timestamp 1694700623
transform 1 0 3680 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_41
timestamp 1694700623
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1694700623
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_69
timestamp 1694700623
transform 1 0 7452 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_76
timestamp 1694700623
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_84
timestamp 1694700623
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp 1694700623
transform 1 0 9476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_99
timestamp 1694700623
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_106
timestamp 1694700623
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1694700623
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_121
timestamp 1694700623
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_133
timestamp 1694700623
transform 1 0 13340 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1694700623
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_215
timestamp 1694700623
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1694700623
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1694700623
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_234
timestamp 1694700623
transform 1 0 22632 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1694700623
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_261
timestamp 1694700623
transform 1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1694700623
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1694700623
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_281
timestamp 1694700623
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_36
timestamp 1694700623
transform 1 0 4416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_43
timestamp 1694700623
transform 1 0 5060 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_48
timestamp 1694700623
transform 1 0 5520 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_60
timestamp 1694700623
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_64
timestamp 1694700623
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1694700623
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_101
timestamp 1694700623
transform 1 0 10396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_119
timestamp 1694700623
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1694700623
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_160
timestamp 1694700623
transform 1 0 15824 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_172
timestamp 1694700623
transform 1 0 16928 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_188
timestamp 1694700623
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_197
timestamp 1694700623
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_213
timestamp 1694700623
transform 1 0 20700 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_230
timestamp 1694700623
transform 1 0 22264 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_238
timestamp 1694700623
transform 1 0 23000 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1694700623
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_253
timestamp 1694700623
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_260
timestamp 1694700623
transform 1 0 25024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_266
timestamp 1694700623
transform 1 0 25576 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_289
timestamp 1694700623
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_297
timestamp 1694700623
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_25
timestamp 1694700623
transform 1 0 3404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_98
timestamp 1694700623
transform 1 0 10120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_107
timestamp 1694700623
transform 1 0 10948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_124
timestamp 1694700623
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_130
timestamp 1694700623
transform 1 0 13064 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_142
timestamp 1694700623
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_150
timestamp 1694700623
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_162
timestamp 1694700623
transform 1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_185
timestamp 1694700623
transform 1 0 18124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_197
timestamp 1694700623
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_203
timestamp 1694700623
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_210
timestamp 1694700623
transform 1 0 20424 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 1694700623
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1694700623
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_242
timestamp 1694700623
transform 1 0 23368 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_265
timestamp 1694700623
transform 1 0 25484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_275
timestamp 1694700623
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1694700623
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_281
timestamp 1694700623
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_287
timestamp 1694700623
transform 1 0 27508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_13
timestamp 1694700623
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_38
timestamp 1694700623
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_45
timestamp 1694700623
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_56
timestamp 1694700623
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_68
timestamp 1694700623
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_72
timestamp 1694700623
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_76
timestamp 1694700623
transform 1 0 8096 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_80
timestamp 1694700623
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1694700623
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_95
timestamp 1694700623
transform 1 0 9844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_103
timestamp 1694700623
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_124
timestamp 1694700623
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1694700623
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1694700623
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_167
timestamp 1694700623
transform 1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_175
timestamp 1694700623
transform 1 0 17204 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1694700623
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_217
timestamp 1694700623
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_223
timestamp 1694700623
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_227
timestamp 1694700623
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_242
timestamp 1694700623
transform 1 0 23368 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1694700623
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_260
timestamp 1694700623
transform 1 0 25024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_272
timestamp 1694700623
transform 1 0 26128 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_280
timestamp 1694700623
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_298
timestamp 1694700623
transform 1 0 28520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_7
timestamp 1694700623
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_25
timestamp 1694700623
transform 1 0 3404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_41
timestamp 1694700623
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_45
timestamp 1694700623
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1694700623
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_71
timestamp 1694700623
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_90
timestamp 1694700623
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1694700623
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_118
timestamp 1694700623
transform 1 0 11960 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_126
timestamp 1694700623
transform 1 0 12696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_133
timestamp 1694700623
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_152
timestamp 1694700623
transform 1 0 15088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1694700623
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1694700623
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_189
timestamp 1694700623
transform 1 0 18492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_201
timestamp 1694700623
transform 1 0 19596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_214
timestamp 1694700623
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 1694700623
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1694700623
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_230
timestamp 1694700623
transform 1 0 22264 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_242
timestamp 1694700623
transform 1 0 23368 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1694700623
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1694700623
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1694700623
transform 1 0 3220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_32
timestamp 1694700623
transform 1 0 4048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp 1694700623
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_99
timestamp 1694700623
transform 1 0 10212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_132
timestamp 1694700623
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_145
timestamp 1694700623
transform 1 0 14444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_157
timestamp 1694700623
transform 1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_172
timestamp 1694700623
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_176
timestamp 1694700623
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_189
timestamp 1694700623
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 1694700623
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_207
timestamp 1694700623
transform 1 0 20148 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_214
timestamp 1694700623
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1694700623
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_253
timestamp 1694700623
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_257
timestamp 1694700623
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_264
timestamp 1694700623
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_268
timestamp 1694700623
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_288
timestamp 1694700623
transform 1 0 27600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_296
timestamp 1694700623
transform 1 0 28336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_28
timestamp 1694700623
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1694700623
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_62
timestamp 1694700623
transform 1 0 6808 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_67
timestamp 1694700623
transform 1 0 7268 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_85
timestamp 1694700623
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_97
timestamp 1694700623
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1694700623
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_113
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1694700623
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_123
timestamp 1694700623
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_127
timestamp 1694700623
transform 1 0 12788 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_149
timestamp 1694700623
transform 1 0 14812 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_158
timestamp 1694700623
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1694700623
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1694700623
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_181
timestamp 1694700623
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1694700623
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_231
timestamp 1694700623
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_235
timestamp 1694700623
transform 1 0 22724 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_241
timestamp 1694700623
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_259
timestamp 1694700623
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_266
timestamp 1694700623
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1694700623
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_289
timestamp 1694700623
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_297
timestamp 1694700623
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 1694700623
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_11
timestamp 1694700623
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1694700623
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_69
timestamp 1694700623
transform 1 0 7452 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_77
timestamp 1694700623
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1694700623
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_113
timestamp 1694700623
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_133
timestamp 1694700623
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_175
timestamp 1694700623
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_187
timestamp 1694700623
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1694700623
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_202
timestamp 1694700623
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_208
timestamp 1694700623
transform 1 0 20240 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_224
timestamp 1694700623
transform 1 0 21712 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_236
timestamp 1694700623
transform 1 0 22816 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 1694700623
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_258
timestamp 1694700623
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_3
timestamp 1694700623
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_16
timestamp 1694700623
transform 1 0 2576 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_23
timestamp 1694700623
transform 1 0 3220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_76
timestamp 1694700623
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_94
timestamp 1694700623
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1694700623
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1694700623
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_128
timestamp 1694700623
transform 1 0 12880 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_136
timestamp 1694700623
transform 1 0 13616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_142
timestamp 1694700623
transform 1 0 14168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_154
timestamp 1694700623
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_161
timestamp 1694700623
transform 1 0 15916 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1694700623
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 1694700623
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_193
timestamp 1694700623
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_201
timestamp 1694700623
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_218
timestamp 1694700623
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_225
timestamp 1694700623
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_232
timestamp 1694700623
transform 1 0 22448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_242
timestamp 1694700623
transform 1 0 23368 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_250
timestamp 1694700623
transform 1 0 24104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1694700623
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_297
timestamp 1694700623
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_3
timestamp 1694700623
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_21
timestamp 1694700623
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1694700623
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1694700623
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1694700623
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_53
timestamp 1694700623
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_59
timestamp 1694700623
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_95
timestamp 1694700623
transform 1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_104
timestamp 1694700623
transform 1 0 10672 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_122
timestamp 1694700623
transform 1 0 12328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_166
timestamp 1694700623
transform 1 0 16376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_177
timestamp 1694700623
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_185
timestamp 1694700623
transform 1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1694700623
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_210
timestamp 1694700623
transform 1 0 20424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_237
timestamp 1694700623
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1694700623
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_286
timestamp 1694700623
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_298
timestamp 1694700623
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_31
timestamp 1694700623
transform 1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_37
timestamp 1694700623
transform 1 0 4508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_46
timestamp 1694700623
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1694700623
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_61
timestamp 1694700623
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_78
timestamp 1694700623
transform 1 0 8280 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_90
timestamp 1694700623
transform 1 0 9384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1694700623
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_121
timestamp 1694700623
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_126
timestamp 1694700623
transform 1 0 12696 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_147
timestamp 1694700623
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_151
timestamp 1694700623
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1694700623
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1694700623
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_183
timestamp 1694700623
transform 1 0 17940 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1694700623
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_212
timestamp 1694700623
transform 1 0 20608 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1694700623
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_237
timestamp 1694700623
transform 1 0 22908 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_265
timestamp 1694700623
transform 1 0 25484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_274
timestamp 1694700623
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1694700623
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_293
timestamp 1694700623
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1694700623
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_55
timestamp 1694700623
transform 1 0 6164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_94
timestamp 1694700623
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_114
timestamp 1694700623
transform 1 0 11592 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_126
timestamp 1694700623
transform 1 0 12696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1694700623
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_167
timestamp 1694700623
transform 1 0 16468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_173
timestamp 1694700623
transform 1 0 17020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1694700623
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_201
timestamp 1694700623
transform 1 0 19596 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_241
timestamp 1694700623
transform 1 0 23276 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1694700623
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1694700623
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_269
timestamp 1694700623
transform 1 0 25852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_281
timestamp 1694700623
transform 1 0 26956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_293
timestamp 1694700623
transform 1 0 28060 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1694700623
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_15
timestamp 1694700623
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_31
timestamp 1694700623
transform 1 0 3956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_45
timestamp 1694700623
transform 1 0 5244 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_51
timestamp 1694700623
transform 1 0 5796 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_80
timestamp 1694700623
transform 1 0 8464 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_92
timestamp 1694700623
transform 1 0 9568 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_104
timestamp 1694700623
transform 1 0 10672 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1694700623
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1694700623
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_144
timestamp 1694700623
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_152
timestamp 1694700623
transform 1 0 15088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_160
timestamp 1694700623
transform 1 0 15824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1694700623
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_179
timestamp 1694700623
transform 1 0 17572 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_187
timestamp 1694700623
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_195
timestamp 1694700623
transform 1 0 19044 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_207
timestamp 1694700623
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_212
timestamp 1694700623
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_237
timestamp 1694700623
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_241
timestamp 1694700623
transform 1 0 23276 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_258
timestamp 1694700623
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_262
timestamp 1694700623
transform 1 0 25208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1694700623
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1694700623
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_293
timestamp 1694700623
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1694700623
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_7
timestamp 1694700623
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_14
timestamp 1694700623
transform 1 0 2392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 1694700623
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1694700623
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 1694700623
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_47
timestamp 1694700623
transform 1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_55
timestamp 1694700623
transform 1 0 6164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_74
timestamp 1694700623
transform 1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_85
timestamp 1694700623
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_96
timestamp 1694700623
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_120
timestamp 1694700623
transform 1 0 12144 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_126
timestamp 1694700623
transform 1 0 12696 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_136
timestamp 1694700623
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_144
timestamp 1694700623
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_154
timestamp 1694700623
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_163
timestamp 1694700623
transform 1 0 16100 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_171
timestamp 1694700623
transform 1 0 16836 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1694700623
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_189
timestamp 1694700623
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_206
timestamp 1694700623
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_222
timestamp 1694700623
transform 1 0 21528 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_234
timestamp 1694700623
transform 1 0 22632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_241
timestamp 1694700623
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_247
timestamp 1694700623
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1694700623
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1694700623
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_261
timestamp 1694700623
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1694700623
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1694700623
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_289
timestamp 1694700623
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_297
timestamp 1694700623
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 1694700623
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_25
timestamp 1694700623
transform 1 0 3404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_42
timestamp 1694700623
transform 1 0 4968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1694700623
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_73
timestamp 1694700623
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_78
timestamp 1694700623
transform 1 0 8280 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_86
timestamp 1694700623
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1694700623
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_120
timestamp 1694700623
transform 1 0 12144 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_126
timestamp 1694700623
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_144
timestamp 1694700623
transform 1 0 14352 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1694700623
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_172
timestamp 1694700623
transform 1 0 16928 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_193
timestamp 1694700623
transform 1 0 18860 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_203
timestamp 1694700623
transform 1 0 19780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1694700623
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_225
timestamp 1694700623
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_246
timestamp 1694700623
transform 1 0 23736 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_258
timestamp 1694700623
transform 1 0 24840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_266
timestamp 1694700623
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_271
timestamp 1694700623
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1694700623
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1694700623
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_293
timestamp 1694700623
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_13
timestamp 1694700623
transform 1 0 2300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_20
timestamp 1694700623
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1694700623
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_61
timestamp 1694700623
transform 1 0 6716 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1694700623
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_97
timestamp 1694700623
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_124
timestamp 1694700623
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_132
timestamp 1694700623
transform 1 0 13248 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1694700623
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_141
timestamp 1694700623
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_150
timestamp 1694700623
transform 1 0 14904 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_179
timestamp 1694700623
transform 1 0 17572 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_185
timestamp 1694700623
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1694700623
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_215
timestamp 1694700623
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_219
timestamp 1694700623
transform 1 0 21252 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_246
timestamp 1694700623
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1694700623
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_290
timestamp 1694700623
transform 1 0 27784 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_298
timestamp 1694700623
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_3
timestamp 1694700623
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1694700623
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_57
timestamp 1694700623
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_67
timestamp 1694700623
transform 1 0 7268 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_88
timestamp 1694700623
transform 1 0 9200 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_100
timestamp 1694700623
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_125
timestamp 1694700623
transform 1 0 12604 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_129
timestamp 1694700623
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_138
timestamp 1694700623
transform 1 0 13800 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_150
timestamp 1694700623
transform 1 0 14904 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_156
timestamp 1694700623
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_169
timestamp 1694700623
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_175
timestamp 1694700623
transform 1 0 17204 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_187
timestamp 1694700623
transform 1 0 18308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_199
timestamp 1694700623
transform 1 0 19412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_219
timestamp 1694700623
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1694700623
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1694700623
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_237
timestamp 1694700623
transform 1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_249
timestamp 1694700623
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_253
timestamp 1694700623
transform 1 0 24380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_260
timestamp 1694700623
transform 1 0 25024 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_268
timestamp 1694700623
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1694700623
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_293
timestamp 1694700623
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_3
timestamp 1694700623
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_11
timestamp 1694700623
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_24
timestamp 1694700623
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_49
timestamp 1694700623
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1694700623
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_104
timestamp 1694700623
transform 1 0 10672 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_111
timestamp 1694700623
transform 1 0 11316 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_123
timestamp 1694700623
transform 1 0 12420 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1694700623
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_148
timestamp 1694700623
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_152
timestamp 1694700623
transform 1 0 15088 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_168
timestamp 1694700623
transform 1 0 16560 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_179
timestamp 1694700623
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_188
timestamp 1694700623
transform 1 0 18400 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1694700623
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_202
timestamp 1694700623
transform 1 0 19688 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_208
timestamp 1694700623
transform 1 0 20240 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_216
timestamp 1694700623
transform 1 0 20976 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_222
timestamp 1694700623
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1694700623
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1694700623
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_269
timestamp 1694700623
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_281
timestamp 1694700623
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_293
timestamp 1694700623
transform 1 0 28060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1694700623
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_7
timestamp 1694700623
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_16
timestamp 1694700623
transform 1 0 2576 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_24
timestamp 1694700623
transform 1 0 3312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_36
timestamp 1694700623
transform 1 0 4416 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_45
timestamp 1694700623
transform 1 0 5244 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1694700623
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_73
timestamp 1694700623
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_77
timestamp 1694700623
transform 1 0 8188 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_98
timestamp 1694700623
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1694700623
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1694700623
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_125
timestamp 1694700623
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_146
timestamp 1694700623
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1694700623
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_179
timestamp 1694700623
transform 1 0 17572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_196
timestamp 1694700623
transform 1 0 19136 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_200
timestamp 1694700623
transform 1 0 19504 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_206
timestamp 1694700623
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_216
timestamp 1694700623
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 1694700623
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_249
timestamp 1694700623
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_255
timestamp 1694700623
transform 1 0 24564 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_275
timestamp 1694700623
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1694700623
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1694700623
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_293
timestamp 1694700623
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_38
timestamp 1694700623
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_59
timestamp 1694700623
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_68
timestamp 1694700623
transform 1 0 7360 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_72
timestamp 1694700623
transform 1 0 7728 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_85
timestamp 1694700623
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_96
timestamp 1694700623
transform 1 0 9936 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_126
timestamp 1694700623
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_130
timestamp 1694700623
transform 1 0 13064 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1694700623
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_149
timestamp 1694700623
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_153
timestamp 1694700623
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_161
timestamp 1694700623
transform 1 0 15916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_173
timestamp 1694700623
transform 1 0 17020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_192
timestamp 1694700623
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_202
timestamp 1694700623
transform 1 0 19688 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_214
timestamp 1694700623
transform 1 0 20792 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_226
timestamp 1694700623
transform 1 0 21896 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_248
timestamp 1694700623
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_269
timestamp 1694700623
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_281
timestamp 1694700623
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_293
timestamp 1694700623
transform 1 0 28060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_3
timestamp 1694700623
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_15
timestamp 1694700623
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_46
timestamp 1694700623
transform 1 0 5336 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1694700623
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_64
timestamp 1694700623
transform 1 0 6992 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_73
timestamp 1694700623
transform 1 0 7820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_84
timestamp 1694700623
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_91
timestamp 1694700623
transform 1 0 9476 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_102
timestamp 1694700623
transform 1 0 10488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_108
timestamp 1694700623
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_118
timestamp 1694700623
transform 1 0 11960 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_122
timestamp 1694700623
transform 1 0 12328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_134
timestamp 1694700623
transform 1 0 13432 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_162
timestamp 1694700623
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_184
timestamp 1694700623
transform 1 0 18032 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_192
timestamp 1694700623
transform 1 0 18768 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1694700623
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_233
timestamp 1694700623
transform 1 0 22540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_245
timestamp 1694700623
transform 1 0 23644 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_249
timestamp 1694700623
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_263
timestamp 1694700623
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1694700623
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1694700623
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1694700623
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_293
timestamp 1694700623
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1694700623
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1694700623
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_35
timestamp 1694700623
transform 1 0 4324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_50
timestamp 1694700623
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_54
timestamp 1694700623
transform 1 0 6072 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_62
timestamp 1694700623
transform 1 0 6808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_95
timestamp 1694700623
transform 1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_122
timestamp 1694700623
transform 1 0 12328 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_150
timestamp 1694700623
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_154
timestamp 1694700623
transform 1 0 15272 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_192
timestamp 1694700623
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_202
timestamp 1694700623
transform 1 0 19688 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_210
timestamp 1694700623
transform 1 0 20424 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1694700623
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_269
timestamp 1694700623
transform 1 0 25852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_281
timestamp 1694700623
transform 1 0 26956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_293
timestamp 1694700623
transform 1 0 28060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_3
timestamp 1694700623
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_46
timestamp 1694700623
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1694700623
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_57
timestamp 1694700623
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_63
timestamp 1694700623
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_70
timestamp 1694700623
transform 1 0 7544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_78
timestamp 1694700623
transform 1 0 8280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_82
timestamp 1694700623
transform 1 0 8648 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_86
timestamp 1694700623
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_90
timestamp 1694700623
transform 1 0 9384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_103
timestamp 1694700623
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1694700623
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1694700623
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_125
timestamp 1694700623
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_131
timestamp 1694700623
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_143
timestamp 1694700623
transform 1 0 14260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_151
timestamp 1694700623
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_169
timestamp 1694700623
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_178
timestamp 1694700623
transform 1 0 17480 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_188
timestamp 1694700623
transform 1 0 18400 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_208
timestamp 1694700623
transform 1 0 20240 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_216
timestamp 1694700623
transform 1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_222
timestamp 1694700623
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_230
timestamp 1694700623
transform 1 0 22264 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_242
timestamp 1694700623
transform 1 0 23368 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_254
timestamp 1694700623
transform 1 0 24472 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_266
timestamp 1694700623
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1694700623
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1694700623
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_293
timestamp 1694700623
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_3
timestamp 1694700623
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1694700623
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 1694700623
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_44
timestamp 1694700623
transform 1 0 5152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_56
timestamp 1694700623
transform 1 0 6256 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_66
timestamp 1694700623
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_78
timestamp 1694700623
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_85
timestamp 1694700623
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_98
timestamp 1694700623
transform 1 0 10120 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_110
timestamp 1694700623
transform 1 0 11224 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1694700623
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1694700623
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1694700623
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_153
timestamp 1694700623
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_160
timestamp 1694700623
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_171
timestamp 1694700623
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1694700623
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_197
timestamp 1694700623
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_203
timestamp 1694700623
transform 1 0 19780 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_211
timestamp 1694700623
transform 1 0 20516 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_229
timestamp 1694700623
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_241
timestamp 1694700623
transform 1 0 23276 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1694700623
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1694700623
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1694700623
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1694700623
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1694700623
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_289
timestamp 1694700623
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_297
timestamp 1694700623
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_18
timestamp 1694700623
transform 1 0 2760 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_27
timestamp 1694700623
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_31
timestamp 1694700623
transform 1 0 3956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_35
timestamp 1694700623
transform 1 0 4324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_43
timestamp 1694700623
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_49
timestamp 1694700623
transform 1 0 5612 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_65
timestamp 1694700623
transform 1 0 7084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_69
timestamp 1694700623
transform 1 0 7452 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_76
timestamp 1694700623
transform 1 0 8096 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_88
timestamp 1694700623
transform 1 0 9200 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_106
timestamp 1694700623
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_113
timestamp 1694700623
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_131
timestamp 1694700623
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_151
timestamp 1694700623
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_160
timestamp 1694700623
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_177
timestamp 1694700623
transform 1 0 17388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_189
timestamp 1694700623
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_193
timestamp 1694700623
transform 1 0 18860 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_215
timestamp 1694700623
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1694700623
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_225
timestamp 1694700623
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_255
timestamp 1694700623
transform 1 0 24564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_267
timestamp 1694700623
transform 1 0 25668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1694700623
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1694700623
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_293
timestamp 1694700623
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_3
timestamp 1694700623
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_15
timestamp 1694700623
transform 1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1694700623
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_44
timestamp 1694700623
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_80
timestamp 1694700623
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_85
timestamp 1694700623
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_90
timestamp 1694700623
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_98
timestamp 1694700623
transform 1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_120
timestamp 1694700623
transform 1 0 12144 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_138
timestamp 1694700623
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_179
timestamp 1694700623
transform 1 0 17572 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_186
timestamp 1694700623
transform 1 0 18216 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1694700623
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_197
timestamp 1694700623
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_206
timestamp 1694700623
transform 1 0 20056 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_216
timestamp 1694700623
transform 1 0 20976 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_222
timestamp 1694700623
transform 1 0 21528 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1694700623
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1694700623
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1694700623
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1694700623
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_289
timestamp 1694700623
transform 1 0 27692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_297
timestamp 1694700623
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_3
timestamp 1694700623
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_15
timestamp 1694700623
transform 1 0 2484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_27
timestamp 1694700623
transform 1 0 3588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1694700623
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1694700623
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_70
timestamp 1694700623
transform 1 0 7544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_82
timestamp 1694700623
transform 1 0 8648 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_93
timestamp 1694700623
transform 1 0 9660 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_99
timestamp 1694700623
transform 1 0 10212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1694700623
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1694700623
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_128
timestamp 1694700623
transform 1 0 12880 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_136
timestamp 1694700623
transform 1 0 13616 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_144
timestamp 1694700623
transform 1 0 14352 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 1694700623
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1694700623
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_169
timestamp 1694700623
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_177
timestamp 1694700623
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_197
timestamp 1694700623
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_201
timestamp 1694700623
transform 1 0 19596 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_205
timestamp 1694700623
transform 1 0 19964 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_241
timestamp 1694700623
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_253
timestamp 1694700623
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_265
timestamp 1694700623
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 1694700623
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1694700623
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_293
timestamp 1694700623
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_3
timestamp 1694700623
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_8
timestamp 1694700623
transform 1 0 1840 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1694700623
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_41
timestamp 1694700623
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_48
timestamp 1694700623
transform 1 0 5520 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_63
timestamp 1694700623
transform 1 0 6900 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_75
timestamp 1694700623
transform 1 0 8004 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_96
timestamp 1694700623
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_119
timestamp 1694700623
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_131
timestamp 1694700623
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_135
timestamp 1694700623
transform 1 0 13524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1694700623
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_141
timestamp 1694700623
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_151
timestamp 1694700623
transform 1 0 14996 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_156
timestamp 1694700623
transform 1 0 15456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_168
timestamp 1694700623
transform 1 0 16560 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_172
timestamp 1694700623
transform 1 0 16928 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_176
timestamp 1694700623
transform 1 0 17296 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_180
timestamp 1694700623
transform 1 0 17664 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_185
timestamp 1694700623
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_193
timestamp 1694700623
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_213
timestamp 1694700623
transform 1 0 20700 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_224
timestamp 1694700623
transform 1 0 21712 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_236
timestamp 1694700623
transform 1 0 22816 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_248
timestamp 1694700623
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1694700623
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1694700623
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1694700623
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_289
timestamp 1694700623
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_297
timestamp 1694700623
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_3
timestamp 1694700623
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_7
timestamp 1694700623
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_13
timestamp 1694700623
transform 1 0 2300 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_24
timestamp 1694700623
transform 1 0 3312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_39
timestamp 1694700623
transform 1 0 4692 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1694700623
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_102
timestamp 1694700623
transform 1 0 10488 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1694700623
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_125
timestamp 1694700623
transform 1 0 12604 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_131
timestamp 1694700623
transform 1 0 13156 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_148
timestamp 1694700623
transform 1 0 14720 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 1694700623
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_197
timestamp 1694700623
transform 1 0 19228 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_215
timestamp 1694700623
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1694700623
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1694700623
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1694700623
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1694700623
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1694700623
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1694700623
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1694700623
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1694700623
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_293
timestamp 1694700623
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_18
timestamp 1694700623
transform 1 0 2760 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1694700623
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_29
timestamp 1694700623
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_35
timestamp 1694700623
transform 1 0 4324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_100
timestamp 1694700623
transform 1 0 10304 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1694700623
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1694700623
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1694700623
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_169
timestamp 1694700623
transform 1 0 16652 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_187
timestamp 1694700623
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1694700623
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1694700623
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1694700623
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1694700623
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1694700623
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1694700623
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1694700623
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1694700623
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1694700623
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1694700623
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_289
timestamp 1694700623
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_297
timestamp 1694700623
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_22
timestamp 1694700623
transform 1 0 3128 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_40
timestamp 1694700623
transform 1 0 4784 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_52
timestamp 1694700623
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_57
timestamp 1694700623
transform 1 0 6348 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_65
timestamp 1694700623
transform 1 0 7084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_77
timestamp 1694700623
transform 1 0 8188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_85
timestamp 1694700623
transform 1 0 8924 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_113
timestamp 1694700623
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_129
timestamp 1694700623
transform 1 0 12972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_141
timestamp 1694700623
transform 1 0 14076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_153
timestamp 1694700623
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_157
timestamp 1694700623
transform 1 0 15548 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1694700623
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1694700623
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1694700623
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1694700623
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1694700623
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1694700623
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1694700623
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1694700623
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1694700623
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1694700623
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1694700623
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1694700623
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1694700623
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1694700623
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1694700623
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_293
timestamp 1694700623
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_3
timestamp 1694700623
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_12
timestamp 1694700623
transform 1 0 2208 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_19
timestamp 1694700623
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1694700623
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_29
timestamp 1694700623
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_44
timestamp 1694700623
transform 1 0 5152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_56
timestamp 1694700623
transform 1 0 6256 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1694700623
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_77
timestamp 1694700623
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_98
timestamp 1694700623
transform 1 0 10120 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_119
timestamp 1694700623
transform 1 0 12052 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_131
timestamp 1694700623
transform 1 0 13156 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1694700623
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1694700623
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1694700623
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1694700623
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1694700623
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1694700623
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1694700623
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1694700623
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1694700623
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1694700623
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1694700623
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1694700623
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1694700623
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1694700623
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1694700623
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1694700623
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_289
timestamp 1694700623
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_297
timestamp 1694700623
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_3
timestamp 1694700623
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_24
timestamp 1694700623
transform 1 0 3312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_45
timestamp 1694700623
transform 1 0 5244 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_62
timestamp 1694700623
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_81
timestamp 1694700623
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_103
timestamp 1694700623
transform 1 0 10580 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 1694700623
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1694700623
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1694700623
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1694700623
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1694700623
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1694700623
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1694700623
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1694700623
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1694700623
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1694700623
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1694700623
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1694700623
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1694700623
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1694700623
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1694700623
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1694700623
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1694700623
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1694700623
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1694700623
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1694700623
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_293
timestamp 1694700623
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1694700623
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1694700623
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1694700623
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_29
timestamp 1694700623
transform 1 0 3772 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_40
timestamp 1694700623
transform 1 0 4784 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_78
timestamp 1694700623
transform 1 0 8280 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_104
timestamp 1694700623
transform 1 0 10672 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_110
timestamp 1694700623
transform 1 0 11224 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_122
timestamp 1694700623
transform 1 0 12328 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_134
timestamp 1694700623
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1694700623
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1694700623
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1694700623
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1694700623
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1694700623
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1694700623
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1694700623
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1694700623
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1694700623
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1694700623
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1694700623
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1694700623
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1694700623
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1694700623
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1694700623
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_289
timestamp 1694700623
transform 1 0 27692 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_297
timestamp 1694700623
transform 1 0 28428 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1694700623
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1694700623
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_27
timestamp 1694700623
transform 1 0 3588 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_29
timestamp 1694700623
transform 1 0 3772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_45
timestamp 1694700623
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_53
timestamp 1694700623
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_67
timestamp 1694700623
transform 1 0 7268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_71
timestamp 1694700623
transform 1 0 7636 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_82
timestamp 1694700623
transform 1 0 8648 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_85
timestamp 1694700623
transform 1 0 8924 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_94
timestamp 1694700623
transform 1 0 9752 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_109
timestamp 1694700623
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1694700623
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1694700623
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_137
timestamp 1694700623
transform 1 0 13708 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_141
timestamp 1694700623
transform 1 0 14076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_153
timestamp 1694700623
transform 1 0 15180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1694700623
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1694700623
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1694700623
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_193
timestamp 1694700623
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_197
timestamp 1694700623
transform 1 0 19228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_209
timestamp 1694700623
transform 1 0 20332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_221
timestamp 1694700623
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1694700623
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1694700623
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_249
timestamp 1694700623
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_253
timestamp 1694700623
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_265
timestamp 1694700623
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_277
timestamp 1694700623
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1694700623
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_293
timestamp 1694700623
transform 1 0 28060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9660 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5888 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1694700623
transform 1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1694700623
transform 1 0 5612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1694700623
transform -1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1694700623
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1694700623
transform -1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1694700623
transform 1 0 8280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1694700623
transform -1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1694700623
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1694700623
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap2
timestamp 1694700623
transform -1 0 15272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap17
timestamp 1694700623
transform -1 0 14352 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap18
timestamp 1694700623
transform 1 0 14260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap20
timestamp 1694700623
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap21
timestamp 1694700623
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap22
timestamp 1694700623
transform -1 0 3036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_58
timestamp 1694700623
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 28888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_59
timestamp 1694700623
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 28888 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_60
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_61
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_62
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_63
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_64
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_65
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_66
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_67
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_68
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_69
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_70
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_71
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_72
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_73
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_74
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_75
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_76
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_77
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_78
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_79
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_80
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_81
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_82
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_83
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_84
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_85
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_86
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1694700623
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_87
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1694700623
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_88
timestamp 1694700623
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1694700623
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_89
timestamp 1694700623
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1694700623
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_90
timestamp 1694700623
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1694700623
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_91
timestamp 1694700623
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1694700623
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_92
timestamp 1694700623
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1694700623
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_93
timestamp 1694700623
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1694700623
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_94
timestamp 1694700623
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1694700623
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_95
timestamp 1694700623
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1694700623
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_96
timestamp 1694700623
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1694700623
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_97
timestamp 1694700623
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1694700623
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_98
timestamp 1694700623
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1694700623
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_99
timestamp 1694700623
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1694700623
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_100
timestamp 1694700623
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1694700623
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_101
timestamp 1694700623
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1694700623
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_102
timestamp 1694700623
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1694700623
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_103
timestamp 1694700623
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1694700623
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_104
timestamp 1694700623
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1694700623
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_105
timestamp 1694700623
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1694700623
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_106
timestamp 1694700623
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1694700623
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_107
timestamp 1694700623
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1694700623
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_108
timestamp 1694700623
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1694700623
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_109
timestamp 1694700623
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1694700623
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_110
timestamp 1694700623
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1694700623
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_111
timestamp 1694700623
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1694700623
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_112
timestamp 1694700623
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1694700623
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_113
timestamp 1694700623
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1694700623
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_114
timestamp 1694700623
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1694700623
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_115
timestamp 1694700623
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1694700623
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_116 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_117
timestamp 1694700623
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_118
timestamp 1694700623
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_119
timestamp 1694700623
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_120
timestamp 1694700623
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_121
timestamp 1694700623
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_122
timestamp 1694700623
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_123
timestamp 1694700623
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_124
timestamp 1694700623
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_125
timestamp 1694700623
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_126
timestamp 1694700623
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_127
timestamp 1694700623
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_128
timestamp 1694700623
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_129
timestamp 1694700623
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_130
timestamp 1694700623
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_131
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_132
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_133
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_134
timestamp 1694700623
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_135
timestamp 1694700623
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_136
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_137
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_138
timestamp 1694700623
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_139
timestamp 1694700623
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_140
timestamp 1694700623
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_141
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_142
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_143
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_144
timestamp 1694700623
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_145
timestamp 1694700623
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_146
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_147
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_148
timestamp 1694700623
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_149
timestamp 1694700623
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_150
timestamp 1694700623
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_151
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_152
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_153
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_154
timestamp 1694700623
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_155
timestamp 1694700623
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_156
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_157
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_158
timestamp 1694700623
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_159
timestamp 1694700623
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_160
timestamp 1694700623
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_161
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_162
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_163
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_164
timestamp 1694700623
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_165
timestamp 1694700623
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_166
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_167
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_168
timestamp 1694700623
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_169
timestamp 1694700623
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_170
timestamp 1694700623
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_171
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_172
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_173
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_174
timestamp 1694700623
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_175
timestamp 1694700623
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_176
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_177
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_178
timestamp 1694700623
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_179
timestamp 1694700623
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_180
timestamp 1694700623
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_181
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_182
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_183
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_184
timestamp 1694700623
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_185
timestamp 1694700623
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_186
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_187
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_188
timestamp 1694700623
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_189
timestamp 1694700623
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_190
timestamp 1694700623
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_191
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_192
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_193
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_194
timestamp 1694700623
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_195
timestamp 1694700623
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_196
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_197
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_198
timestamp 1694700623
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_199
timestamp 1694700623
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_200
timestamp 1694700623
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_201
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_202
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_203
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_204
timestamp 1694700623
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_205
timestamp 1694700623
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_206
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_207
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_208
timestamp 1694700623
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_209
timestamp 1694700623
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_210
timestamp 1694700623
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_211
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_212
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_213
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_214
timestamp 1694700623
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_215
timestamp 1694700623
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_216
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_217
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_218
timestamp 1694700623
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_219
timestamp 1694700623
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_220
timestamp 1694700623
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_221
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_222
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_223
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_224
timestamp 1694700623
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_225
timestamp 1694700623
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_226
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_227
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_228
timestamp 1694700623
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_229
timestamp 1694700623
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_230
timestamp 1694700623
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_231
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_232
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_233
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_234
timestamp 1694700623
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_235
timestamp 1694700623
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_236
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_237
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_238
timestamp 1694700623
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_239
timestamp 1694700623
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_240
timestamp 1694700623
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_241
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_242
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_243
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_244
timestamp 1694700623
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_245
timestamp 1694700623
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_246
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_247
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_248
timestamp 1694700623
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_249
timestamp 1694700623
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_250
timestamp 1694700623
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_251
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_252
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_253
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_254
timestamp 1694700623
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_255
timestamp 1694700623
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_256
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_257
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_258
timestamp 1694700623
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_259
timestamp 1694700623
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_260
timestamp 1694700623
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_261
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_262
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_263
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_264
timestamp 1694700623
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_265
timestamp 1694700623
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_266
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_267
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_268
timestamp 1694700623
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_269
timestamp 1694700623
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_270
timestamp 1694700623
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_271
timestamp 1694700623
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_272
timestamp 1694700623
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_273
timestamp 1694700623
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_274
timestamp 1694700623
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_275
timestamp 1694700623
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_276
timestamp 1694700623
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_277
timestamp 1694700623
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_278
timestamp 1694700623
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_279
timestamp 1694700623
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_280
timestamp 1694700623
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_281
timestamp 1694700623
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_282
timestamp 1694700623
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_283
timestamp 1694700623
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_284
timestamp 1694700623
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_285
timestamp 1694700623
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_286
timestamp 1694700623
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_287
timestamp 1694700623
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_288
timestamp 1694700623
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_289
timestamp 1694700623
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_290
timestamp 1694700623
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_291
timestamp 1694700623
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_292
timestamp 1694700623
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_293
timestamp 1694700623
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_294
timestamp 1694700623
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_295
timestamp 1694700623
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_296
timestamp 1694700623
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_297
timestamp 1694700623
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_298
timestamp 1694700623
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_299
timestamp 1694700623
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_300
timestamp 1694700623
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_301
timestamp 1694700623
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_302
timestamp 1694700623
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_303
timestamp 1694700623
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_304
timestamp 1694700623
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_305
timestamp 1694700623
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_306
timestamp 1694700623
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_307
timestamp 1694700623
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_308
timestamp 1694700623
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_309
timestamp 1694700623
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_310
timestamp 1694700623
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_311
timestamp 1694700623
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_312
timestamp 1694700623
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_313
timestamp 1694700623
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_314
timestamp 1694700623
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_315
timestamp 1694700623
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_316
timestamp 1694700623
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_317
timestamp 1694700623
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_318
timestamp 1694700623
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_319
timestamp 1694700623
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_320
timestamp 1694700623
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_321
timestamp 1694700623
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_322
timestamp 1694700623
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_323
timestamp 1694700623
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_324
timestamp 1694700623
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_325
timestamp 1694700623
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_326
timestamp 1694700623
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_327
timestamp 1694700623
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_328
timestamp 1694700623
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_329
timestamp 1694700623
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_330
timestamp 1694700623
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_331
timestamp 1694700623
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_332
timestamp 1694700623
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_333
timestamp 1694700623
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_334
timestamp 1694700623
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_335
timestamp 1694700623
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_336
timestamp 1694700623
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_337
timestamp 1694700623
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_338
timestamp 1694700623
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_339
timestamp 1694700623
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_340
timestamp 1694700623
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_341
timestamp 1694700623
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_342
timestamp 1694700623
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_343
timestamp 1694700623
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_344
timestamp 1694700623
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_345
timestamp 1694700623
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_346
timestamp 1694700623
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_347
timestamp 1694700623
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_348
timestamp 1694700623
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_349
timestamp 1694700623
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_350
timestamp 1694700623
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_351
timestamp 1694700623
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_352
timestamp 1694700623
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_353
timestamp 1694700623
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_354
timestamp 1694700623
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_355
timestamp 1694700623
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_356
timestamp 1694700623
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_357
timestamp 1694700623
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_358
timestamp 1694700623
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_359
timestamp 1694700623
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_360
timestamp 1694700623
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_361
timestamp 1694700623
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_362
timestamp 1694700623
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_363
timestamp 1694700623
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_364
timestamp 1694700623
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_365
timestamp 1694700623
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_366
timestamp 1694700623
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_367
timestamp 1694700623
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_368
timestamp 1694700623
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_369
timestamp 1694700623
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_370
timestamp 1694700623
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_371
timestamp 1694700623
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_372
timestamp 1694700623
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_373
timestamp 1694700623
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_374
timestamp 1694700623
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_375
timestamp 1694700623
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_376
timestamp 1694700623
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_377
timestamp 1694700623
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_378
timestamp 1694700623
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_379
timestamp 1694700623
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_380
timestamp 1694700623
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_381
timestamp 1694700623
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_382
timestamp 1694700623
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_383
timestamp 1694700623
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_384
timestamp 1694700623
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_385
timestamp 1694700623
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_386
timestamp 1694700623
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_387
timestamp 1694700623
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_388
timestamp 1694700623
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_389
timestamp 1694700623
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_390
timestamp 1694700623
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_391
timestamp 1694700623
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_392
timestamp 1694700623
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_393
timestamp 1694700623
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_394
timestamp 1694700623
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_395
timestamp 1694700623
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_396
timestamp 1694700623
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_397
timestamp 1694700623
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_398
timestamp 1694700623
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_399
timestamp 1694700623
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_400
timestamp 1694700623
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_401
timestamp 1694700623
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_402
timestamp 1694700623
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_403
timestamp 1694700623
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_404
timestamp 1694700623
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_405
timestamp 1694700623
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_406
timestamp 1694700623
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_407
timestamp 1694700623
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_408
timestamp 1694700623
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_409
timestamp 1694700623
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_410
timestamp 1694700623
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_411
timestamp 1694700623
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_412
timestamp 1694700623
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_413
timestamp 1694700623
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_414
timestamp 1694700623
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_415
timestamp 1694700623
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[0\].cap
timestamp 1694700623
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[0\].cap_49 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[1\].cap
timestamp 1694700623
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[1\].cap_56
timestamp 1694700623
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[2\].cap
timestamp 1694700623
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[2\].cap_57
timestamp 1694700623
transform -1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[3\].cap_58
timestamp 1694700623
transform -1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[3\].cap
timestamp 1694700623
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[4\].cap_59
timestamp 1694700623
transform -1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[4\].cap
timestamp 1694700623
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[5\].cap
timestamp 1694700623
transform -1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[5\].cap_60
timestamp 1694700623
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[6\].cap_61
timestamp 1694700623
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[6\].cap
timestamp 1694700623
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[7\].cap_62
timestamp 1694700623
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[7\].cap
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[8\].cap
timestamp 1694700623
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[8\].cap_63
timestamp 1694700623
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[9\].cap_64
timestamp 1694700623
transform -1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[9\].cap
timestamp 1694700623
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[10\].cap_50
timestamp 1694700623
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[10\].cap
timestamp 1694700623
transform 1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[11\].cap_51
timestamp 1694700623
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[11\].cap
timestamp 1694700623
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[12\].cap
timestamp 1694700623
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[12\].cap_52
timestamp 1694700623
transform -1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[13\].cap_53
timestamp 1694700623
transform -1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[13\].cap
timestamp 1694700623
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[14\].cap
timestamp 1694700623
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[14\].cap_54
timestamp 1694700623
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[15\].cap_55
timestamp 1694700623
transform -1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[15\].cap
timestamp 1694700623
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2852 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1694700623
transform 1 0 2852 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1694700623
transform 1 0 1748 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1694700623
transform 1 0 2300 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1694700623
transform 1 0 1380 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1694700623
transform -1 0 2300 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1694700623
transform 1 0 1840 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1694700623
transform -1 0 2852 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1694700623
transform 1 0 2300 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1694700623
transform 1 0 2852 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1694700623
transform 1 0 1380 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1694700623
transform -1 0 2392 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1694700623
transform -1 0 2300 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1694700623
transform 1 0 2392 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1694700623
transform 1 0 4324 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1694700623
transform 1 0 5980 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1694700623
transform 1 0 4784 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1694700623
transform 1 0 5520 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1694700623
transform 1 0 3864 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1694700623
transform 1 0 6440 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1694700623
transform 1 0 4784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1694700623
transform 1 0 6348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1694700623
transform 1 0 3864 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1694700623
transform -1 0 6808 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1694700623
transform 1 0 3864 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1694700623
transform 1 0 5060 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1694700623
transform -1 0 4784 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1694700623
transform 1 0 6808 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1694700623
transform -1 0 4784 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1694700623
transform 1 0 5796 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1694700623
transform 1 0 10948 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1694700623
transform 1 0 10212 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1694700623
transform 1 0 9660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1694700623
transform 1 0 7176 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1694700623
transform 1 0 11592 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1694700623
transform 1 0 7360 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1694700623
transform -1 0 11132 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1694700623
transform 1 0 9752 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1694700623
transform -1 0 11500 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1694700623
transform -1 0 8648 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1694700623
transform 1 0 10212 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1694700623
transform -1 0 8188 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1694700623
transform 1 0 11500 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1694700623
transform 1 0 9292 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1694700623
transform 1 0 9568 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1694700623
transform 1 0 9752 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1694700623
transform 1 0 11592 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1694700623
transform 1 0 9292 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1694700623
transform -1 0 12512 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1694700623
transform -1 0 8832 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1694700623
transform 1 0 10028 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1694700623
transform -1 0 9660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1694700623
transform 1 0 9108 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1694700623
transform -1 0 7360 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1694700623
transform -1 0 12972 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1694700623
transform -1 0 9752 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1694700623
transform 1 0 10488 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1694700623
transform 1 0 7820 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1694700623
transform -1 0 11592 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1694700623
transform 1 0 7636 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1694700623
transform -1 0 11040 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1694700623
transform 1 0 8096 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd_66
timestamp 1694700623
transform 1 0 4508 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1694700623
transform 1 0 3220 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].vref_65
timestamp 1694700623
transform 1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].vref
timestamp 1694700623
transform -1 0 11224 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dcdc
timestamp 1694700623
transform -1 0 3956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  temp1.inv1_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_2
timestamp 1694700623
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_3
timestamp 1694700623
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_4
timestamp 1694700623
transform -1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2
timestamp 1694700623
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire1
timestamp 1694700623
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire12
timestamp 1694700623
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire15
timestamp 1694700623
transform -1 0 14904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire16
timestamp 1694700623
transform -1 0 14168 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire19
timestamp 1694700623
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
<< labels >>
flabel metal3 s 29600 3000 30000 3120 0 FreeSans 480 0 0 0 dbg_delay
port 0 nsew signal tristate
flabel metal3 s 29600 7624 30000 7744 0 FreeSans 480 0 0 0 dbg_result[0]
port 1 nsew signal tristate
flabel metal3 s 29600 12248 30000 12368 0 FreeSans 480 0 0 0 dbg_result[1]
port 2 nsew signal tristate
flabel metal3 s 29600 16872 30000 16992 0 FreeSans 480 0 0 0 dbg_result[2]
port 3 nsew signal tristate
flabel metal3 s 29600 21496 30000 21616 0 FreeSans 480 0 0 0 dbg_result[3]
port 4 nsew signal tristate
flabel metal3 s 29600 26120 30000 26240 0 FreeSans 480 0 0 0 dbg_result[4]
port 5 nsew signal tristate
flabel metal3 s 29600 30744 30000 30864 0 FreeSans 480 0 0 0 dbg_result[5]
port 6 nsew signal tristate
flabel metal3 s 0 2456 400 2576 0 FreeSans 480 0 0 0 io_in[0]
port 7 nsew signal input
flabel metal3 s 0 4360 400 4480 0 FreeSans 480 0 0 0 io_in[1]
port 8 nsew signal input
flabel metal3 s 0 6264 400 6384 0 FreeSans 480 0 0 0 io_in[2]
port 9 nsew signal input
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 io_in[3]
port 10 nsew signal input
flabel metal3 s 0 10072 400 10192 0 FreeSans 480 0 0 0 io_in[4]
port 11 nsew signal input
flabel metal3 s 0 11976 400 12096 0 FreeSans 480 0 0 0 io_in[5]
port 12 nsew signal input
flabel metal3 s 0 13880 400 14000 0 FreeSans 480 0 0 0 io_in[6]
port 13 nsew signal input
flabel metal3 s 0 15784 400 15904 0 FreeSans 480 0 0 0 io_in[7]
port 14 nsew signal input
flabel metal3 s 0 17688 400 17808 0 FreeSans 480 0 0 0 io_out[0]
port 15 nsew signal tristate
flabel metal3 s 0 19592 400 19712 0 FreeSans 480 0 0 0 io_out[1]
port 16 nsew signal tristate
flabel metal3 s 0 21496 400 21616 0 FreeSans 480 0 0 0 io_out[2]
port 17 nsew signal tristate
flabel metal3 s 0 23400 400 23520 0 FreeSans 480 0 0 0 io_out[3]
port 18 nsew signal tristate
flabel metal3 s 0 25304 400 25424 0 FreeSans 480 0 0 0 io_out[4]
port 19 nsew signal tristate
flabel metal3 s 0 27208 400 27328 0 FreeSans 480 0 0 0 io_out[5]
port 20 nsew signal tristate
flabel metal3 s 0 29112 400 29232 0 FreeSans 480 0 0 0 io_out[6]
port 21 nsew signal tristate
flabel metal3 s 0 31016 400 31136 0 FreeSans 480 0 0 0 io_out[7]
port 22 nsew signal tristate
flabel metal4 s 4417 1040 4737 32688 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 11363 1040 11683 32688 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 18309 1040 18629 32688 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 25255 1040 25575 32688 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 7890 1040 8210 32688 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 14836 1040 15156 32688 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 21782 1040 22102 32688 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
flabel metal4 s 28728 1040 29048 32688 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
rlabel metal1 14996 32096 14996 32096 0 vccd1
rlabel via1 15076 32640 15076 32640 0 vssd1
rlabel metal1 2990 9928 2990 9928 0 _0000_
rlabel metal1 7636 16218 7636 16218 0 _0001_
rlabel metal1 8459 16150 8459 16150 0 _0002_
rlabel metal1 9844 15674 9844 15674 0 _0003_
rlabel metal2 11178 15266 11178 15266 0 _0004_
rlabel metal2 12190 17442 12190 17442 0 _0005_
rlabel metal2 12006 26758 12006 26758 0 _0006_
rlabel via1 12645 27438 12645 27438 0 _0007_
rlabel via1 12829 25262 12829 25262 0 _0008_
rlabel metal1 13565 23766 13565 23766 0 _0009_
rlabel metal2 15042 13702 15042 13702 0 _0010_
rlabel metal1 18522 13974 18522 13974 0 _0011_
rlabel metal1 20884 14042 20884 14042 0 _0012_
rlabel via1 22397 13226 22397 13226 0 _0013_
rlabel metal1 24338 12818 24338 12818 0 _0014_
rlabel metal1 25258 13294 25258 13294 0 _0015_
rlabel metal1 15210 12886 15210 12886 0 _0016_
rlabel metal1 17970 12886 17970 12886 0 _0017_
rlabel via1 6660 12886 6660 12886 0 _0018_
rlabel metal1 7774 12682 7774 12682 0 _0019_
rlabel metal2 9798 13090 9798 13090 0 _0020_
rlabel metal2 12558 13668 12558 13668 0 _0021_
rlabel metal1 16560 14586 16560 14586 0 _0022_
rlabel metal1 19166 15402 19166 15402 0 _0023_
rlabel metal1 21466 16490 21466 16490 0 _0024_
rlabel metal1 24292 17238 24292 17238 0 _0025_
rlabel metal1 23547 19414 23547 19414 0 _0026_
rlabel metal2 25438 19618 25438 19618 0 _0027_
rlabel metal2 18814 16966 18814 16966 0 _0028_
rlabel via1 20276 17170 20276 17170 0 _0029_
rlabel metal2 21482 21522 21482 21522 0 _0030_
rlabel metal2 23966 22882 23966 22882 0 _0031_
rlabel metal1 24794 21896 24794 21896 0 _0032_
rlabel metal1 26362 20502 26362 20502 0 _0033_
rlabel metal1 15118 19754 15118 19754 0 _0034_
rlabel metal1 14071 16150 14071 16150 0 _0035_
rlabel via1 7401 14382 7401 14382 0 _0036_
rlabel via1 7677 11118 7677 11118 0 _0037_
rlabel metal1 9782 11798 9782 11798 0 _0038_
rlabel metal1 13294 21114 13294 21114 0 _0039_
rlabel metal2 14674 21726 14674 21726 0 _0040_
rlabel metal2 16698 21794 16698 21794 0 _0041_
rlabel metal2 16606 26962 16606 26962 0 _0042_
rlabel metal1 17618 28662 17618 28662 0 _0043_
rlabel metal1 15451 29206 15451 29206 0 _0044_
rlabel via1 15681 25262 15681 25262 0 _0045_
rlabel metal2 17802 25058 17802 25058 0 _0046_
rlabel metal1 18890 25942 18890 25942 0 _0047_
rlabel metal2 19734 28662 19734 28662 0 _0048_
rlabel metal1 13616 28730 13616 28730 0 _0049_
rlabel metal1 14858 28730 14858 28730 0 _0050_
rlabel metal1 17848 28730 17848 28730 0 _0051_
rlabel metal2 19734 26758 19734 26758 0 _0052_
rlabel metal2 20746 27880 20746 27880 0 _0053_
rlabel metal2 21666 28288 21666 28288 0 _0054_
rlabel metal1 23613 27370 23613 27370 0 _0055_
rlabel metal1 23782 26554 23782 26554 0 _0056_
rlabel metal1 24154 20502 24154 20502 0 _0057_
rlabel via1 22958 19822 22958 19822 0 _0058_
rlabel via1 20649 19754 20649 19754 0 _0059_
rlabel metal1 21781 23834 21781 23834 0 _0060_
rlabel metal1 24272 24106 24272 24106 0 _0061_
rlabel metal1 25054 23766 25054 23766 0 _0062_
rlabel metal1 26082 21658 26082 21658 0 _0063_
rlabel metal1 20071 22712 20071 22712 0 _0064_
rlabel metal2 20654 21726 20654 21726 0 _0065_
rlabel metal2 21666 15198 21666 15198 0 _0066_
rlabel metal1 23828 14586 23828 14586 0 _0067_
rlabel metal2 24794 15878 24794 15878 0 _0068_
rlabel metal2 25530 17442 25530 17442 0 _0069_
rlabel metal1 26756 18326 26756 18326 0 _0070_
rlabel metal1 27503 16150 27503 16150 0 _0071_
rlabel metal2 26450 16354 26450 16354 0 _0072_
rlabel metal2 27462 17442 27462 17442 0 _0073_
rlabel metal1 24686 18326 24686 18326 0 _0074_
rlabel via1 26261 18734 26261 18734 0 _0075_
rlabel via1 17148 18326 17148 18326 0 _0076_
rlabel metal1 18128 16082 18128 16082 0 _0077_
rlabel viali 8413 15062 8413 15062 0 _0078_
rlabel via1 9241 14382 9241 14382 0 _0079_
rlabel via1 10897 14382 10897 14382 0 _0080_
rlabel metal2 12926 22882 12926 22882 0 _0081_
rlabel metal1 17572 23834 17572 23834 0 _0082_
rlabel metal1 19356 24786 19356 24786 0 _0083_
rlabel metal2 21298 25058 21298 25058 0 _0084_
rlabel metal2 22494 25058 22494 25058 0 _0085_
rlabel metal1 24150 24922 24150 24922 0 _0086_
rlabel metal2 21482 26146 21482 26146 0 _0087_
rlabel metal1 17700 26350 17700 26350 0 _0088_
rlabel metal2 19182 28322 19182 28322 0 _0089_
rlabel metal1 18358 28118 18358 28118 0 _0090_
rlabel metal1 15083 28118 15083 28118 0 _0091_
rlabel metal1 13646 27030 13646 27030 0 _0092_
rlabel metal1 14485 24854 14485 24854 0 _0093_
rlabel metal1 15129 23766 15129 23766 0 _0094_
rlabel metal2 15410 17442 15410 17442 0 _0095_
rlabel metal1 12645 14382 12645 14382 0 _0096_
rlabel metal1 13206 11118 13206 11118 0 _0097_
rlabel metal2 12466 9418 12466 9418 0 _0098_
rlabel metal2 12926 9350 12926 9350 0 _0099_
rlabel metal1 14658 10710 14658 10710 0 _0100_
rlabel metal2 16238 10914 16238 10914 0 _0101_
rlabel metal1 19448 11118 19448 11118 0 _0102_
rlabel metal1 20920 11118 20920 11118 0 _0103_
rlabel metal2 21206 9826 21206 9826 0 _0104_
rlabel metal2 18998 9350 18998 9350 0 _0105_
rlabel metal1 17015 9622 17015 9622 0 _0106_
rlabel metal1 19136 9078 19136 9078 0 _0107_
rlabel viali 22121 8466 22121 8466 0 _0108_
rlabel metal2 23322 7650 23322 7650 0 _0109_
rlabel via1 20005 7854 20005 7854 0 _0110_
rlabel metal2 18722 7650 18722 7650 0 _0111_
rlabel metal1 17751 6698 17751 6698 0 _0112_
rlabel metal1 19448 5678 19448 5678 0 _0113_
rlabel metal1 20976 4250 20976 4250 0 _0114_
rlabel metal1 23133 4114 23133 4114 0 _0115_
rlabel metal2 23874 3910 23874 3910 0 _0116_
rlabel metal2 19734 4386 19734 4386 0 _0117_
rlabel metal1 13841 5270 13841 5270 0 _0118_
rlabel metal2 14766 5474 14766 5474 0 _0119_
rlabel metal1 7815 8942 7815 8942 0 _0120_
rlabel metal1 8924 8058 8924 8058 0 _0121_
rlabel metal1 10304 6970 10304 6970 0 _0122_
rlabel metal1 11720 7378 11720 7378 0 _0123_
rlabel metal1 13386 6664 13386 6664 0 _0124_
rlabel metal1 14566 7446 14566 7446 0 _0125_
rlabel metal1 8045 6766 8045 6766 0 _0126_
rlabel metal1 9138 6358 9138 6358 0 _0127_
rlabel metal1 10702 5610 10702 5610 0 _0128_
rlabel via1 11725 3502 11725 3502 0 _0129_
rlabel metal2 12926 3910 12926 3910 0 _0130_
rlabel metal1 14025 4182 14025 4182 0 _0131_
rlabel metal1 8050 3706 8050 3706 0 _0132_
rlabel via1 6573 3502 6573 3502 0 _0133_
rlabel metal1 5377 4114 5377 4114 0 _0134_
rlabel metal2 7038 5474 7038 5474 0 _0135_
rlabel metal1 4354 5610 4354 5610 0 _0136_
rlabel metal1 4814 6358 4814 6358 0 _0137_
rlabel metal1 5469 9622 5469 9622 0 _0138_
rlabel metal1 6389 8942 6389 8942 0 _0139_
rlabel metal1 3894 8874 3894 8874 0 _0140_
rlabel metal1 4794 7378 4794 7378 0 _0141_
rlabel metal2 4922 7650 4922 7650 0 _0142_
rlabel metal1 6711 7446 6711 7446 0 _0143_
rlabel metal1 6792 6358 6792 6358 0 _0144_
rlabel metal1 7942 5270 7942 5270 0 _0145_
rlabel metal1 10212 3162 10212 3162 0 _0146_
rlabel metal1 12082 2346 12082 2346 0 _0147_
rlabel via1 14393 1326 14393 1326 0 _0148_
rlabel metal2 16514 2210 16514 2210 0 _0149_
rlabel metal2 19642 1734 19642 1734 0 _0150_
rlabel metal1 21880 2006 21880 2006 0 _0151_
rlabel metal1 23234 3094 23234 3094 0 _0152_
rlabel metal1 20920 2414 20920 2414 0 _0153_
rlabel metal2 19642 2210 19642 2210 0 _0154_
rlabel metal1 17786 3434 17786 3434 0 _0155_
rlabel metal1 20178 3434 20178 3434 0 _0156_
rlabel metal1 21758 6426 21758 6426 0 _0157_
rlabel metal1 22478 6358 22478 6358 0 _0158_
rlabel metal1 25028 5678 25028 5678 0 _0159_
rlabel via1 26086 5270 26086 5270 0 _0160_
rlabel metal2 26174 6562 26174 6562 0 _0161_
rlabel metal1 27124 7446 27124 7446 0 _0162_
rlabel metal1 24564 6970 24564 6970 0 _0163_
rlabel metal1 24456 8874 24456 8874 0 _0164_
rlabel metal1 25514 8534 25514 8534 0 _0165_
rlabel metal1 26986 8874 26986 8874 0 _0166_
rlabel metal2 27462 15266 27462 15266 0 _0167_
rlabel metal1 26592 14382 26592 14382 0 _0168_
rlabel via1 25893 10030 25893 10030 0 _0169_
rlabel metal2 27554 9826 27554 9826 0 _0170_
rlabel metal2 27462 11526 27462 11526 0 _0171_
rlabel via1 27457 12818 27457 12818 0 _0172_
rlabel metal1 28198 13498 28198 13498 0 _0173_
rlabel metal2 26266 13090 26266 13090 0 _0174_
rlabel metal1 25856 12138 25856 12138 0 _0175_
rlabel metal1 25764 11118 25764 11118 0 _0176_
rlabel metal1 17484 4182 17484 4182 0 _0177_
rlabel metal1 15451 4182 15451 4182 0 _0178_
rlabel metal1 15267 3026 15267 3026 0 _0179_
rlabel metal1 8367 2006 8367 2006 0 _0180_
rlabel metal1 9379 1326 9379 1326 0 _0181_
rlabel via1 10253 2006 10253 2006 0 _0182_
rlabel metal2 12190 1734 12190 1734 0 _0183_
rlabel metal1 14796 2006 14796 2006 0 _0184_
rlabel metal2 17434 1734 17434 1734 0 _0185_
rlabel metal2 7222 2210 7222 2210 0 _0186_
rlabel metal1 7079 10710 7079 10710 0 _0187_
rlabel metal1 5857 10710 5857 10710 0 _0188_
rlabel via1 5745 11118 5745 11118 0 _0189_
rlabel metal1 6470 12138 6470 12138 0 _0190_
rlabel metal1 13192 12818 13192 12818 0 _0191_
rlabel metal1 6394 14994 6394 14994 0 _0192_
rlabel metal1 5612 16490 5612 16490 0 _0193_
rlabel metal1 7176 18802 7176 18802 0 _0194_
rlabel metal1 6394 18258 6394 18258 0 _0195_
rlabel metal2 10718 27268 10718 27268 0 _0196_
rlabel metal1 10350 28186 10350 28186 0 _0197_
rlabel metal1 3634 15674 3634 15674 0 _0198_
rlabel via1 1697 15062 1697 15062 0 _0199_
rlabel via1 1697 12818 1697 12818 0 _0200_
rlabel metal1 4052 10710 4052 10710 0 _0201_
rlabel metal1 2594 14314 2594 14314 0 _0202_
rlabel metal1 3802 12886 3802 12886 0 _0203_
rlabel metal1 4814 13226 4814 13226 0 _0204_
rlabel metal1 4912 14994 4912 14994 0 _0205_
rlabel metal1 6808 26554 6808 26554 0 _0206_
rlabel metal1 4876 27574 4876 27574 0 _0207_
rlabel metal2 5106 29410 5106 29410 0 _0208_
rlabel metal2 6394 29138 6394 29138 0 _0209_
rlabel metal1 7728 28730 7728 28730 0 _0210_
rlabel metal1 9430 28730 9430 28730 0 _0211_
rlabel via1 7217 27370 7217 27370 0 _0212_
rlabel metal1 14858 21114 14858 21114 0 _0213_
rlabel metal1 16652 21522 16652 21522 0 _0214_
rlabel metal1 17250 24786 17250 24786 0 _0215_
rlabel metal1 13662 21896 13662 21896 0 _0216_
rlabel metal1 17158 28526 17158 28526 0 _0217_
rlabel metal1 16008 29818 16008 29818 0 _0218_
rlabel metal2 15778 26180 15778 26180 0 _0219_
rlabel metal1 17986 24854 17986 24854 0 _0220_
rlabel metal1 19090 25466 19090 25466 0 _0221_
rlabel metal1 21068 15878 21068 15878 0 _0222_
rlabel metal1 19964 27642 19964 27642 0 _0223_
rlabel metal1 13984 28526 13984 28526 0 _0224_
rlabel metal1 14720 28526 14720 28526 0 _0225_
rlabel metal1 17434 28560 17434 28560 0 _0226_
rlabel metal1 19274 26350 19274 26350 0 _0227_
rlabel metal1 20792 27438 20792 27438 0 _0228_
rlabel metal2 21482 28084 21482 28084 0 _0229_
rlabel metal1 23966 27472 23966 27472 0 _0230_
rlabel metal1 23230 26350 23230 26350 0 _0231_
rlabel metal1 23644 20910 23644 20910 0 _0232_
rlabel metal1 22678 20400 22678 20400 0 _0233_
rlabel metal1 20148 20026 20148 20026 0 _0234_
rlabel metal1 21390 23290 21390 23290 0 _0235_
rlabel metal1 23690 24208 23690 24208 0 _0236_
rlabel metal1 16836 19278 16836 19278 0 _0237_
rlabel metal1 24748 23698 24748 23698 0 _0238_
rlabel metal2 25806 21801 25806 21801 0 _0239_
rlabel metal1 19688 21930 19688 21930 0 _0240_
rlabel metal1 20700 21998 20700 21998 0 _0241_
rlabel metal1 21666 15470 21666 15470 0 _0242_
rlabel metal1 23690 14416 23690 14416 0 _0243_
rlabel metal2 24978 15300 24978 15300 0 _0244_
rlabel metal1 25484 16762 25484 16762 0 _0245_
rlabel metal1 19642 16048 19642 16048 0 _0246_
rlabel metal1 26220 18258 26220 18258 0 _0247_
rlabel metal1 27232 16558 27232 16558 0 _0248_
rlabel metal1 26496 16082 26496 16082 0 _0249_
rlabel metal1 27508 17170 27508 17170 0 _0250_
rlabel metal1 24380 17850 24380 17850 0 _0251_
rlabel metal2 25898 19142 25898 19142 0 _0252_
rlabel metal1 17388 18734 17388 18734 0 _0253_
rlabel metal1 18446 16592 18446 16592 0 _0254_
rlabel metal1 11086 15436 11086 15436 0 _0255_
rlabel metal1 9522 15130 9522 15130 0 _0256_
rlabel metal1 10580 14042 10580 14042 0 _0257_
rlabel via2 12466 15147 12466 15147 0 _0258_
rlabel metal1 17342 23664 17342 23664 0 _0259_
rlabel metal1 15824 18258 15824 18258 0 _0260_
rlabel metal1 19136 24378 19136 24378 0 _0261_
rlabel metal1 21482 24752 21482 24752 0 _0262_
rlabel metal1 22264 24786 22264 24786 0 _0263_
rlabel metal1 23736 24786 23736 24786 0 _0264_
rlabel metal1 21298 25840 21298 25840 0 _0265_
rlabel metal1 12742 21318 12742 21318 0 _0266_
rlabel metal1 17342 26010 17342 26010 0 _0267_
rlabel metal1 18952 27642 18952 27642 0 _0268_
rlabel metal2 18170 28084 18170 28084 0 _0269_
rlabel metal2 15410 27812 15410 27812 0 _0270_
rlabel metal1 13616 26962 13616 26962 0 _0271_
rlabel metal1 14720 25262 14720 25262 0 _0272_
rlabel metal1 15318 24174 15318 24174 0 _0273_
rlabel metal1 15410 17170 15410 17170 0 _0274_
rlabel metal1 12972 14994 12972 14994 0 _0275_
rlabel metal1 12880 10778 12880 10778 0 _0276_
rlabel metal1 12236 10030 12236 10030 0 _0277_
rlabel metal1 12742 8976 12742 8976 0 _0278_
rlabel metal1 14490 10234 14490 10234 0 _0279_
rlabel metal1 15962 10642 15962 10642 0 _0280_
rlabel metal2 18354 10948 18354 10948 0 _0281_
rlabel metal1 20286 10778 20286 10778 0 _0282_
rlabel metal1 20930 10744 20930 10744 0 _0283_
rlabel metal1 21344 9554 21344 9554 0 _0284_
rlabel metal1 19044 8942 19044 8942 0 _0285_
rlabel metal1 16698 9622 16698 9622 0 _0286_
rlabel metal1 18538 8976 18538 8976 0 _0287_
rlabel metal1 21206 8942 21206 8942 0 _0288_
rlabel metal1 23828 7378 23828 7378 0 _0289_
rlabel metal1 18538 6290 18538 6290 0 _0290_
rlabel metal1 19872 7514 19872 7514 0 _0291_
rlabel metal1 19872 7378 19872 7378 0 _0292_
rlabel metal1 18262 7344 18262 7344 0 _0293_
rlabel metal1 18860 6290 18860 6290 0 _0294_
rlabel metal1 20792 4114 20792 4114 0 _0295_
rlabel metal1 23966 4624 23966 4624 0 _0296_
rlabel metal2 23690 3978 23690 3978 0 _0297_
rlabel metal1 19780 4114 19780 4114 0 _0298_
rlabel metal1 12742 6290 12742 6290 0 _0299_
rlabel metal1 14306 5712 14306 5712 0 _0300_
rlabel metal1 14812 5202 14812 5202 0 _0301_
rlabel metal1 7912 8602 7912 8602 0 _0302_
rlabel metal1 8832 7854 8832 7854 0 _0303_
rlabel metal2 10534 7242 10534 7242 0 _0304_
rlabel metal1 11684 6970 11684 6970 0 _0305_
rlabel metal1 13570 6766 13570 6766 0 _0306_
rlabel metal1 14352 6970 14352 6970 0 _0307_
rlabel metal1 8464 7378 8464 7378 0 _0308_
rlabel metal1 9246 6290 9246 6290 0 _0309_
rlabel metal1 10488 5338 10488 5338 0 _0310_
rlabel metal1 11960 4590 11960 4590 0 _0311_
rlabel metal1 12972 3502 12972 3502 0 _0312_
rlabel metal1 14214 3706 14214 3706 0 _0313_
rlabel metal1 8326 3604 8326 3604 0 _0314_
rlabel metal1 6946 4182 6946 4182 0 _0315_
rlabel metal2 10166 4318 10166 4318 0 _0316_
rlabel metal1 5796 3706 5796 3706 0 _0317_
rlabel metal1 7222 5168 7222 5168 0 _0318_
rlabel metal1 5290 5304 5290 5304 0 _0319_
rlabel metal1 4784 5338 4784 5338 0 _0320_
rlabel metal2 5750 9588 5750 9588 0 _0321_
rlabel metal1 6808 8602 6808 8602 0 _0322_
rlabel metal1 3128 8942 3128 8942 0 _0323_
rlabel metal1 5796 8466 5796 8466 0 _0324_
rlabel metal1 5106 7412 5106 7412 0 _0325_
rlabel metal1 6532 7854 6532 7854 0 _0326_
rlabel metal1 6394 6800 6394 6800 0 _0327_
rlabel metal1 7636 5202 7636 5202 0 _0328_
rlabel metal1 10166 3026 10166 3026 0 _0329_
rlabel metal2 22310 1870 22310 1870 0 _0330_
rlabel metal2 11776 2652 11776 2652 0 _0331_
rlabel metal1 14030 2414 14030 2414 0 _0332_
rlabel metal1 16629 1870 16629 1870 0 _0333_
rlabel metal1 19366 1326 19366 1326 0 _0334_
rlabel metal1 21666 1530 21666 1530 0 _0335_
rlabel metal1 22724 2618 22724 2618 0 _0336_
rlabel metal1 21022 2992 21022 2992 0 _0337_
rlabel metal1 19504 1938 19504 1938 0 _0338_
rlabel metal1 17572 3162 17572 3162 0 _0339_
rlabel metal1 19780 3502 19780 3502 0 _0340_
rlabel metal1 21390 6664 21390 6664 0 _0341_
rlabel metal1 22034 6324 22034 6324 0 _0342_
rlabel metal1 22632 6970 22632 6970 0 _0343_
rlabel metal1 24334 6256 24334 6256 0 _0344_
rlabel metal1 25898 5780 25898 5780 0 _0345_
rlabel metal1 26220 6290 26220 6290 0 _0346_
rlabel metal2 26818 7684 26818 7684 0 _0347_
rlabel metal2 24886 7140 24886 7140 0 _0348_
rlabel metal1 24242 8602 24242 8602 0 _0349_
rlabel metal1 25530 8466 25530 8466 0 _0350_
rlabel metal1 26818 8602 26818 8602 0 _0351_
rlabel metal1 25714 12920 25714 12920 0 _0352_
rlabel metal1 27462 14586 27462 14586 0 _0353_
rlabel metal1 26174 14960 26174 14960 0 _0354_
rlabel metal1 26082 10608 26082 10608 0 _0355_
rlabel metal1 27738 9520 27738 9520 0 _0356_
rlabel metal2 27462 10948 27462 10948 0 _0357_
rlabel metal2 27370 11764 27370 11764 0 _0358_
rlabel metal1 27922 13328 27922 13328 0 _0359_
rlabel metal1 26128 12818 26128 12818 0 _0360_
rlabel metal2 25208 12614 25208 12614 0 _0361_
rlabel metal1 25392 11730 25392 11730 0 _0362_
rlabel metal1 12466 1972 12466 1972 0 _0363_
rlabel metal1 17112 3706 17112 3706 0 _0364_
rlabel metal1 15732 3706 15732 3706 0 _0365_
rlabel metal1 15732 2414 15732 2414 0 _0366_
rlabel metal1 9016 3026 9016 3026 0 _0367_
rlabel metal1 9568 2414 9568 2414 0 _0368_
rlabel metal1 9982 2074 9982 2074 0 _0369_
rlabel metal2 12006 1530 12006 1530 0 _0370_
rlabel metal1 14398 1904 14398 1904 0 _0371_
rlabel metal1 17204 1326 17204 1326 0 _0372_
rlabel metal1 7406 2006 7406 2006 0 _0373_
rlabel metal1 7452 10234 7452 10234 0 _0374_
rlabel metal1 5980 10234 5980 10234 0 _0375_
rlabel metal1 5520 11322 5520 11322 0 _0376_
rlabel metal1 6256 11866 6256 11866 0 _0377_
rlabel metal1 12834 12240 12834 12240 0 _0378_
rlabel metal1 3266 16218 3266 16218 0 _0379_
rlabel metal2 3082 17391 3082 17391 0 _0380_
rlabel metal2 5934 16558 5934 16558 0 _0381_
rlabel metal1 5382 16694 5382 16694 0 _0382_
rlabel metal1 6946 18734 6946 18734 0 _0383_
rlabel metal1 5520 17782 5520 17782 0 _0384_
rlabel metal1 10626 26928 10626 26928 0 _0385_
rlabel metal2 9982 27302 9982 27302 0 _0386_
rlabel metal1 4370 15572 4370 15572 0 _0387_
rlabel metal1 1840 15470 1840 15470 0 _0388_
rlabel metal1 2484 12206 2484 12206 0 _0389_
rlabel metal1 2070 12308 2070 12308 0 _0390_
rlabel metal2 2530 11424 2530 11424 0 _0391_
rlabel metal1 3726 11118 3726 11118 0 _0392_
rlabel metal2 3542 14484 3542 14484 0 _0393_
rlabel metal1 3588 14586 3588 14586 0 _0394_
rlabel metal1 3910 12818 3910 12818 0 _0395_
rlabel metal1 3680 11866 3680 11866 0 _0396_
rlabel metal1 4462 13362 4462 13362 0 _0397_
rlabel metal1 4600 14586 4600 14586 0 _0398_
rlabel metal1 6486 26248 6486 26248 0 _0399_
rlabel metal2 6394 26554 6394 26554 0 _0400_
rlabel metal1 4922 27404 4922 27404 0 _0401_
rlabel metal1 5244 28730 5244 28730 0 _0402_
rlabel metal1 7084 28186 7084 28186 0 _0403_
rlabel metal1 6762 28526 6762 28526 0 _0404_
rlabel metal1 7774 28560 7774 28560 0 _0405_
rlabel metal1 8970 28492 8970 28492 0 _0406_
rlabel metal1 9154 28560 9154 28560 0 _0407_
rlabel metal2 6762 27948 6762 27948 0 _0408_
rlabel metal1 6072 26418 6072 26418 0 _0409_
rlabel metal1 1978 22984 1978 22984 0 _0410_
rlabel metal1 1978 22576 1978 22576 0 _0411_
rlabel metal1 1794 13498 1794 13498 0 _0412_
rlabel metal1 2346 21998 2346 21998 0 _0413_
rlabel metal1 2254 21318 2254 21318 0 _0414_
rlabel metal1 2254 23766 2254 23766 0 _0415_
rlabel metal1 1840 24786 1840 24786 0 _0416_
rlabel metal1 2116 23086 2116 23086 0 _0417_
rlabel metal1 3818 16116 3818 16116 0 _0418_
rlabel metal1 3358 21046 3358 21046 0 _0419_
rlabel metal1 2254 18802 2254 18802 0 _0420_
rlabel metal1 2622 18938 2622 18938 0 _0421_
rlabel metal2 1794 18836 1794 18836 0 _0422_
rlabel metal1 2714 19312 2714 19312 0 _0423_
rlabel metal1 4784 25874 4784 25874 0 _0424_
rlabel metal1 13846 20468 13846 20468 0 _0425_
rlabel metal1 3772 18666 3772 18666 0 _0426_
rlabel metal1 4232 20434 4232 20434 0 _0427_
rlabel metal2 2070 15980 2070 15980 0 _0428_
rlabel metal2 4646 19346 4646 19346 0 _0429_
rlabel metal1 4600 19210 4600 19210 0 _0430_
rlabel metal1 6486 19346 6486 19346 0 _0431_
rlabel metal1 5290 19856 5290 19856 0 _0432_
rlabel metal1 9982 17646 9982 17646 0 _0433_
rlabel metal1 7866 20434 7866 20434 0 _0434_
rlabel metal1 6624 20774 6624 20774 0 _0435_
rlabel metal1 6854 17578 6854 17578 0 _0436_
rlabel metal1 7866 19278 7866 19278 0 _0437_
rlabel metal2 13294 20502 13294 20502 0 _0438_
rlabel metal1 7590 19346 7590 19346 0 _0439_
rlabel metal2 14214 11968 14214 11968 0 _0440_
rlabel metal1 17802 5066 17802 5066 0 _0441_
rlabel metal2 14674 17816 14674 17816 0 _0442_
rlabel viali 20922 15062 20922 15062 0 _0443_
rlabel metal1 21160 6222 21160 6222 0 _0444_
rlabel metal1 17158 8874 17158 8874 0 _0445_
rlabel metal2 13018 20825 13018 20825 0 _0446_
rlabel metal1 13570 20366 13570 20366 0 _0447_
rlabel metal1 14490 20434 14490 20434 0 _0448_
rlabel metal1 22126 11696 22126 11696 0 _0449_
rlabel metal1 16146 8466 16146 8466 0 _0450_
rlabel metal2 13294 8959 13294 8959 0 _0451_
rlabel metal1 20792 18802 20792 18802 0 _0452_
rlabel metal2 18262 19618 18262 19618 0 _0453_
rlabel metal2 19642 17442 19642 17442 0 _0454_
rlabel metal1 16054 14994 16054 14994 0 _0455_
rlabel metal1 21114 13226 21114 13226 0 _0456_
rlabel metal1 20700 11730 20700 11730 0 _0457_
rlabel metal2 21758 11594 21758 11594 0 _0458_
rlabel metal1 20378 18632 20378 18632 0 _0459_
rlabel metal1 21252 22066 21252 22066 0 _0460_
rlabel metal1 18906 19822 18906 19822 0 _0461_
rlabel metal1 18852 18598 18852 18598 0 _0462_
rlabel metal1 22816 23120 22816 23120 0 _0463_
rlabel metal1 17158 18802 17158 18802 0 _0464_
rlabel metal1 22234 21590 22234 21590 0 _0465_
rlabel metal1 17342 23120 17342 23120 0 _0466_
rlabel metal2 16054 19584 16054 19584 0 _0467_
rlabel metal2 17986 20298 17986 20298 0 _0468_
rlabel metal2 23414 23154 23414 23154 0 _0469_
rlabel metal1 23506 23290 23506 23290 0 _0470_
rlabel metal1 22448 18054 22448 18054 0 _0471_
rlabel metal1 14168 18326 14168 18326 0 _0472_
rlabel metal2 23230 17476 23230 17476 0 _0473_
rlabel metal1 17745 19414 17745 19414 0 _0474_
rlabel metal1 18078 15504 18078 15504 0 _0475_
rlabel metal1 21114 5032 21114 5032 0 _0476_
rlabel metal1 17396 14314 17396 14314 0 _0477_
rlabel metal1 23322 4794 23322 4794 0 _0478_
rlabel metal3 23759 16660 23759 16660 0 _0479_
rlabel metal1 22678 17850 22678 17850 0 _0480_
rlabel metal1 13202 15674 13202 15674 0 _0481_
rlabel metal1 17066 24684 17066 24684 0 _0482_
rlabel metal1 15824 21998 15824 21998 0 _0483_
rlabel metal1 16008 21862 16008 21862 0 _0484_
rlabel metal1 14168 20910 14168 20910 0 _0485_
rlabel metal1 15272 23086 15272 23086 0 _0486_
rlabel metal1 16928 13906 16928 13906 0 _0487_
rlabel metal1 15410 27472 15410 27472 0 _0488_
rlabel metal3 18653 26316 18653 26316 0 _0489_
rlabel metal2 17434 18343 17434 18343 0 _0490_
rlabel metal1 15226 18054 15226 18054 0 _0491_
rlabel metal1 16330 17646 16330 17646 0 _0492_
rlabel metal1 13340 7854 13340 7854 0 _0493_
rlabel metal1 10488 9146 10488 9146 0 _0494_
rlabel metal1 15556 20774 15556 20774 0 _0495_
rlabel viali 9233 11118 9233 11118 0 _0496_
rlabel metal1 9890 11118 9890 11118 0 _0497_
rlabel metal1 16238 5780 16238 5780 0 _0498_
rlabel metal1 10212 5814 10212 5814 0 _0499_
rlabel metal2 17158 20332 17158 20332 0 _0500_
rlabel metal1 20562 13940 20562 13940 0 _0501_
rlabel metal1 14030 5678 14030 5678 0 _0502_
rlabel metal1 9154 4794 9154 4794 0 _0503_
rlabel metal2 9706 13005 9706 13005 0 _0504_
rlabel metal1 19274 7752 19274 7752 0 _0505_
rlabel metal1 21160 12342 21160 12342 0 _0506_
rlabel metal2 19274 19176 19274 19176 0 _0507_
rlabel metal1 19458 18054 19458 18054 0 _0508_
rlabel metal1 23966 11152 23966 11152 0 _0509_
rlabel metal1 24058 9996 24058 9996 0 _0510_
rlabel metal1 24334 10234 24334 10234 0 _0511_
rlabel metal1 20470 11560 20470 11560 0 _0512_
rlabel metal2 10258 10812 10258 10812 0 _0513_
rlabel metal1 15272 12138 15272 12138 0 _0514_
rlabel metal1 16928 10642 16928 10642 0 _0515_
rlabel metal2 9890 15300 9890 15300 0 _0516_
rlabel metal1 9660 18394 9660 18394 0 _0517_
rlabel metal2 15134 15844 15134 15844 0 _0518_
rlabel metal1 12466 16592 12466 16592 0 _0519_
rlabel metal1 9476 18394 9476 18394 0 _0520_
rlabel metal1 8786 19346 8786 19346 0 _0521_
rlabel metal2 19688 17204 19688 17204 0 _0522_
rlabel via2 20010 12325 20010 12325 0 _0523_
rlabel metal1 19688 11866 19688 11866 0 _0524_
rlabel metal1 19688 12410 19688 12410 0 _0525_
rlabel metal1 20930 13498 20930 13498 0 _0526_
rlabel metal2 20746 14144 20746 14144 0 _0527_
rlabel metal2 20654 11764 20654 11764 0 _0528_
rlabel metal1 20202 13294 20202 13294 0 _0529_
rlabel metal1 19918 13736 19918 13736 0 _0530_
rlabel metal1 16974 20876 16974 20876 0 _0531_
rlabel metal2 20194 14076 20194 14076 0 _0532_
rlabel metal1 21022 13770 21022 13770 0 _0533_
rlabel metal1 19872 13498 19872 13498 0 _0534_
rlabel metal1 20424 12750 20424 12750 0 _0535_
rlabel metal1 20976 20774 20976 20774 0 _0536_
rlabel metal2 20562 14144 20562 14144 0 _0537_
rlabel metal1 20194 12954 20194 12954 0 _0538_
rlabel metal2 17618 13651 17618 13651 0 _0539_
rlabel metal1 16836 15946 16836 15946 0 _0540_
rlabel metal2 18722 15164 18722 15164 0 _0541_
rlabel metal2 14628 14212 14628 14212 0 _0542_
rlabel metal1 15640 16014 15640 16014 0 _0543_
rlabel metal2 16330 7684 16330 7684 0 _0544_
rlabel metal1 16192 8058 16192 8058 0 _0545_
rlabel metal3 15617 15300 15617 15300 0 _0546_
rlabel metal1 15916 9146 15916 9146 0 _0547_
rlabel metal1 15916 8806 15916 8806 0 _0548_
rlabel metal1 15686 10234 15686 10234 0 _0549_
rlabel metal1 15456 10234 15456 10234 0 _0550_
rlabel metal1 19826 15674 19826 15674 0 _0551_
rlabel metal2 17710 18224 17710 18224 0 _0552_
rlabel metal1 17664 21862 17664 21862 0 _0553_
rlabel metal1 16744 15606 16744 15606 0 _0554_
rlabel metal1 15042 16218 15042 16218 0 _0555_
rlabel metal2 12466 18972 12466 18972 0 _0556_
rlabel metal2 12558 20162 12558 20162 0 _0557_
rlabel metal1 19458 21114 19458 21114 0 _0558_
rlabel metal2 18630 19584 18630 19584 0 _0559_
rlabel metal1 19182 20570 19182 20570 0 _0560_
rlabel metal3 20079 20740 20079 20740 0 _0561_
rlabel metal1 14950 9350 14950 9350 0 _0562_
rlabel metal1 14628 9350 14628 9350 0 _0563_
rlabel metal2 14674 9044 14674 9044 0 _0564_
rlabel metal1 13846 9146 13846 9146 0 _0565_
rlabel metal1 15686 5100 15686 5100 0 _0566_
rlabel metal1 13662 5882 13662 5882 0 _0567_
rlabel metal2 12926 5508 12926 5508 0 _0568_
rlabel metal2 13202 7446 13202 7446 0 _0569_
rlabel metal1 13064 7514 13064 7514 0 _0570_
rlabel metal2 12926 6970 12926 6970 0 _0571_
rlabel metal1 12650 7990 12650 7990 0 _0572_
rlabel metal1 12834 8058 12834 8058 0 _0573_
rlabel metal1 13202 9078 13202 9078 0 _0574_
rlabel metal1 14076 13906 14076 13906 0 _0575_
rlabel metal2 13478 15912 13478 15912 0 _0576_
rlabel metal2 17204 21284 17204 21284 0 _0577_
rlabel metal1 17204 22950 17204 22950 0 _0578_
rlabel metal1 18032 19958 18032 19958 0 _0579_
rlabel metal2 17526 19652 17526 19652 0 _0580_
rlabel metal1 17112 19958 17112 19958 0 _0581_
rlabel metal1 17250 20026 17250 20026 0 _0582_
rlabel metal1 20516 6086 20516 6086 0 _0583_
rlabel metal2 20562 5780 20562 5780 0 _0584_
rlabel metal1 20562 5882 20562 5882 0 _0585_
rlabel metal1 19090 14926 19090 14926 0 _0586_
rlabel metal1 13340 18190 13340 18190 0 _0587_
rlabel metal1 11592 16762 11592 16762 0 _0588_
rlabel metal1 10902 19244 10902 19244 0 _0589_
rlabel metal1 10626 18768 10626 18768 0 _0590_
rlabel metal1 9522 19312 9522 19312 0 _0591_
rlabel metal1 9384 20910 9384 20910 0 _0592_
rlabel metal1 18078 13294 18078 13294 0 _0593_
rlabel metal2 17894 9792 17894 9792 0 _0594_
rlabel metal1 17710 13906 17710 13906 0 _0595_
rlabel metal1 16606 13328 16606 13328 0 _0596_
rlabel metal1 17112 13838 17112 13838 0 _0597_
rlabel via3 17227 13124 17227 13124 0 _0598_
rlabel metal2 16974 14552 16974 14552 0 _0599_
rlabel metal2 16698 13600 16698 13600 0 _0600_
rlabel metal2 17158 12988 17158 12988 0 _0601_
rlabel metal1 16790 12818 16790 12818 0 _0602_
rlabel metal3 16905 12580 16905 12580 0 _0603_
rlabel metal2 16698 12954 16698 12954 0 _0604_
rlabel metal2 18308 12852 18308 12852 0 _0605_
rlabel metal1 19090 16694 19090 16694 0 _0606_
rlabel metal2 18078 10404 18078 10404 0 _0607_
rlabel metal1 17434 13192 17434 13192 0 _0608_
rlabel metal2 12006 15708 12006 15708 0 _0609_
rlabel metal1 17986 17782 17986 17782 0 _0610_
rlabel metal2 16790 17952 16790 17952 0 _0611_
rlabel metal2 19918 18156 19918 18156 0 _0612_
rlabel metal2 16606 17034 16606 17034 0 _0613_
rlabel metal1 16790 5814 16790 5814 0 _0614_
rlabel metal1 18446 5780 18446 5780 0 _0615_
rlabel metal1 16606 5338 16606 5338 0 _0616_
rlabel metal2 16882 16711 16882 16711 0 _0617_
rlabel metal1 19044 22610 19044 22610 0 _0618_
rlabel metal2 18952 22542 18952 22542 0 _0619_
rlabel metal1 18814 22610 18814 22610 0 _0620_
rlabel metal1 16790 16660 16790 16660 0 _0621_
rlabel metal1 17296 8602 17296 8602 0 _0622_
rlabel metal1 17526 10506 17526 10506 0 _0623_
rlabel metal1 16974 10778 16974 10778 0 _0624_
rlabel metal1 12190 16660 12190 16660 0 _0625_
rlabel metal1 9660 19346 9660 19346 0 _0626_
rlabel metal2 9154 21216 9154 21216 0 _0627_
rlabel metal1 11592 19278 11592 19278 0 _0628_
rlabel metal2 10212 19142 10212 19142 0 _0629_
rlabel metal1 10028 21522 10028 21522 0 _0630_
rlabel metal1 11822 21420 11822 21420 0 _0631_
rlabel metal1 22632 8058 22632 8058 0 _0632_
rlabel metal1 22356 9690 22356 9690 0 _0633_
rlabel metal2 22218 10336 22218 10336 0 _0634_
rlabel metal1 22402 10778 22402 10778 0 _0635_
rlabel metal2 22862 21216 22862 21216 0 _0636_
rlabel metal1 22540 21386 22540 21386 0 _0637_
rlabel metal1 23000 21862 23000 21862 0 _0638_
rlabel metal2 22402 20128 22402 20128 0 _0639_
rlabel metal2 22862 18156 22862 18156 0 _0640_
rlabel metal3 23023 18020 23023 18020 0 _0641_
rlabel metal1 22862 18292 22862 18292 0 _0642_
rlabel metal2 22586 18564 22586 18564 0 _0643_
rlabel metal1 15456 22746 15456 22746 0 _0644_
rlabel metal1 15548 23290 15548 23290 0 _0645_
rlabel metal1 15180 23222 15180 23222 0 _0646_
rlabel metal1 22126 18632 22126 18632 0 _0647_
rlabel metal4 22724 15504 22724 15504 0 _0648_
rlabel metal1 11316 8466 11316 8466 0 _0649_
rlabel metal2 12144 10574 12144 10574 0 _0650_
rlabel metal1 11132 8330 11132 8330 0 _0651_
rlabel metal1 12190 13158 12190 13158 0 _0652_
rlabel metal1 11132 10234 11132 10234 0 _0653_
rlabel metal1 12466 10472 12466 10472 0 _0654_
rlabel metal1 12696 5882 12696 5882 0 _0655_
rlabel metal2 23736 15130 23736 15130 0 _0656_
rlabel metal1 22034 8602 22034 8602 0 _0657_
rlabel metal2 23782 9656 23782 9656 0 _0658_
rlabel metal1 20838 10064 20838 10064 0 _0659_
rlabel metal2 12282 11832 12282 11832 0 _0660_
rlabel metal1 12236 12954 12236 12954 0 _0661_
rlabel metal1 10028 17782 10028 17782 0 _0662_
rlabel metal1 10718 17680 10718 17680 0 _0663_
rlabel metal1 10764 20910 10764 20910 0 _0664_
rlabel metal1 12282 22168 12282 22168 0 _0665_
rlabel metal1 11132 19890 11132 19890 0 _0666_
rlabel metal1 10626 20026 10626 20026 0 _0667_
rlabel via1 11362 19827 11362 19827 0 _0668_
rlabel metal1 10304 17850 10304 17850 0 _0669_
rlabel metal1 10534 20808 10534 20808 0 _0670_
rlabel metal1 12328 21658 12328 21658 0 _0671_
rlabel metal1 10718 21964 10718 21964 0 _0672_
rlabel metal1 11638 20026 11638 20026 0 _0673_
rlabel metal1 11638 22202 11638 22202 0 _0674_
rlabel metal1 10948 23766 10948 23766 0 _0675_
rlabel metal1 11132 20570 11132 20570 0 _0676_
rlabel metal1 9384 21454 9384 21454 0 _0677_
rlabel metal1 10902 21012 10902 21012 0 _0678_
rlabel metal1 12006 22406 12006 22406 0 _0679_
rlabel metal1 9752 18802 9752 18802 0 _0680_
rlabel metal1 10626 23834 10626 23834 0 _0681_
rlabel metal1 10120 24174 10120 24174 0 _0682_
rlabel viali 21850 11732 21850 11732 0 _0683_
rlabel metal1 21804 17170 21804 17170 0 _0684_
rlabel metal2 22310 23562 22310 23562 0 _0685_
rlabel metal1 22586 22950 22586 22950 0 _0686_
rlabel metal1 21942 5100 21942 5100 0 _0687_
rlabel metal3 23575 15300 23575 15300 0 _0688_
rlabel metal1 22678 16762 22678 16762 0 _0689_
rlabel metal1 16698 26996 16698 26996 0 _0690_
rlabel metal2 16882 19965 16882 19965 0 _0691_
rlabel metal1 20378 17204 20378 17204 0 _0692_
rlabel metal1 9844 9146 9844 9146 0 _0693_
rlabel metal1 10764 9690 10764 9690 0 _0694_
rlabel viali 23966 10644 23966 10644 0 _0695_
rlabel metal1 23322 10540 23322 10540 0 _0696_
rlabel metal1 9338 10132 9338 10132 0 _0697_
rlabel metal1 9384 12614 9384 12614 0 _0698_
rlabel metal1 9430 6834 9430 6834 0 _0699_
rlabel metal1 9108 4114 9108 4114 0 _0700_
rlabel metal2 9522 10472 9522 10472 0 _0701_
rlabel metal1 10350 16626 10350 16626 0 _0702_
rlabel metal1 10028 16762 10028 16762 0 _0703_
rlabel metal1 9016 20026 9016 20026 0 _0704_
rlabel metal1 10442 24208 10442 24208 0 _0705_
rlabel metal1 12328 25262 12328 25262 0 _0706_
rlabel metal1 11362 24242 11362 24242 0 _0707_
rlabel metal1 12282 24208 12282 24208 0 _0708_
rlabel metal1 12052 22202 12052 22202 0 _0709_
rlabel metal1 11316 23086 11316 23086 0 _0710_
rlabel metal1 11822 24174 11822 24174 0 _0711_
rlabel metal1 10672 24174 10672 24174 0 _0712_
rlabel metal2 9614 24820 9614 24820 0 _0713_
rlabel metal1 9844 25262 9844 25262 0 _0714_
rlabel metal1 9660 21658 9660 21658 0 _0715_
rlabel via1 9702 19482 9702 19482 0 _0716_
rlabel metal1 10626 23120 10626 23120 0 _0717_
rlabel metal1 10166 24752 10166 24752 0 _0718_
rlabel metal1 10028 25670 10028 25670 0 _0719_
rlabel metal1 6578 24038 6578 24038 0 _0720_
rlabel metal1 9016 25330 9016 25330 0 _0721_
rlabel metal1 7360 25262 7360 25262 0 _0722_
rlabel metal1 9200 24174 9200 24174 0 _0723_
rlabel metal2 7774 25568 7774 25568 0 _0724_
rlabel metal1 9476 23290 9476 23290 0 _0725_
rlabel metal1 9936 23290 9936 23290 0 _0726_
rlabel metal1 9154 24752 9154 24752 0 _0727_
rlabel metal1 8293 22950 8293 22950 0 _0728_
rlabel metal1 11684 25398 11684 25398 0 _0729_
rlabel metal1 12052 24922 12052 24922 0 _0730_
rlabel metal1 11362 25330 11362 25330 0 _0731_
rlabel metal1 10810 25296 10810 25296 0 _0732_
rlabel metal1 7682 25228 7682 25228 0 _0733_
rlabel metal1 8050 25398 8050 25398 0 _0734_
rlabel metal1 7084 21114 7084 21114 0 _0735_
rlabel metal2 5842 20332 5842 20332 0 _0736_
rlabel metal1 4002 21964 4002 21964 0 _0737_
rlabel metal1 5060 20026 5060 20026 0 _0738_
rlabel metal1 4922 19924 4922 19924 0 _0739_
rlabel via1 5124 19346 5124 19346 0 _0740_
rlabel metal1 4370 17646 4370 17646 0 _0741_
rlabel metal1 3726 19380 3726 19380 0 _0742_
rlabel metal1 2024 18734 2024 18734 0 _0743_
rlabel metal1 3082 18666 3082 18666 0 _0744_
rlabel metal1 2852 19414 2852 19414 0 _0745_
rlabel metal1 2346 21114 2346 21114 0 _0746_
rlabel metal2 4830 20060 4830 20060 0 _0747_
rlabel metal1 8004 25874 8004 25874 0 _0748_
rlabel metal1 8142 25806 8142 25806 0 _0749_
rlabel metal1 6486 25194 6486 25194 0 _0750_
rlabel metal2 6854 24990 6854 24990 0 _0751_
rlabel metal1 7498 24208 7498 24208 0 _0752_
rlabel metal1 3910 22032 3910 22032 0 _0753_
rlabel metal1 2806 17272 2806 17272 0 _0754_
rlabel metal1 7958 21556 7958 21556 0 _0755_
rlabel metal1 4646 21930 4646 21930 0 _0756_
rlabel metal1 4462 22032 4462 22032 0 _0757_
rlabel metal1 5106 22066 5106 22066 0 _0758_
rlabel metal1 5060 20434 5060 20434 0 _0759_
rlabel metal1 4554 20468 4554 20468 0 _0760_
rlabel metal1 2990 19822 2990 19822 0 _0761_
rlabel metal2 2346 20332 2346 20332 0 _0762_
rlabel metal1 1748 21930 1748 21930 0 _0763_
rlabel metal1 8326 19482 8326 19482 0 _0764_
rlabel metal1 8418 19822 8418 19822 0 _0765_
rlabel metal2 8786 20434 8786 20434 0 _0766_
rlabel metal1 6946 20230 6946 20230 0 _0767_
rlabel metal1 5106 20808 5106 20808 0 _0768_
rlabel metal2 5198 20740 5198 20740 0 _0769_
rlabel metal1 3772 21114 3772 21114 0 _0770_
rlabel metal1 3082 21590 3082 21590 0 _0771_
rlabel metal1 2484 21522 2484 21522 0 _0772_
rlabel metal1 5060 24038 5060 24038 0 _0773_
rlabel metal2 8510 22950 8510 22950 0 _0774_
rlabel metal1 8602 22440 8602 22440 0 _0775_
rlabel metal1 7682 23494 7682 23494 0 _0776_
rlabel metal1 7636 21522 7636 21522 0 _0777_
rlabel metal1 7038 21590 7038 21590 0 _0778_
rlabel metal1 6982 21488 6982 21488 0 _0779_
rlabel metal1 4692 21590 4692 21590 0 _0780_
rlabel viali 4277 21522 4277 21522 0 _0781_
rlabel metal1 3542 21658 3542 21658 0 _0782_
rlabel metal1 2806 22576 2806 22576 0 _0783_
rlabel metal2 2714 25092 2714 25092 0 _0784_
rlabel metal1 8556 21658 8556 21658 0 _0785_
rlabel metal1 7314 22678 7314 22678 0 _0786_
rlabel metal1 6394 21318 6394 21318 0 _0787_
rlabel metal1 6348 22610 6348 22610 0 _0788_
rlabel metal1 4876 22746 4876 22746 0 _0789_
rlabel metal1 4048 17850 4048 17850 0 _0790_
rlabel metal1 3220 23834 3220 23834 0 _0791_
rlabel metal1 6394 25296 6394 25296 0 _0792_
rlabel metal1 5750 24752 5750 24752 0 _0793_
rlabel metal1 7774 21386 7774 21386 0 _0794_
rlabel metal1 5888 24786 5888 24786 0 _0795_
rlabel metal1 5290 24242 5290 24242 0 _0796_
rlabel metal1 5428 24174 5428 24174 0 _0797_
rlabel metal1 4968 24378 4968 24378 0 _0798_
rlabel metal1 4370 24922 4370 24922 0 _0799_
rlabel metal2 3358 26758 3358 26758 0 _0800_
rlabel metal2 2346 25670 2346 25670 0 _0801_
rlabel metal1 4002 25330 4002 25330 0 _0802_
rlabel metal1 3680 25262 3680 25262 0 _0803_
rlabel metal1 2599 23494 2599 23494 0 _0804_
rlabel metal1 3772 20570 3772 20570 0 _0805_
rlabel metal1 3450 24378 3450 24378 0 _0806_
rlabel metal1 3082 25228 3082 25228 0 _0807_
rlabel metal1 3910 13260 3910 13260 0 _0808_
rlabel metal1 4830 14416 4830 14416 0 _0809_
rlabel metal1 5244 14382 5244 14382 0 _0810_
rlabel metal2 4646 15079 4646 15079 0 _0811_
rlabel metal1 5290 28560 5290 28560 0 _0812_
rlabel metal1 5888 29138 5888 29138 0 _0813_
rlabel metal1 5704 29274 5704 29274 0 _0814_
rlabel metal2 8510 28730 8510 28730 0 _0815_
rlabel metal2 9338 27642 9338 27642 0 _0816_
rlabel metal1 2484 27438 2484 27438 0 _0817_
rlabel metal1 5750 23290 5750 23290 0 _0818_
rlabel metal1 8280 21318 8280 21318 0 _0819_
rlabel metal1 6026 23630 6026 23630 0 _0820_
rlabel metal1 5060 23834 5060 23834 0 _0821_
rlabel metal1 4416 23834 4416 23834 0 _0822_
rlabel metal1 3450 24038 3450 24038 0 _0823_
rlabel metal1 2438 28118 2438 28118 0 _0824_
rlabel via1 1789 28186 1789 28186 0 _0825_
rlabel metal1 4738 27030 4738 27030 0 _0826_
rlabel metal1 6072 23766 6072 23766 0 _0827_
rlabel metal1 4508 25466 4508 25466 0 _0828_
rlabel metal1 4140 26010 4140 26010 0 _0829_
rlabel metal1 3588 27302 3588 27302 0 _0830_
rlabel metal1 2162 30668 2162 30668 0 _0831_
rlabel metal1 2576 28526 2576 28526 0 _0832_
rlabel metal1 2300 30158 2300 30158 0 _0833_
rlabel metal1 4646 30362 4646 30362 0 _0834_
rlabel metal1 4738 29002 4738 29002 0 _0835_
rlabel metal2 12834 17374 12834 17374 0 _0836_
rlabel metal1 1886 9996 1886 9996 0 _0837_
rlabel metal1 13432 21998 13432 21998 0 _0838_
rlabel metal2 7498 27353 7498 27353 0 _0839_
rlabel metal1 7406 16048 7406 16048 0 _0840_
rlabel metal1 8924 16490 8924 16490 0 _0841_
rlabel metal1 8878 17136 8878 17136 0 _0842_
rlabel metal1 9568 15470 9568 15470 0 _0843_
rlabel metal1 11316 14994 11316 14994 0 _0844_
rlabel metal1 12880 16762 12880 16762 0 _0845_
rlabel metal1 12328 18394 12328 18394 0 _0846_
rlabel metal1 12788 26554 12788 26554 0 _0847_
rlabel metal1 13202 25874 13202 25874 0 _0848_
rlabel metal1 13938 24208 13938 24208 0 _0849_
rlabel metal1 22954 4522 22954 4522 0 _0850_
rlabel metal1 14536 14314 14536 14314 0 _0851_
rlabel metal2 15226 13770 15226 13770 0 _0852_
rlabel metal1 18124 14382 18124 14382 0 _0853_
rlabel metal1 20654 13974 20654 13974 0 _0854_
rlabel metal2 22034 13668 22034 13668 0 _0855_
rlabel metal1 23598 12206 23598 12206 0 _0856_
rlabel metal1 23920 13498 23920 13498 0 _0857_
rlabel metal1 14766 12818 14766 12818 0 _0858_
rlabel metal1 17526 12410 17526 12410 0 _0859_
rlabel metal1 9614 13294 9614 13294 0 _0860_
rlabel metal1 7912 12818 7912 12818 0 _0861_
rlabel metal1 9522 12818 9522 12818 0 _0862_
rlabel metal1 14628 22474 14628 22474 0 _0863_
rlabel metal2 12006 13430 12006 13430 0 _0864_
rlabel metal1 15318 14382 15318 14382 0 _0865_
rlabel metal1 18584 15470 18584 15470 0 _0866_
rlabel metal1 20930 16218 20930 16218 0 _0867_
rlabel metal1 23920 16762 23920 16762 0 _0868_
rlabel metal2 23782 19380 23782 19380 0 _0869_
rlabel metal1 25208 19346 25208 19346 0 _0870_
rlabel metal1 18676 16558 18676 16558 0 _0871_
rlabel metal1 18998 21862 18998 21862 0 _0872_
rlabel metal1 20056 16762 20056 16762 0 _0873_
rlabel metal1 21252 20910 21252 20910 0 _0874_
rlabel metal1 23736 22610 23736 22610 0 _0875_
rlabel metal1 24794 21998 24794 21998 0 _0876_
rlabel metal1 25162 20910 25162 20910 0 _0877_
rlabel metal1 14766 19924 14766 19924 0 _0878_
rlabel metal1 14536 15674 14536 15674 0 _0879_
rlabel metal1 13294 15368 13294 15368 0 _0880_
rlabel metal1 8050 11696 8050 11696 0 _0881_
rlabel metal1 9430 11696 9430 11696 0 _0882_
rlabel metal3 13639 20740 13639 20740 0 _0883_
rlabel metal1 14582 9690 14582 9690 0 cal_lut\[100\]
rlabel metal2 16698 17612 16698 17612 0 cal_lut\[101\]
rlabel metal1 17158 10982 17158 10982 0 cal_lut\[102\]
rlabel metal1 20792 10982 20792 10982 0 cal_lut\[103\]
rlabel metal2 21114 11220 21114 11220 0 cal_lut\[104\]
rlabel metal1 20654 9962 20654 9962 0 cal_lut\[105\]
rlabel metal1 17296 9554 17296 9554 0 cal_lut\[106\]
rlabel metal1 18032 9690 18032 9690 0 cal_lut\[107\]
rlabel via1 20746 9690 20746 9690 0 cal_lut\[108\]
rlabel metal1 23966 8568 23966 8568 0 cal_lut\[109\]
rlabel metal1 15042 14314 15042 14314 0 cal_lut\[10\]
rlabel metal1 24150 11050 24150 11050 0 cal_lut\[110\]
rlabel metal1 21160 8058 21160 8058 0 cal_lut\[111\]
rlabel metal1 16744 7990 16744 7990 0 cal_lut\[112\]
rlabel metal1 18400 6970 18400 6970 0 cal_lut\[113\]
rlabel metal1 21160 12954 21160 12954 0 cal_lut\[114\]
rlabel metal1 22540 4590 22540 4590 0 cal_lut\[115\]
rlabel metal2 23506 4896 23506 4896 0 cal_lut\[116\]
rlabel metal2 19458 3842 19458 3842 0 cal_lut\[117\]
rlabel metal1 20930 5814 20930 5814 0 cal_lut\[118\]
rlabel metal1 15042 6154 15042 6154 0 cal_lut\[119\]
rlabel metal1 16744 14042 16744 14042 0 cal_lut\[11\]
rlabel metal1 8234 8500 8234 8500 0 cal_lut\[120\]
rlabel metal2 8786 9384 8786 9384 0 cal_lut\[121\]
rlabel metal2 9982 8126 9982 8126 0 cal_lut\[122\]
rlabel metal1 11500 7514 11500 7514 0 cal_lut\[123\]
rlabel metal1 13018 7718 13018 7718 0 cal_lut\[124\]
rlabel metal1 15502 7752 15502 7752 0 cal_lut\[125\]
rlabel metal1 15502 9146 15502 9146 0 cal_lut\[126\]
rlabel metal1 9338 6664 9338 6664 0 cal_lut\[127\]
rlabel metal2 10442 5678 10442 5678 0 cal_lut\[128\]
rlabel metal1 12236 5814 12236 5814 0 cal_lut\[129\]
rlabel metal1 19872 14586 19872 14586 0 cal_lut\[12\]
rlabel metal2 12742 4216 12742 4216 0 cal_lut\[130\]
rlabel metal1 14674 3638 14674 3638 0 cal_lut\[131\]
rlabel metal1 15042 4182 15042 4182 0 cal_lut\[132\]
rlabel metal1 8786 4250 8786 4250 0 cal_lut\[133\]
rlabel metal1 8648 3366 8648 3366 0 cal_lut\[134\]
rlabel metal1 6808 5270 6808 5270 0 cal_lut\[135\]
rlabel metal1 12581 4998 12581 4998 0 cal_lut\[136\]
rlabel metal1 14674 6188 14674 6188 0 cal_lut\[137\]
rlabel metal1 12834 7208 12834 7208 0 cal_lut\[138\]
rlabel metal1 7912 9418 7912 9418 0 cal_lut\[139\]
rlabel metal1 22034 13430 22034 13430 0 cal_lut\[13\]
rlabel metal1 6624 9146 6624 9146 0 cal_lut\[140\]
rlabel metal1 5474 8466 5474 8466 0 cal_lut\[141\]
rlabel metal1 4416 7990 4416 7990 0 cal_lut\[142\]
rlabel metal1 14582 6936 14582 6936 0 cal_lut\[143\]
rlabel metal2 12742 7718 12742 7718 0 cal_lut\[144\]
rlabel metal1 8326 6426 8326 6426 0 cal_lut\[145\]
rlabel metal2 9246 4454 9246 4454 0 cal_lut\[146\]
rlabel metal1 11776 3706 11776 3706 0 cal_lut\[147\]
rlabel metal1 13340 2618 13340 2618 0 cal_lut\[148\]
rlabel metal1 15962 1530 15962 1530 0 cal_lut\[149\]
rlabel metal2 23414 12920 23414 12920 0 cal_lut\[14\]
rlabel metal1 18584 2618 18584 2618 0 cal_lut\[150\]
rlabel metal1 22126 1462 22126 1462 0 cal_lut\[151\]
rlabel metal1 22816 2550 22816 2550 0 cal_lut\[152\]
rlabel metal2 22494 6154 22494 6154 0 cal_lut\[153\]
rlabel metal1 20930 2618 20930 2618 0 cal_lut\[154\]
rlabel metal1 18676 2550 18676 2550 0 cal_lut\[155\]
rlabel metal2 19090 4352 19090 4352 0 cal_lut\[156\]
rlabel metal1 21022 6868 21022 6868 0 cal_lut\[157\]
rlabel metal1 22816 6630 22816 6630 0 cal_lut\[158\]
rlabel metal1 23598 6426 23598 6426 0 cal_lut\[159\]
rlabel metal1 23828 12682 23828 12682 0 cal_lut\[15\]
rlabel metal1 20838 6188 20838 6188 0 cal_lut\[160\]
rlabel metal1 20378 5644 20378 5644 0 cal_lut\[161\]
rlabel metal1 20378 12070 20378 12070 0 cal_lut\[162\]
rlabel metal1 24288 7242 24288 7242 0 cal_lut\[163\]
rlabel metal2 24610 8126 24610 8126 0 cal_lut\[164\]
rlabel metal1 25116 9146 25116 9146 0 cal_lut\[165\]
rlabel metal1 25668 8262 25668 8262 0 cal_lut\[166\]
rlabel metal1 18814 10472 18814 10472 0 cal_lut\[167\]
rlabel metal1 22034 15946 22034 15946 0 cal_lut\[168\]
rlabel metal1 24702 10540 24702 10540 0 cal_lut\[169\]
rlabel metal1 15272 13226 15272 13226 0 cal_lut\[16\]
rlabel metal1 26036 9894 26036 9894 0 cal_lut\[170\]
rlabel metal1 26542 10506 26542 10506 0 cal_lut\[171\]
rlabel metal1 27186 11288 27186 11288 0 cal_lut\[172\]
rlabel metal2 17342 13447 17342 13447 0 cal_lut\[173\]
rlabel metal1 24058 13770 24058 13770 0 cal_lut\[174\]
rlabel metal1 25254 12682 25254 12682 0 cal_lut\[175\]
rlabel metal1 24012 11594 24012 11594 0 cal_lut\[176\]
rlabel metal1 16974 3604 16974 3604 0 cal_lut\[177\]
rlabel metal1 15732 3638 15732 3638 0 cal_lut\[178\]
rlabel metal2 16514 4624 16514 4624 0 cal_lut\[179\]
rlabel metal1 16882 12206 16882 12206 0 cal_lut\[17\]
rlabel metal1 9591 2890 9591 2890 0 cal_lut\[180\]
rlabel metal1 9246 2584 9246 2584 0 cal_lut\[181\]
rlabel metal1 9844 1802 9844 1802 0 cal_lut\[182\]
rlabel metal1 11638 1802 11638 1802 0 cal_lut\[183\]
rlabel metal1 13616 1734 13616 1734 0 cal_lut\[184\]
rlabel metal1 18124 1462 18124 1462 0 cal_lut\[185\]
rlabel metal1 13570 2380 13570 2380 0 cal_lut\[186\]
rlabel metal1 7958 2618 7958 2618 0 cal_lut\[187\]
rlabel metal1 6900 10438 6900 10438 0 cal_lut\[188\]
rlabel metal1 4876 10438 4876 10438 0 cal_lut\[189\]
rlabel metal2 20010 13158 20010 13158 0 cal_lut\[18\]
rlabel metal1 6716 11594 6716 11594 0 cal_lut\[190\]
rlabel metal1 16146 12376 16146 12376 0 cal_lut\[191\]
rlabel metal1 14950 12410 14950 12410 0 cal_lut\[192\]
rlabel metal1 8372 12614 8372 12614 0 cal_lut\[19\]
rlabel metal1 6762 15912 6762 15912 0 cal_lut\[1\]
rlabel metal1 9016 13498 9016 13498 0 cal_lut\[20\]
rlabel via1 11454 13294 11454 13294 0 cal_lut\[21\]
rlabel metal1 14306 13974 14306 13974 0 cal_lut\[22\]
rlabel metal1 18216 15130 18216 15130 0 cal_lut\[23\]
rlabel metal1 20562 15334 20562 15334 0 cal_lut\[24\]
rlabel metal1 23138 16456 23138 16456 0 cal_lut\[25\]
rlabel metal1 23322 17680 23322 17680 0 cal_lut\[26\]
rlabel metal2 24610 19040 24610 19040 0 cal_lut\[27\]
rlabel metal1 18630 19992 18630 19992 0 cal_lut\[28\]
rlabel metal2 19918 16762 19918 16762 0 cal_lut\[29\]
rlabel metal1 8970 16762 8970 16762 0 cal_lut\[2\]
rlabel metal1 21252 17306 21252 17306 0 cal_lut\[30\]
rlabel metal1 23506 22508 23506 22508 0 cal_lut\[31\]
rlabel metal1 24932 22474 24932 22474 0 cal_lut\[32\]
rlabel metal2 24886 21658 24886 21658 0 cal_lut\[33\]
rlabel metal1 17710 19856 17710 19856 0 cal_lut\[34\]
rlabel metal1 16284 19686 16284 19686 0 cal_lut\[35\]
rlabel metal2 15042 15742 15042 15742 0 cal_lut\[36\]
rlabel metal1 8510 11594 8510 11594 0 cal_lut\[37\]
rlabel metal2 9062 11390 9062 11390 0 cal_lut\[38\]
rlabel metal1 11546 11594 11546 11594 0 cal_lut\[39\]
rlabel metal2 9430 17170 9430 17170 0 cal_lut\[3\]
rlabel metal1 14812 20910 14812 20910 0 cal_lut\[40\]
rlabel metal1 16284 21522 16284 21522 0 cal_lut\[41\]
rlabel metal2 17526 21488 17526 21488 0 cal_lut\[42\]
rlabel metal1 17480 27574 17480 27574 0 cal_lut\[43\]
rlabel metal1 16008 29750 16008 29750 0 cal_lut\[44\]
rlabel metal1 16008 25738 16008 25738 0 cal_lut\[45\]
rlabel metal1 17066 25160 17066 25160 0 cal_lut\[46\]
rlabel metal1 18814 25126 18814 25126 0 cal_lut\[47\]
rlabel metal1 20010 25670 20010 25670 0 cal_lut\[48\]
rlabel metal1 14306 29716 14306 29716 0 cal_lut\[49\]
rlabel metal2 10994 16354 10994 16354 0 cal_lut\[4\]
rlabel metal2 14582 28798 14582 28798 0 cal_lut\[50\]
rlabel metal1 15778 29478 15778 29478 0 cal_lut\[51\]
rlabel metal1 19228 20774 19228 20774 0 cal_lut\[52\]
rlabel metal2 20194 20509 20194 20509 0 cal_lut\[53\]
rlabel metal1 20884 21114 20884 21114 0 cal_lut\[54\]
rlabel metal1 22724 27846 22724 27846 0 cal_lut\[55\]
rlabel metal2 22954 25296 22954 25296 0 cal_lut\[56\]
rlabel metal1 23092 21114 23092 21114 0 cal_lut\[57\]
rlabel metal1 18814 20298 18814 20298 0 cal_lut\[58\]
rlabel metal1 20332 19754 20332 19754 0 cal_lut\[59\]
rlabel metal1 12466 16456 12466 16456 0 cal_lut\[5\]
rlabel metal1 21574 20026 21574 20026 0 cal_lut\[60\]
rlabel via1 23230 24174 23230 24174 0 cal_lut\[61\]
rlabel metal2 24978 23868 24978 23868 0 cal_lut\[62\]
rlabel metal1 25990 22474 25990 22474 0 cal_lut\[63\]
rlabel metal1 20102 21998 20102 21998 0 cal_lut\[64\]
rlabel metal1 19780 22134 19780 22134 0 cal_lut\[65\]
rlabel metal1 21344 15470 21344 15470 0 cal_lut\[66\]
rlabel metal1 23690 14518 23690 14518 0 cal_lut\[67\]
rlabel metal1 24978 14858 24978 14858 0 cal_lut\[68\]
rlabel metal2 25898 15742 25898 15742 0 cal_lut\[69\]
rlabel metal2 12650 18054 12650 18054 0 cal_lut\[6\]
rlabel metal2 18722 18734 18722 18734 0 cal_lut\[70\]
rlabel metal1 26128 17646 26128 17646 0 cal_lut\[71\]
rlabel metal1 26174 16048 26174 16048 0 cal_lut\[72\]
rlabel metal1 26542 16422 26542 16422 0 cal_lut\[73\]
rlabel metal1 24886 17646 24886 17646 0 cal_lut\[74\]
rlabel metal1 25990 18326 25990 18326 0 cal_lut\[75\]
rlabel metal1 17710 19176 17710 19176 0 cal_lut\[76\]
rlabel metal1 17940 16490 17940 16490 0 cal_lut\[77\]
rlabel metal1 16652 16218 16652 16218 0 cal_lut\[78\]
rlabel metal1 9430 14790 9430 14790 0 cal_lut\[79\]
rlabel metal1 13938 26758 13938 26758 0 cal_lut\[7\]
rlabel metal1 10166 13906 10166 13906 0 cal_lut\[80\]
rlabel metal1 11868 14246 11868 14246 0 cal_lut\[81\]
rlabel metal1 17250 23086 17250 23086 0 cal_lut\[82\]
rlabel metal1 19090 24106 19090 24106 0 cal_lut\[83\]
rlabel metal1 20102 24582 20102 24582 0 cal_lut\[84\]
rlabel metal1 22034 24752 22034 24752 0 cal_lut\[85\]
rlabel metal1 23598 25160 23598 25160 0 cal_lut\[86\]
rlabel metal1 22356 21454 22356 21454 0 cal_lut\[87\]
rlabel metal2 17342 26146 17342 26146 0 cal_lut\[88\]
rlabel metal1 18906 26248 18906 26248 0 cal_lut\[89\]
rlabel metal1 13478 27302 13478 27302 0 cal_lut\[8\]
rlabel metal2 20654 25840 20654 25840 0 cal_lut\[90\]
rlabel metal1 16846 27030 16846 27030 0 cal_lut\[91\]
rlabel metal1 15088 27846 15088 27846 0 cal_lut\[92\]
rlabel metal1 14628 25398 14628 25398 0 cal_lut\[93\]
rlabel metal1 16192 24650 16192 24650 0 cal_lut\[94\]
rlabel metal1 15824 18326 15824 18326 0 cal_lut\[95\]
rlabel metal1 16238 16048 16238 16048 0 cal_lut\[96\]
rlabel metal1 13386 14246 13386 14246 0 cal_lut\[97\]
rlabel metal2 12006 10574 12006 10574 0 cal_lut\[98\]
rlabel metal1 12006 8534 12006 8534 0 cal_lut\[99\]
rlabel metal1 13754 24310 13754 24310 0 cal_lut\[9\]
rlabel metal1 8004 19822 8004 19822 0 clknet_0__0380_
rlabel metal1 6900 20570 6900 20570 0 clknet_0_io_in[0]
rlabel metal1 5336 17306 5336 17306 0 clknet_0_net67
rlabel metal1 3036 8602 3036 8602 0 clknet_0_temp1.dcdel_capnode_notouch_
rlabel metal1 3726 24582 3726 24582 0 clknet_0_temp1.i_precharge_n
rlabel metal1 6578 17136 6578 17136 0 clknet_1_0__leaf__0380_
rlabel metal1 1426 12852 1426 12852 0 clknet_1_0__leaf_io_in[0]
rlabel metal1 3358 15470 3358 15470 0 clknet_1_0__leaf_net67
rlabel metal1 1656 6766 1656 6766 0 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_
rlabel metal1 2944 24106 2944 24106 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal1 8280 19414 8280 19414 0 clknet_1_1__leaf__0380_
rlabel metal1 1794 21590 1794 21590 0 clknet_1_1__leaf_io_in[0]
rlabel metal2 3634 16558 3634 16558 0 clknet_1_1__leaf_net67
rlabel metal1 2438 10676 2438 10676 0 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_
rlabel metal2 2162 26112 2162 26112 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal2 2714 14382 2714 14382 0 ctr\[0\]
rlabel metal1 7544 29206 7544 29206 0 ctr\[10\]
rlabel via3 6739 21828 6739 21828 0 ctr\[11\]
rlabel metal1 8142 26894 8142 26894 0 ctr\[12\]
rlabel metal2 4830 21760 4830 21760 0 ctr\[1\]
rlabel metal1 3542 14382 3542 14382 0 ctr\[2\]
rlabel metal1 3266 14246 3266 14246 0 ctr\[3\]
rlabel metal1 5750 22644 5750 22644 0 ctr\[4\]
rlabel metal1 6256 13498 6256 13498 0 ctr\[5\]
rlabel metal1 5290 15538 5290 15538 0 ctr\[6\]
rlabel metal1 7084 26894 7084 26894 0 ctr\[7\]
rlabel metal1 5336 26350 5336 26350 0 ctr\[8\]
rlabel metal1 5980 21998 5980 21998 0 ctr\[9\]
rlabel metal1 13478 3944 13478 3944 0 dbg_delay
rlabel metal2 14260 9452 14260 9452 0 dbg_result[0]
rlabel metal1 14122 17578 14122 17578 0 dbg_result[1]
rlabel metal1 21942 18836 21942 18836 0 dbg_result[2]
rlabel metal1 19918 19448 19918 19448 0 dbg_result[3]
rlabel metal1 17618 21522 17618 21522 0 dbg_result[4]
rlabel metal1 14306 28424 14306 28424 0 dbg_result[5]
rlabel metal1 8740 24718 8740 24718 0 dec1.i_ones
rlabel metal3 3419 2516 3419 2516 0 io_in[0]
rlabel metal3 544 4420 544 4420 0 io_in[1]
rlabel metal3 544 6324 544 6324 0 io_in[2]
rlabel metal3 866 8228 866 8228 0 io_in[3]
rlabel metal3 544 10132 544 10132 0 io_in[4]
rlabel metal3 544 12036 544 12036 0 io_in[5]
rlabel metal3 544 13940 544 13940 0 io_in[6]
rlabel metal3 544 15844 544 15844 0 io_in[7]
rlabel metal2 2806 18479 2806 18479 0 io_out[0]
rlabel metal3 544 19652 544 19652 0 io_out[1]
rlabel metal3 820 21556 820 21556 0 io_out[2]
rlabel metal1 2507 22678 2507 22678 0 io_out[3]
rlabel metal3 567 25364 567 25364 0 io_out[4]
rlabel metal2 2806 26299 2806 26299 0 io_out[5]
rlabel metal2 1610 28951 1610 28951 0 io_out[6]
rlabel metal1 1518 30906 1518 30906 0 io_out[7]
rlabel metal1 2254 9520 2254 9520 0 net1
rlabel metal1 10074 31858 10074 31858 0 net10
rlabel metal1 9062 31858 9062 31858 0 net11
rlabel metal1 10488 17646 10488 17646 0 net12
rlabel metal1 11684 30226 11684 30226 0 net13
rlabel metal1 10258 30838 10258 30838 0 net14
rlabel metal1 13432 18802 13432 18802 0 net15
rlabel metal1 12834 18700 12834 18700 0 net16
rlabel metal3 14191 20740 14191 20740 0 net17
rlabel metal1 23552 17170 23552 17170 0 net18
rlabel metal2 21252 12614 21252 12614 0 net19
rlabel metal1 3542 7786 3542 7786 0 net2
rlabel metal1 19696 14246 19696 14246 0 net20
rlabel metal1 5244 19278 5244 19278 0 net21
rlabel metal1 1978 19754 1978 19754 0 net22
rlabel metal1 8832 6222 8832 6222 0 net23
rlabel metal1 4554 7990 4554 7990 0 net24
rlabel metal1 14122 1292 14122 1292 0 net25
rlabel metal1 14628 1870 14628 1870 0 net26
rlabel metal2 6394 12585 6394 12585 0 net27
rlabel metal1 6808 13362 6808 13362 0 net28
rlabel metal1 12696 9554 12696 9554 0 net29
rlabel metal2 2806 9282 2806 9282 0 net3
rlabel metal2 13018 13566 13018 13566 0 net30
rlabel metal1 17204 2414 17204 2414 0 net31
rlabel metal1 19734 7820 19734 7820 0 net32
rlabel metal1 21942 4046 21942 4046 0 net33
rlabel metal1 23230 6800 23230 6800 0 net34
rlabel metal1 18216 13838 18216 13838 0 net35
rlabel metal1 25024 12818 25024 12818 0 net36
rlabel metal1 22632 15334 22632 15334 0 net37
rlabel metal1 19228 15470 19228 15470 0 net38
rlabel metal1 17388 7378 17388 7378 0 net39
rlabel metal2 1610 10336 1610 10336 0 net4
rlabel metal1 14720 29138 14720 29138 0 net40
rlabel metal1 13662 15980 13662 15980 0 net41
rlabel metal1 21482 17510 21482 17510 0 net42
rlabel metal2 22586 20672 22586 20672 0 net43
rlabel metal1 17894 22032 17894 22032 0 net44
rlabel metal1 21068 25262 21068 25262 0 net45
rlabel metal1 17526 26316 17526 26316 0 net46
rlabel metal2 21666 26724 21666 26724 0 net47
rlabel via2 16698 16541 16698 16541 0 net48
rlabel metal1 2898 7310 2898 7310 0 net49
rlabel metal1 1886 16966 1886 16966 0 net5
rlabel metal1 2622 10710 2622 10710 0 net50
rlabel metal1 2622 10098 2622 10098 0 net51
rlabel metal1 1932 8466 1932 8466 0 net52
rlabel metal1 1886 8874 1886 8874 0 net53
rlabel metal2 1794 7582 1794 7582 0 net54
rlabel metal1 2254 8976 2254 8976 0 net55
rlabel metal1 2254 6358 2254 6358 0 net56
rlabel metal1 2576 8942 2576 8942 0 net57
rlabel metal1 2024 9554 2024 9554 0 net58
rlabel metal1 2254 7310 2254 7310 0 net59
rlabel metal2 1610 15538 1610 15538 0 net6
rlabel metal1 2898 7446 2898 7446 0 net60
rlabel metal1 1886 6358 1886 6358 0 net61
rlabel metal2 1610 9792 1610 9792 0 net62
rlabel metal1 2346 7446 2346 7446 0 net63
rlabel metal1 1702 8976 1702 8976 0 net64
rlabel metal1 11132 31858 11132 31858 0 net65
rlabel metal1 4094 30090 4094 30090 0 net66
rlabel metal2 3864 16524 3864 16524 0 net67
rlabel metal1 4278 15504 4278 15504 0 net68
rlabel metal1 3910 16218 3910 16218 0 net69
rlabel metal1 1840 17238 1840 17238 0 net7
rlabel metal2 3358 27676 3358 27676 0 net70
rlabel metal1 7866 28458 7866 28458 0 net71
rlabel metal2 5198 13311 5198 13311 0 net72
rlabel metal1 7636 28050 7636 28050 0 net73
rlabel metal1 5934 28152 5934 28152 0 net74
rlabel metal1 4600 11730 4600 11730 0 net75
rlabel metal1 7084 26350 7084 26350 0 net76
rlabel metal1 5014 14348 5014 14348 0 net77
rlabel metal1 8832 28526 8832 28526 0 net78
rlabel metal1 5474 28492 5474 28492 0 net79
rlabel metal1 12926 30124 12926 30124 0 net8
rlabel metal1 17710 13260 17710 13260 0 net80
rlabel metal1 15423 22950 15423 22950 0 net81
rlabel metal1 11914 30702 11914 30702 0 net9
rlabel metal2 2162 28288 2162 28288 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal1 2300 28526 2300 28526 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal1 3266 28084 3266 28084 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal1 2070 27506 2070 27506 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 2254 26384 2254 26384 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal1 1978 26894 1978 26894 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal2 1886 30124 1886 30124 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal1 2484 30770 2484 30770 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel via1 2162 21845 2162 21845 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 3956 31790 3956 31790 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal1 5060 31790 5060 31790 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal1 4784 32334 4784 32334 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 9798 30124 9798 30124 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal1 8832 31790 8832 31790 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal1 10258 29818 10258 29818 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal1 3358 29818 3358 29818 0 temp1.dac.vdac_single.en_pupd
rlabel metal1 4324 32198 4324 32198 0 temp1.dac_vout_notouch_
rlabel metal3 3887 9588 3887 9588 0 temp1.dcdel_capnode_notouch_
rlabel metal1 2714 24752 2714 24752 0 temp1.i_precharge_n
rlabel metal1 4278 15980 4278 15980 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>

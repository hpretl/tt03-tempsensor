* PEX produced on Wed Dec 27 09:39:50 AM CET 2023 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from hpretl_tt03_temperature_sensor.ext - technology: sky130A

.subckt hpretl_tt03_temperature_sensor
+ io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ dbg_result[0] dbg_result[1] dbg_result[2] dbg_result[3] dbg_result[4] dbg_result[5]
+ dbg_delay
+ vccd1 vssd1
X0 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 vccd1 _0111_ a_18673_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2 vccd1 a_15963_28853# a_15879_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3 a_13639_2589# a_13459_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4 a_15439_2388# _0366_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5 a_9963_9295# _0493_ a_10141_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 cal_lut\[149\] a_15135_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_14829_27497# cal_lut\[49\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X8 a_22361_21807# a_21371_21807# a_22235_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9 a_24477_15113# a_23487_14741# a_24351_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10 a_27253_9661# a_26983_9295# a_27163_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11 vssd1 a_18482_12533# a_18440_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 vssd1 a_2271_14735# a_2439_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_9096_27221# _0816_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X16 a_8533_22671# _0776_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X17 cal_lut\[94\] a_15043_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 _0467_ a_15370_19407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_12407_10901# a_12691_10901# a_12626_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X20 a_15623_26324# _0219_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X21 vccd1 _0680_ _0682_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X22 a_4348_20495# _0427_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X23 a_26519_7119# a_26339_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
R0 temp1.dac.vdac_single.einvp_batch\[0\].vref_65.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X24 vccd1 a_22863_23413# a_22779_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X25 a_12962_27359# a_12794_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X27 vssd1 a_4963_10601# a_4970_10505# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X28 vccd1 net8 a_11619_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X29 _0455_ _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X30 vccd1 a_17381_15425# _0554_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X32 a_2695_20969# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X33 vccd1 a_15779_13621# a_15695_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X34 vssd1 _0283_ a_19333_9991# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 vccd1 a_3399_10601# a_3406_10505# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X36 cal_lut\[94\] a_15043_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_13722_20175# a_13942_20149# _0485_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 vssd1 a_22403_16635# a_22361_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X39 a_4797_29423# _0208_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X41 a_10659_3829# cal_lut\[132\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X42 a_16179_29397# a_16355_29397# a_16307_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X44 a_14913_13653# a_14747_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 a_22855_27247# a_22726_27521# a_22435_27221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X46 vccd1 a_4912_8439# net24 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X47 a_20893_9839# a_20727_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X49 vccd1 a_20132_19394# a_19915_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.0672 ps=0.74 w=0.42 l=0.15
X50 _0168_ a_26155_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X51 vssd1 a_23211_6575# net33 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X52 a_21591_10205# a_20727_9839# a_21334_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X53 vssd1 _0467_ a_15177_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X54 vssd1 a_3851_25045# _0803_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X55 a_19126_16885# a_18958_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X56 a_14674_9295# _0563_ a_14594_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X57 a_8300_31375# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X58 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X59 a_23631_17143# a_23922_17033# a_23873_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X60 a_21889_4943# _0687_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X61 a_12162_5737# _0502_ a_12162_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X63 a_16679_28879# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X64 a_22291_2589# _0330_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X67 a_17213_9295# a_16679_9301# a_17118_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X68 a_14385_10927# cal_lut\[172\] a_14313_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X69 vccd1 a_24455_13255# cal_lut\[16\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X72 a_7492_27247# a_7093_27247# a_7366_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X75 vssd1 net45 a_21831_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X76 vssd1 _0290_ a_14331_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X77 _0631_ _0627_ a_10521_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X79 a_14591_3855# a_13809_3861# a_14507_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X81 a_21261_10205# a_20727_9839# a_21166_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X82 cal_lut\[9\] a_13571_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X83 cal_lut\[110\] a_23875_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X84 a_4472_21807# _0747_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X85 vccd1 a_3891_17455# _0755_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X86 _0219_ a_15479_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X87 a_27161_10927# a_26891_11293# a_27071_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X88 a_13512_13621# _0575_ a_13904_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X89 net26 a_10659_7637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X90 vssd1 _0323_ a_2971_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X94 vssd1 net25 a_9963_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X95 a_22185_8207# _0108_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X96 a_26210_9951# a_26042_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X98 _0439_ _0438_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X99 vssd1 net25 a_12079_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X100 a_1932_17271# net5 a_1860_17271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X101 a_23351_7338# _0289_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X102 a_6319_11293# a_5621_10927# a_6062_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X103 a_3781_12565# a_3615_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X105 a_23147_3855# a_22365_3861# a_23063_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X106 _0648_ a_22383_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X107 a_13674_7235# _0299_ a_13592_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X108 a_28057_15279# a_27510_15553# a_27710_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X109 vssd1 _0456_ a_20992_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X111 vssd1 a_11030_27383# a_10968_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X112 a_8104_18543# a_7111_18543# a_7975_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X113 vccd1 a_17651_8181# _0450_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X114 vssd1 a_6633_26703# a_6739_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X115 _0067_ a_23671_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X116 a_27978_13647# a_27731_14025# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X118 vccd1 _0277_ a_12263_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X119 a_8483_31849# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X120 a_9117_14191# a_8951_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X121 _0397_ ctr\[4\] a_3974_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X122 a_24573_7125# a_24407_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X124 a_25755_20393# net43 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X125 a_12659_26703# a_11877_26709# a_12575_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 a_10764_29967# a_10515_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X127 a_5158_6031# a_4885_6037# a_5073_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X128 vccd1 a_21115_21237# a_21031_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X129 a_15469_3855# _0178_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X130 a_22438_8181# a_22270_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X131 a_3965_8751# a_3799_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X132 vccd1 a_10570_3423# a_10497_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X134 a_11001_22923# _0675_ a_10915_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X135 vssd1 _0418_ a_4708_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X136 vssd1 a_21334_2335# a_21292_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X137 vccd1 _0378_ a_12815_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X138 a_26861_13103# a_26307_13077# a_26514_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X139 a_12289_21807# _0671_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X140 a_17283_28853# cal_lut\[43\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X141 a_15356_15529# _0505_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X142 a_9209_22895# _0704_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X143 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X145 a_24972_25071# a_24573_25071# a_24846_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X146 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X147 vccd1 _0874_ a_21279_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X148 vccd1 a_21878_17143# _0692_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X149 a_14139_4943# a_13275_4949# a_13882_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X151 a_16307_29423# cal_lut\[44\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X152 a_18475_19783# _0453_ a_18709_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X153 a_2376_30199# _0801_ a_2518_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X154 _0646_ a_14287_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X155 a_16281_20541# cal_lut\[41\] a_16209_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X157 a_24971_19631# a_24835_19605# a_24551_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X158 _0148_ a_14103_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X159 _0372_ a_16859_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X160 a_1573_12565# a_1407_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X161 a_16761_24847# cal_lut\[94\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X162 a_5326_14709# a_5158_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X163 a_1656_29673# a_1407_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X164 io_out[5] a_2564_25045# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X165 vccd1 a_20287_28603# a_20203_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X166 a_15737_2057# a_14747_1685# a_15611_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X167 vssd1 net33 a_21831_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X168 vccd1 a_17459_29185# a_17283_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X169 a_9769_17705# cal_lut\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X172 a_7157_19319# clknet_1_1__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 vccd1 a_10379_6740# _0122_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X174 a_18617_5309# cal_lut\[156\] a_18545_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X176 _0030_ a_21279_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X177 vssd1 a_9558_1247# a_9516_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X178 vssd1 _0567_ a_13241_5633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X179 a_7101_23439# _0750_ a_6955_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X180 temp1.capload\[1\].cap.Y clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X181 vccd1 a_4951_7338# _0142_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X182 vssd1 a_24823_15444# _0068_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X183 vccd1 ctr\[10\] a_7381_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X184 vssd1 _0474_ a_18455_18337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X185 a_19977_14709# _0459_ a_20223_15073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X186 a_14855_12265# _0514_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X187 a_10313_19203# _0589_ a_10241_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X188 a_28031_17821# a_27333_17455# a_27774_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X189 a_20847_1679# a_20065_1685# a_20763_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X190 vccd1 a_6519_21495# _0780_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X191 net7 a_1407_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X192 a_18045_3311# _0155_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X193 a_22645_6031# _0158_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X194 vssd1 a_20322_7775# a_20280_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X195 a_23565_19087# _0026_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X196 a_23355_10615# _0695_ a_23683_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X199 _0173_ a_27903_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X200 a_8688_15113# a_8289_14741# a_8562_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X201 a_4679_10615# a_4970_10505# a_4921_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X203 a_8769_17999# _0520_ a_8645_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.235 ps=1.47 w=1 l=0.15
X205 vccd1 _0414_ _0415_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X206 vccd1 cal_lut\[71\] a_19303_17607# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X207 vssd1 a_20451_23439# _0460_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X208 vccd1 a_23535_17143# cal_lut\[26\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X209 vssd1 cal_lut\[142\] a_4253_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X210 vccd1 a_10699_4399# _0850_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X211 a_25355_25437# a_24573_25071# a_25271_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 vssd1 clknet_1_1__leaf_io_in[0] a_4443_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X213 vccd1 a_18355_25339# a_18271_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X214 vssd1 _0380_ a_7102_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X215 a_4824_5487# a_4425_5487# a_4698_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X216 vccd1 a_5105_25045# a_5135_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X217 vccd1 a_16640_4373# net31 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X218 a_27639_15279# a_27510_15553# a_27219_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X219 cal_lut\[118\] a_20287_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X220 a_11970_9117# a_11723_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X221 a_7373_25071# _0722_ a_7071_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X224 vccd1 dbg_result[1] a_20543_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X225 vccd1 cal_lut\[113\] a_18107_8439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X226 a_16734_21919# a_16566_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X228 vssd1 net71 _0405_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X229 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X230 vccd1 a_14331_29397# a_14155_29397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X231 a_10247_21583# _0591_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X232 a_16574_17455# cal_lut\[101\] a_16493_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X233 a_27203_22173# a_26505_21807# a_26946_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X234 a_22089_14741# a_21923_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X235 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_2596_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X236 vssd1 a_3175_14459# ctr\[3\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X237 _0369_ a_9591_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X238 temp1.capload\[10\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X239 a_6019_27247# a_5890_27521# a_5599_27221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X240 vccd1 net40 a_12355_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X242 a_19797_13353# _0525_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X243 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X244 a_25471_11989# a_25762_12289# a_25713_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X245 a_19862_15391# a_19694_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X246 vccd1 net31 a_20727_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X247 cal_lut\[32\] a_25439_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X248 vccd1 a_1639_15444# _0199_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X249 a_22898_6005# a_22730_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X250 vssd1 a_25014_7093# a_24972_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X252 vccd1 a_28199_17723# a_28115_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X254 a_18409_12559# a_17875_12565# a_18314_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X255 _0058_ a_22659_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X256 _0698_ a_8951_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X257 vccd1 net67 a_3882_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X258 _0348_ a_24035_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X259 vccd1 a_15335_7119# a_15503_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X260 vccd1 ctr\[6\] a_3991_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X261 vccd1 a_24827_24501# _0238_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X263 a_9876_4399# _0502_ a_9385_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X264 _0506_ a_20943_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X265 vccd1 ctr\[3\] a_5359_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X266 a_8123_16911# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X267 vccd1 a_12723_21807# _0237_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X269 a_21218_27497# _0222_ a_21136_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X270 vccd1 a_7959_27515# dec1.i_ones vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X271 a_15531_24135# _0460_ a_15765_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X272 vccd1 a_21334_9951# a_21261_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X273 vccd1 _0352_ a_25327_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_10975_20969# _0678_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X275 vccd1 cal_lut\[78\] a_17812_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X276 a_6007_8029# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X277 vssd1 a_15427_10383# a_15595_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R1 vssd1 net53 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X278 vssd1 _0863_ a_8351_11777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X279 vssd1 _0783_ a_2287_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X280 vssd1 a_14415_26703# a_14583_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X282 vssd1 a_15535_24501# _0273_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X283 vssd1 a_22235_22173# a_22403_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X284 vssd1 a_12355_21271# _0266_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 vccd1 cal_lut\[6\] a_12545_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X286 vccd1 a_22247_9991# _0634_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X287 a_18397_19453# cal_lut\[70\] a_18325_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X289 vssd1 _0491_ _0515_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X290 _0184_ a_14379_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X291 a_4435_30511# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X292 vssd1 a_11765_17973# _0589_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X293 _0737_ _0421_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X295 a_4187_28918# _0800_ a_4115_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X296 vssd1 a_4461_25913# a_4395_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X297 a_27106_17027# _0246_ a_27024_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X298 a_20947_3677# a_20083_3311# a_20690_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X299 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X300 vssd1 a_12955_3476# _0130_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X301 a_22319_16733# a_21537_16367# a_22235_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X302 a_25891_12015# a_25762_12289# a_25471_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X304 a_18489_28169# a_17942_27913# a_18142_28068# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X306 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6835_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X307 vssd1 net8 a_10975_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X309 vssd1 a_16423_25339# a_16381_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X310 a_18685_16917# a_18519_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X311 vccd1 a_8532_31751# a_8483_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X312 a_21166_25437# a_20727_25071# a_21081_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X313 vssd1 a_17095_16055# cal_lut\[78\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X314 vccd1 _0441_ a_16757_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 vssd1 a_2235_9303# _0838_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X316 vssd1 a_18669_22325# _0621_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X317 a_14465_9839# a_14195_10205# a_14375_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X319 temp1.dac_vout_notouch_ net13 a_10764_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X320 a_5801_26409# ctr\[9\] a_5547_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X322 a_4805_19407# _0427_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X323 a_12525_14191# _0096_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X324 a_7987_9514# _0302_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X325 vccd1 _0266_ a_11711_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X326 vssd1 a_17498_29397# a_17427_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X327 vccd1 _0839_ a_10423_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X328 vssd1 _0519_ a_12437_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 a_12981_9301# a_12815_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X331 vccd1 a_24915_21959# cal_lut\[33\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X332 vccd1 cal_lut\[124\] a_13028_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X333 a_14353_18793# _0447_ a_14103_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X334 a_27606_11471# a_27167_11477# a_27521_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X335 a_24101_27081# a_23547_26921# a_23754_26980# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X336 a_22813_19631# a_22259_19605# a_22466_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X337 a_14277_13647# _0456_ a_14131_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X338 vssd1 a_4647_12533# a_4605_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X339 a_15377_19631# _0034_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X340 vssd1 a_5897_28335# a_6003_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X341 vssd1 _0800_ _0801_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X342 vccd1 _0467_ a_16035_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X343 a_18335_6031# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X344 vssd1 _0176_ a_25757_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X346 vccd1 a_18142_28068# a_18071_28169# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X347 vssd1 _0590_ a_9933_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X349 a_19343_3855# a_19163_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X350 a_3859_7337# net24 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X352 a_7826_9117# a_7553_8751# a_7741_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X353 _0380_ a_2879_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X354 vccd1 cal_lut\[160\] a_24771_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X355 _0356_ a_27163_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X357 a_22181_17027# _0689_ a_22109_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X358 a_21292_10927# a_20893_10927# a_21166_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X359 a_5399_8029# a_4535_7663# a_5142_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X360 a_19537_17455# cal_lut\[71\] a_19465_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X361 a_27590_7093# a_27422_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X362 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_1656_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X363 _0379_ a_3575_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X364 a_14223_28879# a_13441_28885# a_14139_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X365 _0332_ a_13639_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X366 _0632_ a_22291_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X367 a_22649_24233# _0469_ a_22503_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X368 _0469_ a_19287_21835# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X370 a_20758_5059# _0283_ a_20676_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X371 vssd1 a_15135_7931# a_15093_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X372 a_7277_2589# a_6743_2223# a_7182_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X373 vssd1 a_25991_23413# a_25949_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X374 _0177_ a_16955_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X375 vssd1 net41 a_14931_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X376 vssd1 a_21683_14557# a_21851_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X378 vssd1 _0448_ a_14747_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X379 a_24846_7119# a_24407_7125# a_24761_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X381 vccd1 a_12035_26324# _0006_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X382 a_4774_27765# a_4606_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X383 a_15356_14441# cal_lut\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X384 a_5031_27791# a_4333_27797# a_4774_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X385 a_19785_25993# a_18795_25621# a_19659_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X386 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X387 vccd1 net37 a_23487_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X389 a_19820_24905# a_19421_24533# a_19694_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X391 a_6729_30199# _0814_ a_6892_30083# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X392 a_6458_20175# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X393 a_8293_15823# _0002_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X394 _0437_ a_7111_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X395 vssd1 _0686_ a_21878_17143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X396 a_3990_19631# _0420_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.12 ps=1.04 w=0.65 l=0.15
X397 a_20992_13103# cal_lut\[18\] a_20417_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X400 _0322_ a_6555_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X401 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_5264_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X402 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X403 vccd1 ctr\[5\] a_5077_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X404 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X405 a_20161_22351# _0064_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X406 a_5897_28335# a_5661_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X407 a_23167_26935# a_23263_26935# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X408 a_7073_25589# _0733_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X409 _0194_ _0383_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X410 vssd1 a_18723_3579# a_18681_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X411 a_1741_30199# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X412 vccd1 _0443_ a_19287_21835# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X413 _0293_ a_16996_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X414 vssd1 a_16734_27359# a_16692_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X415 vccd1 net2 a_3155_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X416 vccd1 a_8268_24501# _0722_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X417 vssd1 _0434_ a_6705_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.266 pd=2.12 as=0.091 ps=0.93 w=0.65 l=0.15
X420 a_10570_7093# a_10402_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X421 a_23707_8029# a_23009_7663# a_23450_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X424 a_27847_7119# a_27149_7125# a_27590_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X425 vssd1 _0624_ a_16373_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X426 vssd1 a_4866_5599# a_4824_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X427 a_7308_10761# a_6909_10389# a_7182_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X428 a_16807_11293# a_16109_10927# a_16550_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X429 a_12525_3855# _0130_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X430 vccd1 _0463_ a_22457_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X431 a_5971_15253# ctr\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X432 a_10033_6409# a_9043_6037# a_9907_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X434 vccd1 _0722_ a_7079_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X435 a_4892_20175# _0759_ a_4719_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X436 a_23959_20553# a_23823_20393# a_23539_20407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 cal_lut\[79\] a_9155_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X439 vccd1 _0441_ a_12539_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X440 vccd1 cal_lut\[29\] a_19303_16519# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X441 a_11796_30511# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X442 _0245_ a_25047_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X443 a_8025_21263# _0755_ _0794_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X444 a_5639_16911# clknet_1_0__leaf__0380_ _0381_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X445 a_2317_27497# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X447 vccd1 _0755_ a_5547_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X448 vccd1 a_17682_16100# a_17611_16201# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X449 vccd1 a_17095_10004# _0106_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X450 vssd1 cal_lut\[189\] a_5173_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X451 vssd1 a_19681_12161# _0525_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X452 vssd1 a_10659_3829# _0314_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X453 vccd1 dec1.i_ones _0720_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X455 vccd1 _0873_ a_19991_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X456 a_19609_10927# _0102_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X457 vccd1 _0462_ a_21983_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X458 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X459 vccd1 a_15722_12533# a_15649_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X460 vssd1 _0425_ a_13091_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X461 vccd1 a_8987_14735# a_9155_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X463 vssd1 a_1461_21781# _0763_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X464 vccd1 a_18698_19319# _0461_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X465 a_18979_21376# cal_lut\[64\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X466 a_17710_15529# _0552_ a_17630_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X467 vssd1 a_27215_13879# cal_lut\[174\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X468 a_20338_1679# a_19899_1685# a_20253_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X469 net68 clknet_1_0__leaf_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X470 a_18689_13647# _0011_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X472 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X474 a_20937_18365# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X476 vccd1 _0141_ a_4413_7497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X477 _0505_ a_17323_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X478 a_5123_5853# a_4425_5487# a_4866_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X479 a_12310_10615# _0659_ a_12613_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X481 a_10659_25321# _0718_ a_10197_25223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X482 vssd1 a_14151_4564# _0131_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X483 a_22269_11791# cal_lut\[157\] a_21831_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X484 _0262_ a_20907_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X485 vccd1 a_13052_15797# _0519_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X486 a_11711_11471# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X487 a_4087_21263# _0781_ a_3885_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X488 a_10773_5487# a_10607_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X489 vccd1 _0561_ a_13341_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X490 cal_lut\[2\] a_8419_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X491 vccd1 a_7067_5162# _0135_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X492 a_20705_9673# a_19715_9301# a_20579_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X493 vssd1 net41 a_15023_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X494 vssd1 _0353_ a_27259_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X495 a_25014_8863# a_24846_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X496 vccd1 a_24099_4073# a_24106_3977# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X497 a_4163_8029# a_3983_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X498 cal_lut\[70\] a_26267_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X499 a_10659_3829# a_10835_4161# a_10787_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X500 vssd1 _0482_ a_15829_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X501 a_28149_14025# a_27595_13865# a_27802_13924# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X503 vccd1 cal_lut\[63\] a_23351_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X504 a_12649_11293# a_12311_11079# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X505 a_9043_11177# _0496_ a_9126_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X506 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4351_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X507 vssd1 a_15623_26324# _0045_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X509 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X510 vssd1 a_26467_10205# a_26635_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X511 vccd1 _0754_ a_3891_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X512 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X513 a_16117_15279# _0454_ a_16035_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X515 vssd1 _0460_ _0590_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X516 a_22988_4917# _0478_ a_23117_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X517 a_16731_1653# cal_lut\[149\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X518 vssd1 a_13514_21237# a_13472_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X519 a_15101_13647# _0010_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X520 a_13161_14191# a_12171_14191# a_13035_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X521 a_16991_27613# a_16127_27247# a_16734_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X522 vssd1 a_18107_7338# _0112_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X523 a_5507_22325# _0747_ a_5725_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X525 a_14616_14709# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X526 a_17930_1653# a_17762_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X527 a_17680_10703# cal_lut\[107\] a_17105_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X528 a_7093_27247# a_6927_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X529 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X530 vccd1 _0422_ a_3785_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X531 a_7323_14735# a_6541_14741# a_7239_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X532 vccd1 a_21897_12533# _0683_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X533 vssd1 a_15354_13621# a_15312_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X534 vccd1 a_5326_6005# a_5253_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X535 vccd1 a_21879_6250# _0157_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X536 vssd1 a_23443_20407# cal_lut\[58\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X537 vssd1 a_24519_14709# a_24477_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X538 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X539 a_5173_10927# a_4903_11293# a_5083_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X540 vssd1 a_14523_6549# _0307_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X541 vssd1 _0216_ a_17459_29185# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X542 vssd1 _0433_ _0435_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X543 vccd1 _0418_ a_1917_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X544 vccd1 net35 a_19715_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X545 vccd1 _0531_ a_15023_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X546 a_13771_21263# a_13073_21269# a_13514_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X547 a_16661_27613# a_16127_27247# a_16566_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X548 vssd1 a_19255_19631# _0462_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X549 vccd1 a_20867_2986# _0153_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X550 a_13606_12533# a_13438_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X551 vccd1 net30 a_12171_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X552 vccd1 a_14307_4917# a_14223_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X554 vssd1 a_19793_21959# _0240_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X555 vccd1 ctr\[1\] a_2695_14013# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0746 ps=0.775 w=0.42 l=0.15
X558 a_16761_26703# _0484_ a_16845_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X559 _0694_ a_9963_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X560 vssd1 a_22431_13866# _0013_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X561 a_23915_17129# net42 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X562 a_24972_7497# a_24573_7125# a_24846_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X564 vssd1 a_8419_29691# a_8377_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X566 vssd1 a_8175_11445# _0881_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X567 vccd1 a_17555_19319# _0580_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X568 vccd1 _0266_ a_17875_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X569 a_6814_12381# a_6375_12015# a_6729_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X571 vssd1 _0462_ a_20329_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X572 a_8951_6825# _0498_ a_9034_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X573 vssd1 _0455_ a_16311_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X574 a_11422_20969# _0676_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X575 a_14833_18115# dbg_result[1] a_14737_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X576 a_8533_22671# _0774_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X577 vccd1 clknet_0_net67 a_3869_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X578 _0211_ _0407_ a_9037_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.127 ps=1.25 w=1 l=0.15
X579 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X580 vssd1 a_24030_20452# a_23959_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X581 a_12437_22671# _0665_ _0707_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X582 a_13438_12559# a_13165_12565# a_13353_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X583 a_11508_20719# a_10975_20969# _0679_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 _0759_ a_3995_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X585 _0840_ a_6647_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X586 vssd1 a_5324_4373# net23 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X587 cal_lut\[55\] a_22863_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X588 vccd1 a_4491_13879# _0809_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X589 a_21081_2223# _0153_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X591 _0147_ a_11711_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X592 vccd1 a_22339_27399# cal_lut\[56\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X594 a_21155_26133# net45 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X595 a_24262_10383# cal_lut\[169\] a_24105_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X596 vccd1 _0237_ a_24867_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X597 a_7231_3677# a_6449_3311# a_7147_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X598 a_19100_22351# _0618_ a_18998_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X599 vccd1 a_17783_21271# _0531_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X600 a_24964_9839# _0510_ a_24473_9813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X601 vccd1 _0863_ a_24591_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X602 a_22983_15431# _0531_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X603 vssd1 a_11794_8725# a_11723_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X604 a_11303_8725# a_11594_9025# a_11545_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X605 a_13172_7663# cal_lut\[124\] a_12597_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X606 cal_lut\[149\] a_15135_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X607 a_13422_9269# a_13254_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X608 vssd1 a_20119_11293# a_20287_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X610 vccd1 _0236_ a_23671_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X611 a_12962_27359# a_12794_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X612 a_11632_15279# a_11233_15279# a_11506_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X613 cal_lut\[107\] a_17711_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X614 a_9305_1135# _0181_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X615 vssd1 a_15727_21959# _0484_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X616 a_20400_15939# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X617 a_17313_14191# _0454_ a_17231_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X618 vssd1 a_3072_19637# _0747_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X619 a_20893_2223# a_20727_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X620 a_22891_20871# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X621 vccd1 a_9563_28487# _0406_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X622 vccd1 net16 a_12455_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X623 vccd1 a_10827_3677# a_10995_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X624 a_7912_31055# a_7663_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X625 vssd1 a_5416_23413# _0821_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X626 a_20069_7663# _0110_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X627 a_5507_22325# _0788_ a_5938_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X628 vccd1 _0352_ a_27167_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X630 vccd1 net45 a_17323_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X631 a_10777_27247# _0196_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X632 a_22469_22895# cal_lut\[85\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X633 vssd1 a_11579_3829# _0363_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X634 _0192_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X635 _0857_ a_23759_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X636 vssd1 a_2014_12533# a_1972_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X637 a_14177_3855# a_13643_3861# a_14082_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X638 a_25875_13647# a_25695_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X639 cal_lut\[76\] a_27003_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X642 _0688_ a_21889_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.172 ps=1.35 w=1 l=0.15
X643 vccd1 a_19862_28447# a_19789_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X644 vccd1 a_11029_17429# _0663_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X645 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X646 vssd1 _0838_ a_1945_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X647 a_20464_2057# a_20065_1685# a_20338_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X650 vssd1 a_9319_26159# a_9767_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0683 ps=0.745 w=0.42 l=0.15
X651 a_10883_25071# _0729_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.219 ps=1.33 w=0.65 l=0.15
X652 a_19303_23047# _0465_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X653 _0250_ a_27024_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X654 a_7550_14557# a_7277_14191# a_7465_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X655 a_22365_3861# a_22199_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X656 a_14741_6397# a_14471_6031# a_14651_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X657 _0300_ a_13040_6147# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X658 a_21626_6941# a_21187_6575# a_21541_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X659 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2879_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X661 a_12318_26677# a_12150_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X662 vssd1 a_2288_17973# _0420_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X663 a_19793_26703# _0052_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X664 _0446_ a_12815_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X665 a_22150_12879# cal_lut\[175\] a_22060_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X666 a_10793_19203# _0626_ a_10697_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X667 vssd1 _0817_ _0826_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X668 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X669 vccd1 a_12559_7093# a_12475_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X670 vssd1 _0277_ a_12263_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X671 a_22596_10383# _0632_ a_22494_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X672 a_2009_30676# _0831_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X673 vssd1 net9 a_12163_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X674 a_12625_4399# a_12355_4765# a_12535_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X675 vssd1 a_12955_25834# _0008_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X676 vssd1 cal_lut\[148\] a_13729_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X677 a_20359_20719# cal_lut\[54\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X678 vccd1 _0320_ a_4443_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X679 a_4140_31055# a_3891_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X680 a_11067_6941# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X681 a_15496_17455# a_15097_17455# a_15370_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X682 vssd1 a_7147_3677# a_7315_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X683 vssd1 _0306_ a_13183_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X685 vccd1 _0422_ a_3238_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0567 ps=0.69 w=0.42 l=0.15
X686 a_17651_8181# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X687 vccd1 _0706_ a_11882_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X688 _0843_ a_9223_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X689 _0290_ a_17875_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X690 a_22787_14735# a_22089_14741# a_22530_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X691 cal_lut\[131\] a_13203_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X692 a_4406_9951# a_4238_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X693 a_5253_6031# a_4719_6037# a_5158_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X694 a_6879_6549# _0316_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X695 a_13438_12559# a_12999_12565# a_13353_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X696 a_10347_25071# _0731_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X697 _0413_ a_1773_22467# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X698 _0113_ a_18887_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X699 a_6729_7119# _0143_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X700 vccd1 cal_lut\[99\] a_12259_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X701 a_14151_11079# _0440_ a_14385_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X702 a_8390_23439# clknet_0__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X704 _0815_ a_7847_28992# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X705 vssd1 a_22971_13469# a_23139_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X706 _0419_ _0414_ a_2695_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 vccd1 a_20775_5639# _0585_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X708 vssd1 _0409_ _0410_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X709 a_5837_23983# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X710 vssd1 cal_lut\[73\] a_27024_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X711 a_20690_3423# a_20522_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X712 a_17589_5487# _0445_ a_17507_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X713 vccd1 _0476_ a_9963_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X714 cal_lut\[47\] a_18355_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X715 vccd1 a_2839_27221# _0831_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X716 a_5460_17999# clknet_1_0__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X717 vssd1 _0754_ a_3891_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X718 vssd1 _0838_ a_13459_22359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X719 a_9928_6825# cal_lut\[127\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X720 a_18942_13621# a_18774_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X722 vccd1 _0763_ a_1959_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X723 vssd1 cal_lut\[173\] a_27621_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X724 vssd1 cal_lut\[93\] a_14373_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X725 vccd1 _0671_ _0707_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X727 vssd1 _0420_ a_3615_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X728 a_9899_1501# a_9117_1135# a_9815_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X729 vccd1 cal_lut\[170\] a_27163_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X730 vccd1 a_16734_27359# a_16661_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X731 vssd1 net44 a_16863_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X732 a_10844_31029# net9 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X733 a_23903_27069# a_23683_27081# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X734 net22 a_2747_18517# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X736 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X737 a_9643_21046# _0626_ a_9184_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X738 vccd1 a_7994_8863# a_7921_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X739 a_7952_10927# a_7553_10927# a_7826_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X740 a_23391_22351# a_23211_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X741 a_6245_21781# _0431_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X742 _0233_ a_21872_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X744 _0730_ _0711_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X745 _0434_ net7 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X746 a_17811_2589# a_17029_2223# a_17727_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X748 vccd1 a_5567_7931# a_5483_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X749 _0352_ a_24683_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X750 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9496_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X752 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd _0784_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X753 vccd1 _0414_ a_2485_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X754 a_27333_15829# a_27167_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X755 vssd1 _0850_ a_24407_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X756 a_10784_23983# _0681_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X757 a_6537_19605# clknet_0__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X758 vssd1 a_10699_4399# _0850_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X759 a_12893_25071# _0008_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X760 a_19915_19087# a_19715_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X761 vccd1 cal_lut\[31\] a_23391_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X762 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10028_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X764 vssd1 a_14345_9269# _0565_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X765 a_18843_13131# net80 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X766 a_20690_21237# a_20522_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X767 net32 a_17783_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X768 a_12778_14303# a_12610_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X769 a_6633_26703# a_6397_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X770 a_12843_17821# a_12061_17455# a_12759_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X771 a_13129_16911# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X772 a_3969_12559# _0203_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X773 a_14821_23445# a_14655_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X774 a_4709_19881# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X775 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd a_9687_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X776 vssd1 _0495_ a_16281_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X777 _0123_ a_11527_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X778 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X779 a_27461_15645# a_27123_15431# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X780 vssd1 a_13035_14557# a_13203_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X781 a_19878_28879# a_19439_28885# a_19793_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X782 vssd1 cal_lut\[69\] a_25137_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X783 vccd1 a_17743_2741# _0339_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X784 ctr\[2\] a_2947_10615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X785 vssd1 a_19126_16885# a_19084_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X786 vssd1 cal_lut\[126\] a_7980_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X787 vccd1 a_6487_11195# a_6403_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X788 vccd1 a_6445_29111# net79 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X789 a_13291_18543# _0438_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X790 a_22861_2767# a_22523_2999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X791 vccd1 a_18119_7637# a_18126_7937# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X792 vccd1 a_27491_11092# _0171_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X793 a_10938_28471# a_10779_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X794 a_1471_19319# _0422_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X795 a_2125_15829# a_1959_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X796 a_25695_13647# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X797 vssd1 _0746_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X798 _0082_ a_17323_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X799 a_10129_9295# cal_lut\[121\] a_10045_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X800 vccd1 a_21591_11293# a_21759_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X802 a_7618_26935# ctr\[10\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X803 a_7753_26819# ctr\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X804 a_25187_15041# _0237_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X806 vccd1 a_21851_14459# a_21767_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X807 a_11046_14557# a_10773_14191# a_10961_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X808 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X809 a_9311_30761# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X810 a_2797_21583# _0770_ a_2701_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X811 a_21181_11791# cal_lut\[104\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X812 vssd1 net40 a_12355_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X813 vccd1 a_18187_1679# a_18355_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X814 vssd1 _0714_ a_9431_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X815 a_23579_16733# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X816 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7912_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X817 temp_delay_last a_2991_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X818 vssd1 _0414_ _0784_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X819 vccd1 ctr\[8\] a_5081_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X820 vccd1 dbg_result[1] a_14103_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X821 vssd1 clknet_1_0__leaf__0380_ a_4733_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X822 vssd1 _0515_ a_13512_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X823 a_9117_13353# cal_lut\[80\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X825 _0446_ a_12815_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X826 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X827 a_6244_25045# _0805_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X828 _0481_ a_12263_20495# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X829 _0485_ _0438_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X830 cal_lut\[127\] a_8419_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X831 a_14373_25071# a_14103_25437# a_14283_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X832 _0556_ net4 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X833 vssd1 a_8971_1653# a_8929_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X834 vssd1 a_1735_27765# _0825_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X835 a_21362_26133# a_21162_26433# a_21511_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X836 a_14733_5487# _0119_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X837 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X838 a_8979_18543# _0439_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X839 vccd1 a_5751_14709# ctr\[6\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X840 vssd1 a_11207_14954# _0004_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X841 vssd1 a_23063_3855# a_23231_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X842 a_25230_21807# a_24915_21959# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X843 a_19820_10927# a_19421_10927# a_19694_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X844 a_21334_9951# a_21166_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X845 vssd1 net8 a_11619_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X846 cal_lut\[90\] a_20287_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X847 a_2309_14191# a_2143_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X848 a_28157_12937# a_27167_12565# a_28031_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X849 a_2409_7663# net63 temp1.capload\[8\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X850 a_10827_7119# a_9963_7125# a_10570_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X851 a_3335_12559# _0390_ a_3117_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X853 vssd1 a_12962_27359# a_12920_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X854 a_5621_10927# a_5455_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X855 vssd1 net40 a_14931_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X856 vccd1 _0876_ a_24591_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X857 a_15972_10089# _0547_ a_15870_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X858 a_4726_24566# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X859 a_12851_2589# a_11987_2223# a_12594_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X860 a_4613_5487# _0136_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X861 a_5377_18319# clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X862 a_23407_17705# cal_lut\[74\] a_23205_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X863 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4140_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X864 _0220_ a_16904_25321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X865 vccd1 a_26819_6843# a_26735_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X866 a_21752_6575# a_21353_6575# a_21626_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X867 a_18119_7637# net32 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X868 a_5250_9295# a_4811_9301# a_5165_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X869 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8300_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X870 a_6463_22057# _0755_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X871 vssd1 net41 a_12907_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X875 vssd1 cal_lut\[101\] a_15524_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X876 vssd1 a_6699_13268# _0018_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X877 a_17762_25437# a_17489_25071# a_17677_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X878 vccd1 _0759_ a_4283_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X879 vssd1 _0756_ _0757_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X880 vssd1 a_20690_21237# a_20648_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X882 vccd1 a_9096_27221# _0817_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X883 vssd1 _0787_ a_7021_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X884 a_14604_20969# _0872_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X885 vssd1 net29 a_14747_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X886 vccd1 cal_lut\[156\] a_18383_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X887 a_11049_10499# _0696_ a_10977_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X888 a_11303_8725# a_11587_8725# a_11522_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X889 vccd1 a_5871_10004# _0138_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X890 vccd1 a_23351_21959# _0638_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X892 a_13679_9295# a_12981_9301# a_13422_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X893 vssd1 a_19827_25589# a_19785_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X894 a_21936_16367# a_21537_16367# a_21810_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X895 a_15371_15823# _0550_ a_15289_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X896 a_21029_6369# _0441_ a_20943_6369# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X897 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X898 vccd1 cal_lut\[25\] a_23021_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X899 vssd1 a_21879_6250# _0157_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X900 vssd1 _0447_ _0485_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X901 a_10137_17705# net12 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X902 vssd1 _0206_ a_6437_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X903 vssd1 a_11759_4564# _0129_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X904 vssd1 a_6729_30199# _0404_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X905 vssd1 _0507_ a_18397_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X906 a_7921_9117# a_7387_8751# a_7826_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X907 net2 a_1407_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X908 vccd1 net34 a_25419_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X909 a_20947_21263# a_20249_21269# a_20690_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X910 a_27606_17821# a_27333_17455# a_27521_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X911 a_16116_9839# cal_lut\[102\] a_15541_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X912 cal_lut\[191\] a_7407_12283# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X913 a_4277_23957# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X914 vccd1 cal_lut\[73\] a_27106_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X915 vccd1 a_22955_14709# a_22871_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R2 vccd1 temp1.capload\[2\].cap_57.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X917 _0855_ a_21735_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X918 a_27521_12559# _0172_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X919 a_21975_19605# a_22266_19905# a_22217_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X920 a_4406_8863# a_4238_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X921 _0755_ a_3891_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X922 a_3424_30287# temp1.dac.vdac_single.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X923 a_13955_23439# a_13091_23445# a_13698_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X925 vssd1 _0111_ a_18673_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X926 vssd1 _0474_ a_22961_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X927 a_2503_31375# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X928 a_20663_8029# a_19881_7663# a_20579_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X929 vssd1 _0422_ a_3799_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.109 ps=1.36 w=0.42 l=0.15
X931 _0214_ a_16076_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X932 vssd1 a_9765_6727# _0309_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X933 a_27337_7119# _0162_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X934 vccd1 net76 _0399_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X937 a_9899_14557# a_9117_14191# a_9815_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X938 vccd1 a_2439_12533# a_2355_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X939 a_22898_6005# a_22730_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X940 vccd1 clknet_1_0__leaf_io_in[0] a_3615_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X941 a_5541_3311# a_5271_3677# a_5451_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X942 _0088_ a_17231_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X943 vssd1 net67 a_3882_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X945 vssd1 clknet_0__0380_ a_8390_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X947 net18 a_14287_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X948 a_17168_13647# _0487_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X949 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X950 _0213_ a_14604_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X951 vssd1 a_25755_20393# a_25762_20297# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X952 vssd1 a_3859_7337# a_3866_7241# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X953 a_17893_27791# a_17555_28023# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X954 a_18371_26525# a_17673_26159# a_18114_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X955 vssd1 a_26743_16733# a_26911_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X956 a_16731_1653# a_16907_1985# a_16859_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X957 vccd1 _0863_ a_8767_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X959 a_20470_6031# _0584_ a_20390_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X961 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X964 vssd1 a_22903_21959# _0463_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X965 net39 a_3155_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X967 a_3236_15055# _0393_ a_2933_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X968 vccd1 a_9360_30663# a_9311_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X969 vssd1 a_5675_3855# a_5843_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X970 vccd1 _0258_ a_12723_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X971 _0509_ a_23151_10955# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X972 a_10028_31849# a_9779_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X973 a_24551_19605# a_24842_19905# a_24793_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X974 vccd1 cal_lut\[126\] a_8062_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X975 vssd1 clknet_1_0__leaf_io_in[0] a_1407_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X976 a_11874_3677# a_11601_3311# a_11789_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X977 a_10851_11079# _0460_ a_11025_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X978 vssd1 a_7994_8863# a_7952_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X979 a_13253_13103# a_12263_13103# a_13127_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X980 vssd1 _0737_ _0795_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X981 a_12889_27613# a_12355_27247# a_12794_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X982 vccd1 a_5644_12533# a_5404_12797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.41 as=0.217 ps=2.17 w=0.82 l=0.25
X983 a_13892_19407# a_13838_19319# a_13796_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X984 vssd1 _0598_ a_16737_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X985 vssd1 a_17095_5639# _0614_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X986 vssd1 a_6703_6549# _0327_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X987 a_6081_8751# a_5915_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X988 net74 a_6003_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X989 vssd1 _0803_ a_2959_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
X990 _0267_ a_17135_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X992 a_15473_27497# _0484_ a_15557_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X993 a_13508_18517# dbg_result[1] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X994 vssd1 _0451_ a_23763_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X995 vssd1 a_27774_11445# a_27732_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X996 vssd1 a_7959_27515# a_7917_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X997 a_8303_16911# a_8123_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X998 vccd1 _0495_ a_15667_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X999 a_2805_19407# _0418_ a_2709_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1001 vccd1 a_18669_22325# _0621_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1002 a_23683_10383# cal_lut\[67\] a_23481_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1004 _0651_ a_10699_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1005 vccd1 net42 a_24591_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1007 a_22695_27791# a_21997_27797# a_22438_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1008 a_4584_24759# dbg_result[5] a_4726_24566# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1009 vccd1 cal_lut\[27\] a_24863_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1010 vccd1 clknet_1_0__leaf_io_in[0] a_4719_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1011 a_20175_5056# cal_lut\[154\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1012 a_6256_31849# a_6007_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1013 a_22438_23413# a_22270_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1014 vccd1 net1 a_2235_9303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1015 a_17286_9269# a_17118_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1016 a_27548_18377# a_27149_18005# a_27422_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1017 vssd1 _0320_ a_4443_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1019 vssd1 cal_lut\[53\] a_20308_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1020 vccd1 _0422_ a_3785_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1021 a_23811_15431# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1023 vccd1 _0452_ a_16127_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1024 vccd1 _0288_ a_21371_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1025 vssd1 _0835_ a_6835_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1026 vssd1 _0236_ a_23671_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1027 vccd1 cal_lut\[156\] a_19435_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1028 a_8543_30485# temp1.dac.parallel_cells\[4\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1029 vccd1 _0817_ a_2317_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1032 a_23811_15431# _0460_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1033 vssd1 _0027_ a_25389_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1035 a_11693_8207# cal_lut\[99\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1036 a_11233_15279# a_11067_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1037 _0113_ a_18887_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1038 vccd1 a_10659_7637# net26 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1039 _0103_ a_20175_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1041 vccd1 _0418_ a_5555_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1042 vssd1 a_21794_6687# a_21752_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1043 vssd1 a_27583_9514# _0170_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1044 a_2024_27497# a_1775_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1045 a_5376_9673# a_4977_9301# a_5250_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1046 a_7929_29245# ctr\[10\] a_7847_28992# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1047 a_26225_17455# a_25235_17455# a_26099_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1048 a_5621_10927# a_5455_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1049 vccd1 a_10809_19605# a_10839_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1050 _0442_ a_14523_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1051 vssd1 a_9447_8207# a_9615_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1052 a_22633_11445# _0456_ a_22790_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1053 vccd1 a_25271_23261# a_25439_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1054 vccd1 io_in[5] a_1407_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1055 a_14633_16201# a_13643_15829# a_14507_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1056 a_8101_14191# a_7111_14191# a_7975_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1057 a_5123_5853# a_4259_5487# a_4866_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1058 a_17003_7691# net17 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1059 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1061 a_4679_19319# net21 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1062 vssd1 a_27491_17130# _0073_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1063 vccd1 a_18475_5639# _0615_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1064 a_19225_11837# cal_lut\[186\] a_19153_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1065 _0849_ a_13363_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X1067 a_27149_7125# a_26983_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1069 vccd1 cal_lut\[123\] a_11247_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1070 a_18698_19319# a_19167_19061# a_19111_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X1071 vccd1 cal_lut\[63\] a_25415_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1072 a_7093_27247# a_6927_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1073 a_7439_4373# net1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1074 a_8013_4949# a_7847_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1075 vssd1 a_11527_9303# net29 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1076 vssd1 a_19333_13255# _0860_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1077 vccd1 net28 a_7111_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1078 a_8263_15444# _0255_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1079 cal_lut\[127\] a_8419_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1080 net78 a_8671_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1082 a_23027_12559# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1083 a_20893_25071# a_20727_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1084 vssd1 a_2376_30199# _0833_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1085 a_5341_17429# clknet_0_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1086 vccd1 _0268_ a_18979_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1087 vccd1 a_15711_24833# a_15535_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1088 a_17325_20291# _0578_ a_17229_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1089 vssd1 _0475_ a_23200_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1090 a_8653_4233# a_7663_3861# a_8527_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1091 a_6460_26159# _0400_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1092 vccd1 a_14747_20175# net20 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1093 vccd1 a_6979_19061# _0383_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X1094 a_21997_23445# a_21831_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1095 vssd1 _0468_ a_17772_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1096 a_9559_26481# ctr\[7\] a_9487_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0578 ps=0.695 w=0.42 l=0.15
X1097 vssd1 _0394_ a_3236_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1098 a_15097_17455# a_14931_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1099 _0294_ a_18515_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X1101 a_16189_15279# cal_lut\[35\] a_16117_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1102 a_25271_9117# a_24407_8751# a_25014_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1103 a_20203_11293# a_19421_10927# a_20119_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1104 a_27521_11471# _0171_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1105 a_8979_18543# _0520_ _0680_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1107 a_16845_9301# a_16679_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1108 a_5547_26409# ctr\[8\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1111 a_14283_3311# cal_lut\[131\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X1112 a_8758_10383# _0496_ a_8758_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X1113 _0089_ a_18979_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1114 a_15956_25071# a_15557_25071# a_15830_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1115 vccd1 a_14243_16532# _0035_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1116 a_4977_9301# a_4811_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1117 vccd1 a_10851_11079# _0496_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1118 a_27333_12565# a_27167_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1119 a_14103_18793# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1121 vccd1 a_14967_8029# a_15135_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1122 a_11797_25071# _0708_ a_11579_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1123 vccd1 a_6516_20871# _0736_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1124 a_5324_4373# net39 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1125 a_6459_32143# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1126 vssd1 net31 a_19255_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1127 a_17578_6941# a_17305_6575# a_17493_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1128 a_19681_12161# _0522_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1129 a_6644_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1130 a_11224_29967# a_10975_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1131 a_21155_26133# net45 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1132 vccd1 a_15979_3855# a_16147_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1133 vssd1 _0486_ a_14449_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1134 a_20298_22057# _0222_ a_20216_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1136 a_13809_15829# a_13643_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1137 a_1941_14735# a_1407_14741# a_1846_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1138 vssd1 cal_lut\[183\] a_11797_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1139 a_24846_7119# a_24573_7125# a_24761_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1140 a_24573_25071# a_24407_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1141 vssd1 _0384_ _0195_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1142 vssd1 cal_lut\[184\] a_13913_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1144 vccd1 _0841_ a_8951_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1145 a_22903_2985# net33 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1146 a_7365_12937# a_6375_12565# a_7239_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1147 a_16189_6397# cal_lut\[119\] a_16117_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1148 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1149 vssd1 a_22503_24135# _0685_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1150 a_23513_21807# _0443_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1151 _0650_ a_11527_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1152 vccd1 a_10239_31055# net14 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1154 a_3479_7351# a_3575_7351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1155 _0286_ a_16168_9411# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1156 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1157 _0398_ _0809_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1159 a_13838_19319# _0442_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1160 vccd1 _0380_ a_7102_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1161 a_2116_29673# a_1867_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1163 _0495_ a_13714_19407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X1164 a_20249_3311# a_20083_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1166 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1167 vccd1 _0862_ a_9595_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1168 a_5250_13469# a_4977_13103# a_5165_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1169 a_19987_13353# _0534_ a_19881_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.19 ps=1.38 w=1 l=0.15
X1170 vccd1 a_2377_28500# temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1171 a_16339_25437# a_15557_25071# a_16255_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1172 a_11471_14557# a_10773_14191# a_11214_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1173 vssd1 _0628_ _0716_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1174 a_24298_16911# a_24051_17289# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1176 vccd1 cal_lut\[110\] a_19619_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1177 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1178 a_1741_30199# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1179 a_4091_15529# net68 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X1180 vccd1 a_7410_14709# dbg_result[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X1181 vssd1 _0174_ a_26861_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1182 a_20114_10499# _0260_ a_20032_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1183 ctr\[5\] a_5843_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1184 vccd1 cal_lut\[82\] a_16951_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1185 _0418_ a_2327_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1186 a_15611_13647# a_14913_13653# a_15354_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1188 vssd1 a_15611_1679# a_15779_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1189 vccd1 a_23155_6031# a_23323_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1190 a_23056_17999# _0640_ a_22954_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1191 a_26059_8751# cal_lut\[165\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X1192 a_9853_13103# a_9687_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1193 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6256_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1194 vssd1 a_23547_26921# a_23554_26825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1195 vccd1 a_2931_22325# _0783_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1197 vssd1 a_21223_19997# a_21391_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 a_25713_20175# a_25375_20407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1199 vccd1 _0309_ a_8767_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1200 a_17078_7235# _0283_ a_16996_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1201 a_14116_27081# a_13717_26709# a_13990_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1202 a_18114_26271# a_17946_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1203 vccd1 _0720_ a_6619_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1204 vccd1 _0451_ a_22843_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1205 vccd1 a_2000_26935# a_1951_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1207 vssd1 _0495_ a_12693_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1208 vssd1 a_23167_26935# cal_lut\[57\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1209 vccd1 a_8251_9117# a_8419_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1210 vssd1 a_27491_11092# _0171_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1211 vssd1 a_19439_21263# _0459_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1214 a_9499_3133# cal_lut\[180\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X1215 a_17385_14191# cal_lut\[23\] a_17313_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1216 _0476_ a_23763_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1217 a_15439_2388# _0366_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1218 _0703_ a_9749_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.373 ps=1.75 w=1 l=0.15
X1219 vssd1 _0838_ a_13459_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1220 vssd1 a_8987_14735# a_9155_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1221 vccd1 a_10995_7093# a_10911_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1222 vssd1 a_13127_13469# a_13295_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1223 vssd1 _0260_ a_19333_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1224 a_5099_20969# _0769_ a_4897_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1225 a_17543_14735# a_16845_14741# a_17286_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1226 a_24094_14709# a_23926_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1227 a_11214_5599# a_11046_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1228 vssd1 io_in[3] a_1407_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1229 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1230 vccd1 clknet_0_temp1.i_precharge_n a_1753_26133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1231 _0428_ _0411_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1233 vccd1 cal_lut\[3\] a_9223_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1235 a_25014_8863# a_24846_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1236 vssd1 a_17286_9269# a_17244_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1237 a_23197_7663# _0109_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1238 a_7097_10383# _0187_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1239 a_7826_13469# a_7553_13103# a_7741_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1240 vssd1 _0653_ a_11527_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1241 vccd1 _0266_ a_17691_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1243 net2 a_1407_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1244 a_23351_8439# _0450_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1245 _0028_ a_18611_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1246 a_25007_5175# a_25103_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1247 a_11214_5599# a_11046_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1248 dbg_result[3] a_7410_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X1249 vssd1 a_21759_11195# a_21717_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1250 vccd1 net32 a_19255_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1252 _0530_ a_15299_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1253 cal_lut\[83\] a_18355_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1254 a_15695_1679# a_14913_1685# a_15611_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1255 a_5271_10205# _0836_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1256 vssd1 net1 a_3155_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1257 a_17647_29423# a_17427_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1258 a_26946_21919# a_26778_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1263 a_18313_25071# a_17323_25071# a_18187_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1264 a_22619_2999# a_22903_2985# a_22838_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1265 vssd1 a_25143_6031# _0341_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1266 a_18671_9513# net35 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1268 a_9591_1679# a_9411_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1269 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1270 vssd1 _0872_ a_14733_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1271 a_8297_20765# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1272 a_19167_19061# dbg_result[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X1273 vccd1 a_27847_17999# a_28015_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1274 a_2947_10615# a_3115_10615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1275 a_10865_19203# _0589_ a_10793_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1276 a_17397_2589# a_16863_2223# a_17302_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1277 _0346_ a_25783_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X1279 _0114_ a_20727_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1281 vssd1 temp1.i_precharge_n a_2778_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1282 a_3885_21263# _0780_ a_4087_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1283 a_14457_1135# _0148_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1284 vssd1 a_2023_19319# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X1285 vccd1 a_3175_14459# ctr\[3\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1286 a_6791_4074# _0315_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1287 a_13035_3855# a_12171_3861# a_12778_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1289 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1290 vssd1 a_26578_18655# a_26536_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1291 a_25842_17567# a_25674_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1292 vccd1 a_8251_16733# a_8419_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1293 vssd1 a_9983_1403# a_9941_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1294 a_10677_13103# a_9687_13103# a_10551_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1295 temp1.capload\[9\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1296 _0284_ a_20952_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1297 _0097_ a_12815_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1298 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1299 vssd1 a_26099_17821# a_26267_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1300 a_7718_14303# a_7550_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1301 a_23481_21629# a_23211_21263# a_23391_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X1302 a_20874_27765# a_20706_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1303 a_23282_8029# a_22843_7663# a_23197_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1304 vssd1 a_7975_14557# a_8143_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1305 a_27422_7119# a_26983_7125# a_27337_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1306 a_16925_8751# cal_lut\[125\] a_16853_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1307 a_21537_16367# a_21371_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1308 vssd1 a_13537_15431# _0255_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1310 temp1.dac_vout_notouch_ net13 a_11224_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1311 vccd1 a_15630_19743# a_15557_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1312 vssd1 cal_lut\[76\] a_17225_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1313 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1314 vssd1 _0258_ a_12723_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1315 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1316 vssd1 a_22863_23413# a_22821_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1317 vssd1 _0854_ a_20635_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1318 vccd1 _0773_ a_3749_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1319 vccd1 ctr\[2\] a_2071_11791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X1320 vccd1 cal_lut\[29\] a_19838_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1321 vccd1 _0863_ a_24499_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1322 _0590_ net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1323 vccd1 _0159_ a_25389_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1324 a_4224_30333# _0800_ a_4003_30006# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1325 vssd1 dbg_result[4] _0453_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1326 vccd1 a_10938_28471# a_10872_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X1327 _0067_ a_23671_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1328 a_22741_8751# _0450_ a_22659_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1330 vssd1 a_28199_12533# a_28157_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1331 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1333 a_25773_8207# _0165_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1334 a_23351_8439# _0450_ a_23585_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1335 a_15093_27247# cal_lut\[49\] a_14747_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1336 _0488_ a_14103_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1337 a_20430_16911# a_19991_16917# a_20345_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1338 vssd1 _0731_ a_10883_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.219 pd=1.33 as=0.101 ps=0.96 w=0.65 l=0.15
X1339 io_out[1] a_1551_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1340 _0429_ a_3615_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1341 vssd1 _0683_ a_21831_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1342 vssd1 a_20141_6005# _0586_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X1343 a_18475_7663# a_18255_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1345 a_4484_32375# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1346 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_2116_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1347 a_18348_29257# a_17949_28885# a_18222_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1349 vccd1 _0841_ a_7571_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1352 a_9868_5487# _0451_ a_9678_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X1353 vccd1 a_22988_4917# _0479_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1354 vssd1 _0378_ a_12815_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1355 vccd1 dec1.i_ones a_8055_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X1356 a_3882_22895# clknet_0_temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1357 vssd1 _0508_ a_23549_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1358 a_11422_20969# _0678_ _0679_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1359 _0435_ _0434_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1360 vssd1 a_2419_12015# _0390_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1361 a_5759_9295# a_4977_9301# a_5675_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1362 a_15603_29789# a_14821_29423# a_15519_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1363 a_27774_9951# a_27606_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1364 vssd1 _0058_ a_22813_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1365 vccd1 a_28199_10107# a_28115_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1366 a_19973_22357# a_19807_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1367 vssd1 a_11287_27613# a_11458_27500# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1368 vccd1 cal_lut\[48\] a_19746_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1370 _0148_ a_14103_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1371 a_23117_5263# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X1373 _0644_ a_15023_22464# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1374 vccd1 a_23915_17129# a_23922_17033# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1375 vssd1 a_13606_12533# a_13564_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1377 a_8055_25321# _0713_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X1379 vssd1 a_22806_25183# a_22764_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1380 a_5693_21781# _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1381 a_10843_2197# cal_lut\[186\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X1382 vssd1 a_10379_6740# _0122_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1383 a_21009_5487# cal_lut\[118\] a_20937_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1384 vccd1 _0676_ a_11422_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1385 a_17996_13647# _0475_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1386 _0204_ _0397_ a_4345_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.127 ps=1.25 w=1 l=0.15
X1387 a_15829_3145# a_14839_2773# a_15703_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1388 _0649_ a_10699_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1389 a_7952_29423# a_7553_29423# a_7826_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1390 _0492_ _0491_ a_15959_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1391 vssd1 _0246_ a_13537_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1392 a_15243_5853# a_14545_5487# a_14986_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1394 vccd1 a_8351_11777# a_8175_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1395 vccd1 cal_lut\[146\] a_10051_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1396 vccd1 a_19759_3073# a_19583_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1397 vssd1 cal_lut\[16\] a_14604_13353# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1400 vssd1 _0267_ a_17231_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1401 a_20727_24527# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1402 vssd1 a_22247_9991# _0634_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1403 vccd1 a_21327_24746# _0084_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1404 a_6920_18377# a_6541_18005# a_6823_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X1406 _0303_ a_8164_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1407 a_16737_12533# _0601_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1408 a_6905_29423# a_5915_29423# a_6779_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1409 a_10914_16617# _0519_ a_10832_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1410 vccd1 temp_delay_last a_4351_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X1412 a_8164_8323# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1413 a_24919_10901# a_25203_10901# a_25138_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1414 a_13245_10927# a_12691_10901# a_12898_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1415 vccd1 net44 a_22291_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1416 a_21003_11471# _0449_ a_21181_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1418 a_11799_22057# _0664_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1420 a_23205_17705# _0473_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X1422 vccd1 a_21683_14557# a_21851_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1423 a_17286_9269# a_17118_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1424 a_18998_22351# _0619_ a_18918_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1425 a_15193_2767# _0179_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1426 vssd1 a_14967_8029# a_15135_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1427 a_15009_23439# _0094_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1428 vssd1 _0633_ a_22165_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X1429 vssd1 a_3615_17999# _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1430 a_20407_16519# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1431 a_17225_19453# a_16955_19087# a_17135_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X1432 a_21327_24746# _0262_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1433 a_8251_13469# a_7553_13103# a_7994_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1435 a_5323_4917# cal_lut\[136\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X1437 cal_lut\[64\] a_27371_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1438 a_5894_11293# a_5621_10927# a_5809_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1439 cal_lut\[17\] a_16147_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1441 a_21131_27791# a_20267_27797# a_20874_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1443 ctr\[2\] a_2947_10615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1444 vccd1 _0327_ a_6375_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1445 a_12052_17999# _0576_ a_11950_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X1446 a_24665_15829# a_24499_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1447 a_11214_14303# a_11046_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1448 temp1.capload\[2\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1449 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1451 vccd1 a_17711_14709# a_17627_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1452 cal_lut\[17\] a_16147_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1453 a_19793_28879# _0048_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1454 vssd1 a_5475_29691# a_5433_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1455 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1457 a_6541_12565# a_6375_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1459 a_12610_3855# a_12171_3861# a_12525_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1461 a_10781_8751# _0451_ a_10699_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1462 vssd1 _0735_ a_6929_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1463 vccd1 a_9907_6031# a_10075_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1464 a_11799_22057# _0673_ a_11581_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1465 vccd1 a_18597_13077# _0456_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1466 cal_lut\[146\] a_8879_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1467 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_8951_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1468 _0380_ a_2879_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1469 cal_lut\[69\] a_25531_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1470 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_2327_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1471 vssd1 _0710_ a_11001_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1472 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1473 vssd1 a_12502_17567# a_12460_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1474 vccd1 a_5291_5755# a_5207_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1475 a_20249_8029# a_19715_7663# a_20154_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1476 a_15959_18793# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1477 a_1945_15431# _0428_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X1478 vssd1 a_18555_3677# a_18723_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1479 a_8845_28023# _0406_ a_9008_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1480 _0023_ a_18611_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1481 a_5995_23983# ctr\[5\] _0773_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1483 vccd1 _0744_ a_2605_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1485 a_15630_19743# a_15462_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1486 a_23930_26703# a_23683_27081# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1487 a_26873_22173# a_26339_21807# a_26778_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1488 vccd1 net23 a_8951_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1489 _0420_ a_2288_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1490 vssd1 _0288_ a_21371_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1491 vssd1 cal_lut\[54\] a_21136_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1492 a_5264_28879# _0402_ _0208_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1493 _0826_ _0817_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1494 vssd1 _0560_ a_19426_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X1495 a_21541_6575# _0157_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1496 vccd1 a_6090_27221# a_6019_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1498 a_10043_27069# _0460_ a_9835_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.173 ps=1.25 w=0.42 l=0.15
X1499 a_21725_21807# _0030_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1500 a_2489_17455# _0422_ a_2931_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1501 a_22457_6037# a_22291_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1502 _0876_ a_24679_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1503 _0058_ a_22659_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1504 _0288_ a_20676_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1505 _0845_ a_12856_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1506 a_24455_12925# a_24235_12937# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1507 _0226_ a_16859_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1508 vccd1 a_9671_21495# _0677_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X1509 vccd1 _0810_ a_5179_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1510 a_17930_1653# a_17762_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1511 vccd1 a_2419_12015# _0390_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1512 vccd1 a_27003_18811# a_26919_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1513 _0421_ a_3155_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1516 a_21721_18909# a_21555_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X1517 a_19303_17607# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1518 _0310_ a_10280_5059# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1519 a_23408_7663# a_23009_7663# a_23282_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1520 _0449_ a_17907_10955# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1521 _0402_ _0812_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1522 a_19763_4074# _0298_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1523 a_27548_7497# a_27149_7125# a_27422_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1524 a_12097_23983# a_11896_24233# _0712_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1525 _0410_ _0409_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1526 vssd1 _0495_ a_17109_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1527 vssd1 a_18187_25437# a_18355_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1528 vssd1 _0501_ a_20440_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1529 _0831_ a_2839_27221# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1530 a_17857_1679# a_17323_1685# a_17762_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1531 a_15186_1679# a_14747_1685# a_15101_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1532 vssd1 a_19303_23047# _0619_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1534 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1535 vssd1 a_12985_10615# _0276_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1536 vccd1 a_17746_6687# a_17673_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1537 vssd1 a_3707_9303# net27 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1540 cal_lut\[8\] a_13387_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1541 cal_lut\[70\] a_26267_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1542 vssd1 _0282_ a_20175_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1543 _0431_ a_1773_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1544 a_4663_9117# a_3799_8751# a_4406_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1545 vccd1 net7 _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1546 a_18326_7637# a_18126_7937# a_18475_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1547 vccd1 cal_lut\[108\] a_20758_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1548 vccd1 net40 a_14011_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1549 vssd1 _0808_ _0393_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1550 a_6453_5487# _0135_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1551 a_27330_9117# a_27057_8751# a_27245_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1552 a_7987_9514# _0302_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1553 vccd1 a_20039_18695# _0612_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1554 a_1641_28500# _0825_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1555 vccd1 _0863_ a_23303_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1556 vssd1 net42 a_27167_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1557 vssd1 _0309_ a_8767_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1558 a_16063_12559# a_15281_12565# a_15979_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1559 vccd1 a_17831_24746# _0046_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1560 a_7656_18543# a_7277_18543# a_7559_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X1561 a_17428_18377# a_17029_18005# a_17302_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1563 vccd1 _0360_ a_26063_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1564 vssd1 _0707_ a_10784_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1567 a_13466_18543# a_13091_18543# a_13375_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.064 ps=0.725 w=0.42 l=0.15
X1568 a_18187_1679# a_17489_1685# a_17930_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1569 cal_lut\[52\] a_18815_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1570 vssd1 cal_lut\[109\] a_23804_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
R3 temp1.capload\[5\].cap_60.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1572 a_1846_12559# a_1573_12565# a_1761_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1573 vccd1 _0211_ a_10025_29257# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1574 vssd1 cal_lut\[120\] a_7704_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 vssd1 ctr\[7\] a_6397_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1576 a_12759_17821# a_11895_17455# a_12502_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1577 vssd1 a_11671_2741# _0331_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1578 a_19930_12265# _0524_ a_19681_12161# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X1579 a_10699_8320# cal_lut\[135\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1581 vssd1 cal_lut\[65\] a_20216_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1582 vssd1 _0706_ a_12097_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1583 temp_delay_last a_2991_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1584 a_17812_15529# _0475_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1585 vccd1 a_23231_25339# a_23147_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1586 a_25949_23817# a_24959_23445# a_25823_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1587 a_25447_15823# a_24665_15829# a_25363_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1588 a_4593_8439# net24 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1589 a_15531_24135# _0481_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1590 vssd1 a_15963_17723# a_15921_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1592 a_15554_3855# a_15115_3861# a_15469_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1593 temp1.capload\[3\].cap.Y net58 a_1769_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1594 a_3007_14557# a_2309_14191# a_2750_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1595 a_3782_10383# a_3535_10761# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1596 a_22821_2057# a_21831_1685# a_22695_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1597 _0515_ _0514_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1598 vccd1 a_18647_28879# a_18815_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1599 a_25271_24349# a_24573_23983# a_25014_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1600 a_2505_9839# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1601 a_6737_22351# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X1602 vssd1 a_7067_5162# _0135_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1603 vssd1 a_15335_7119# a_15503_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1604 a_13091_9001# _0573_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1605 a_3755_10749# a_3535_10761# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1606 vccd1 cal_lut\[45\] a_15479_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1607 a_15725_15797# _0542_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1608 a_11233_15279# a_11067_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1609 a_23631_11079# cal_lut\[110\] a_23757_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1610 a_17555_19319# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1611 a_13649_13647# cal_lut\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1612 vccd1 cal_lut\[141\] a_5359_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1613 vccd1 a_13459_21807# _0216_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1614 _0281_ a_18055_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1615 vccd1 a_12863_14954# _0096_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1616 a_9431_25071# _0713_ a_9235_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1617 a_22235_22173# a_21371_21807# a_21978_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1618 vssd1 _0799_ a_4069_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X1619 vssd1 _0222_ a_19793_21959# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1620 vssd1 cal_lut\[30\] a_20860_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1621 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6552_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1622 vssd1 a_6982_7093# a_6940_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1623 vssd1 a_14250_15797# a_14208_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1624 a_19199_13647# a_18501_13653# a_18942_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1625 a_27951_14013# a_27731_14025# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1626 a_16127_20288# cal_lut\[41\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1627 vssd1 a_25014_25183# a_24972_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1628 temp1.i_precharge_n a_1683_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1629 vccd1 a_12263_20495# _0481_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1631 a_3418_25321# _0806_ a_2564_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1632 vccd1 _0438_ a_15207_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0746 ps=0.775 w=0.42 l=0.15
X1634 a_5813_22895# _0434_ _0818_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1635 _0810_ a_4843_15307# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1636 vccd1 net36 a_24407_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1637 a_16585_13353# _0596_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X1638 vssd1 cal_lut\[75\] a_25552_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1641 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1642 a_10046_9001# _0493_ a_10046_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X1643 vccd1 a_20119_28701# a_20287_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1644 vssd1 _0418_ a_4431_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0894 ps=0.925 w=0.65 l=0.15
X1645 a_7255_20871# _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1646 a_13997_3855# _0131_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1648 _0447_ a_14103_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1649 a_12736_4233# a_12337_3861# a_12610_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1650 vccd1 a_26946_21919# a_26873_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1651 vssd1 a_9615_8181# a_9573_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1652 a_10505_22895# _0716_ _0718_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1653 vssd1 a_10857_21781# _0675_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X1654 vssd1 _0873_ a_19991_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1655 a_8175_11445# a_8351_11777# a_8303_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1656 vccd1 a_17283_28853# _0217_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1657 a_4333_27797# a_4167_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1658 a_13672_5737# _0502_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1659 vccd1 _0459_ a_19977_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1660 vssd1 _0330_ a_17919_3073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1661 vssd1 _0444_ a_21441_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1662 vssd1 a_7407_12533# a_7365_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1664 vccd1 clknet_0__0380_ a_6537_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1666 io_out[5] a_2564_25045# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1667 a_23205_17705# _0475_ a_23407_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1668 a_13269_9001# _0569_ a_13173_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1669 a_14618_24501# a_14450_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1670 vssd1 _0755_ a_8478_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X1671 a_4406_8863# a_4238_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1672 a_4798_21263# _0747_ a_4495_21495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X1673 a_6522_8863# a_6354_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1674 vccd1 a_8419_11195# a_8335_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1676 a_2835_30006# _0801_ a_2376_30199# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1677 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1678 a_18629_9295# a_18291_9527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1679 _0682_ _0675_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X1681 a_21217_18543# dbg_result[3] a_21133_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.0878 ps=0.92 w=0.65 l=0.15
X1682 a_15097_17455# a_14931_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1683 a_21073_3311# a_20083_3311# a_20947_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1684 a_17033_9295# _0106_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1685 vccd1 a_24099_12777# a_24106_12681# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1686 a_7994_13215# a_7826_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1687 vccd1 a_6375_19095# _0432_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1688 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1690 _0817_ a_9096_27221# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1691 cal_lut\[4\] a_10627_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1693 a_10975_20969# _0678_ a_10975_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X1694 vssd1 _0465_ a_19225_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1695 a_7975_18909# a_7277_18543# a_7718_18679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X1696 vccd1 a_13203_3829# a_13119_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1697 vccd1 a_25410_10901# a_25339_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1698 a_9223_24527# _0725_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1699 vssd1 net34 a_26983_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1700 a_1846_12559# a_1407_12565# a_1761_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1701 a_25524_23817# a_25125_23445# a_25398_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1702 vccd1 a_19667_18517# a_19303_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X1703 a_17555_19319# _0464_ a_17789_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1704 vccd1 a_3852_14165# _0394_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1705 _0150_ a_19439_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1706 a_17673_6941# a_17139_6575# a_17578_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1708 temp1.dac_vout_notouch_ net66 a_3424_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1709 vssd1 _0420_ a_3990_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1710 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2503_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1711 _0734_ dec1.i_ones a_8229_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1712 a_22051_6941# a_21187_6575# a_21794_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1713 a_24941_7119# a_24407_7125# a_24846_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1714 vssd1 a_23450_7775# a_23408_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1715 vccd1 a_22523_5175# _0687_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1716 _0458_ a_21003_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1717 vssd1 cal_lut\[21\] a_11797_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1718 a_9053_22895# _0712_ a_8971_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1720 vccd1 a_21883_1109# _0335_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1722 vccd1 a_7239_12381# a_7407_12283# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1724 vssd1 a_16055_19899# a_16013_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1725 a_18698_19319# a_19057_19319# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1726 a_24827_24501# a_25003_24833# a_24955_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1727 a_17397_20291# _0582_ a_17325_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1728 vssd1 net37 a_21923_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1729 a_15312_2057# a_14913_1685# a_15186_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1732 vccd1 a_9429_19605# a_9459_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1733 a_19303_16519# net18 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1734 a_8539_2986# _0367_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1735 a_6055_10602# _0375_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1736 vssd1 clknet_0__0380_ a_8390_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1737 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1738 vssd1 a_1919_20693# _0762_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1740 a_12153_2223# a_11987_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1742 a_7553_10927# a_7387_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1743 a_23207_12559# a_23027_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1744 a_25387_5161# net33 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1746 vssd1 a_17291_29397# a_17298_29697# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1747 vccd1 a_3325_8903# _0323_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X1748 a_9864_30511# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1749 vccd1 _0728_ a_7939_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1750 a_25502_21781# a_25302_22081# a_25651_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1751 a_5675_13469# a_4977_13103# a_5418_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1752 vssd1 net35 a_16679_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1753 vccd1 cal_lut\[189\] a_5083_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1754 a_10423_26703# _0385_ _0196_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1755 cal_lut\[24\] a_20287_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1757 a_18709_5487# cal_lut\[161\] a_18637_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1758 a_18673_7663# a_18119_7637# a_18326_7637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1759 vccd1 a_18475_19783# _0579_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1760 a_20303_28879# a_19605_28885# a_20046_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1761 vssd1 a_10784_23983# _0708_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1762 a_8419_25071# _0714_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1763 a_2288_17973# net7 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1764 a_8303_11837# cal_lut\[37\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X1765 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1766 a_10975_20719# _0676_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1768 a_20942_20969# _0872_ a_20860_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1769 a_12597_7809# _0572_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1771 vccd1 a_9551_2388# _0181_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1772 vccd1 _0014_ a_24653_12937# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1773 _0465_ a_21721_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.104 ps=1 w=0.65 l=0.15
X1774 a_12015_15645# a_11233_15279# a_11931_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1776 _0342_ a_20815_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
R4 temp1.capload\[3\].cap_58.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1777 vssd1 net78 _0407_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1778 a_23585_21807# cal_lut\[63\] a_23513_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1779 _0411_ a_1651_14165# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1780 a_6909_2223# a_6743_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1781 vccd1 cal_lut\[109\] a_23886_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1782 a_19027_9661# a_18807_9673# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1783 a_14729_10389# a_14563_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1785 _0025_ a_23763_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1786 _0156_ a_19807_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1788 vccd1 cal_lut\[120\] a_7786_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1789 a_3517_19087# _0419_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1790 a_3606_10660# a_3399_10601# a_3782_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1791 vccd1 net32 a_17139_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1792 vccd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ temp1.capload\[8\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1793 a_25634_18793# _0246_ a_25552_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1794 a_15680_4233# a_15281_3861# a_15554_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1795 _0147_ a_11711_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1796 _0476_ a_23763_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1798 cal_lut\[101\] a_15595_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1799 a_4222_12533# a_4054_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1800 vccd1 a_8565_28879# a_8671_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X1801 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1802 a_12827_10927# a_12698_11201# a_12407_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1804 a_24271_17277# a_24051_17289# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1805 a_14913_1685# a_14747_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1806 a_25566_23413# a_25398_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1807 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1808 a_13139_7351# _0441_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1809 a_24761_22895# _0031_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1810 vccd1 a_24485_17607# _0251_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X1811 a_5181_16617# _0382_ a_4816_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1812 vssd1 a_20499_8439# _0583_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1813 vccd1 cal_lut\[103\] a_20114_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1814 a_3535_10761# a_3399_10601# a_3115_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1815 a_6277_24233# _0429_ _0797_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1817 vssd1 clknet_0_net67 a_3685_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1818 vccd1 net30 a_11527_9303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1819 a_15557_27497# cal_lut\[92\] a_15473_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1820 a_18291_16532# _0254_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1822 a_5801_4233# a_4811_3861# a_5675_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1823 a_11797_12925# a_11527_12559# a_11707_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X1824 a_10543_15823# a_9761_15829# a_10459_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1825 a_1477_10901# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1826 a_22441_21237# _0636_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1827 vssd1 a_5323_4917# _0319_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1828 a_3974_21807# _0753_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X1829 vccd1 _0543_ a_15477_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1830 a_22779_8207# a_21997_8213# a_22695_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1831 _0836_ a_3155_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1832 vccd1 a_27498_8863# a_27425_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1833 a_4054_12559# a_3781_12565# a_3969_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1834 vccd1 a_13035_14557# a_13203_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1835 a_5324_4373# net39 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1836 vssd1 cal_lut\[99\] a_12349_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1837 a_19421_10927# a_19255_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1838 a_14082_15823# a_13643_15829# a_13997_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1839 _0295_ a_20676_5059# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1840 vccd1 a_2773_9991# _0837_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X1841 vccd1 a_19367_13621# a_19283_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1842 vssd1 net25 a_12171_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1843 vccd1 _0472_ a_15483_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1844 a_5554_19631# _0737_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1845 vccd1 a_13291_18909# _0474_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1846 a_18958_16911# a_18519_16917# a_18873_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1847 a_18958_16911# a_18685_16917# a_18873_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1848 vssd1 _0477_ a_17385_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1849 a_18501_13653# a_18335_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1852 a_17075_27613# a_16293_27247# a_16991_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1853 a_12141_8751# a_11594_9025# a_11794_8725# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1854 a_20522_3677# a_20249_3311# a_20437_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1855 vccd1 _0358_ a_27351_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1856 vssd1 _0668_ a_11277_19659# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1857 _0159_ a_24315_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1858 a_4912_8439# net39 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X1859 vccd1 a_24105_10357# _0695_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X1860 a_20308_27497# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1861 a_5105_25045# _0747_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1862 vccd1 _0681_ a_11142_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1863 vssd1 a_18475_18695# _0605_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 a_21831_11471# _0449_ a_22009_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1865 _0515_ _0491_ a_14855_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1866 vccd1 a_5013_24825# a_5043_24566# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1867 a_10943_23671# _0675_ a_11117_23777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1869 _0483_ a_15207_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=1.62 w=1 l=0.15
X1870 a_9275_28023# _0815_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1871 vccd1 net29 a_11067_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1872 a_20245_28335# a_19255_28335# a_20119_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1873 a_27531_13469# a_27351_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1874 a_4898_10749# a_4583_10615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1876 _0729_ _0708_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1877 a_15649_3855# a_15115_3861# a_15554_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1878 a_21537_16367# a_21371_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1879 vccd1 a_24407_15279# _0246_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1880 vssd1 a_15163_9527# _0562_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1881 vssd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1882 _0800_ a_4678_26311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X1884 vccd1 a_7618_26935# _0409_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X1885 a_10603_23439# _0679_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1886 vssd1 cal_lut\[187\] a_7381_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1887 a_14151_11079# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1888 vccd1 net35 a_20819_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1889 vccd1 a_11639_14459# a_11555_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1890 vssd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1892 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1893 vssd1 a_13403_23261# a_13571_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1894 vssd1 dbg_result[1] a_20543_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1895 a_13139_7351# _0441_ a_13373_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1896 _0316_ a_10108_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1897 vssd1 a_21362_26133# a_21291_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1898 vccd1 io_in[1] a_1407_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1899 vccd1 _0440_ a_17599_6039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1900 _0679_ a_10975_20969# a_11508_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1901 _0754_ a_2417_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X1902 vssd1 a_7239_14735# a_7410_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1903 _0748_ _0721_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.114 ps=1 w=0.65 l=0.15
X1905 a_15903_3285# cal_lut\[179\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X1907 vssd1 a_3851_15253# _0198_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.0878 ps=0.92 w=0.65 l=0.15
X1908 vccd1 a_25042_5461# a_24971_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1909 a_14959_24527# a_14177_24533# a_14875_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1911 cal_lut\[133\] a_8695_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1912 a_24630_10089# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X1914 vccd1 a_7369_28879# a_7475_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X1915 a_17677_23983# _0082_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1916 _0868_ a_23759_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1917 vccd1 net45 a_20727_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1919 a_22339_27399# a_22435_27221# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1920 vssd1 cal_lut\[62\] a_23489_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1921 vssd1 a_16991_27613# a_17159_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1922 _0228_ a_20308_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1923 _0824_ a_2563_23957# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1924 a_21166_11293# a_20893_10927# a_21081_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1925 dbg_result[1] a_6674_16620# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
R5 vssd1 net55 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1926 vccd1 a_25962_11989# a_25891_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1927 a_7111_28585# ctr\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X1928 vccd1 a_27847_7119# a_28015_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1929 a_4479_12559# a_3781_12565# a_4222_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1930 vssd1 _0866_ a_18611_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1931 _0145_ a_7571_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1933 a_2947_10615# a_3115_10615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1934 a_2234_28157# _0824_ a_1735_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X1936 a_20119_11293# a_19255_10927# a_19862_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1937 a_4054_12559# a_3615_12565# a_3969_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1938 _0680_ _0520_ a_8979_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
X1939 vccd1 _0454_ a_18611_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1940 a_6182_22895# clknet_0_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1941 a_28157_17455# a_27167_17455# a_28031_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1942 a_13490_5737# _0568_ a_13241_5633# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X1943 a_7553_10927# a_7387_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1944 vccd1 net37 a_27167_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1945 a_4679_19319# _0425_ a_4805_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1947 vccd1 a_4831_9019# a_4747_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1948 vccd1 a_7895_12778# _0019_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1949 _0253_ a_17135_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X1950 a_14821_27797# a_14655_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1952 a_20499_8439# _0441_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1953 a_11302_16519# _0625_ a_11516_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X1954 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1955 _0870_ a_24863_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1957 vssd1 _0817_ temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1958 vccd1 a_22466_19605# a_22395_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1959 a_17732_14441# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1960 vccd1 a_20471_28853# a_20387_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1961 vccd1 _0420_ a_2900_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 vssd1 a_17895_17973# a_17853_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1963 vssd1 _0452_ a_16889_22689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1964 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1965 vssd1 net47 a_24407_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1967 a_23776_19465# a_23377_19093# a_23650_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1968 vssd1 _0235_ a_21279_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1969 vccd1 net2 a_6927_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1970 a_14273_15431# _0872_ a_14436_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1971 a_10360_10383# _0492_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1972 net14 a_10239_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1973 cal_lut\[92\] a_15687_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1974 a_1917_19881# _0428_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.585 pd=2.17 as=0.135 ps=1.27 w=1 l=0.15
X1975 a_17543_9295# a_16679_9301# a_17286_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1976 _0552_ a_16955_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1977 a_20119_5853# a_19421_5487# a_19862_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1979 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1980 _0123_ a_11527_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1981 vccd1 a_14331_3285# a_14155_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1982 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1983 vccd1 a_20690_21237# a_20617_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1984 a_12525_14191# _0096_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1985 a_27425_9117# a_26891_8751# a_27330_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1987 a_6703_6549# cal_lut\[144\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X1988 a_7097_6031# _0144_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1989 _0808_ a_2695_14013# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.175 ps=1.26 w=0.65 l=0.15
X1990 a_11756_22671# _0709_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.127 ps=1.04 w=0.65 l=0.15
X1991 a_27329_21807# a_26339_21807# a_27203_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1992 a_2489_17455# _0422_ a_2931_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1994 _0060_ a_21279_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1995 vccd1 a_6674_16620# a_6587_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X1996 a_10977_10499# _0694_ a_10881_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1997 vccd1 a_19333_25223# _0221_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X1998 a_7021_22671# _0786_ a_6611_22583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1999 a_9429_19605# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2002 vssd1 a_15687_29691# a_15645_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2003 vccd1 a_26743_16733# a_26911_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2004 a_9201_3829# _0476_ a_9454_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X2006 vssd1 _0449_ a_17680_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X2007 net48 a_6927_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2008 a_26226_6941# a_25953_6575# a_26141_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2009 vssd1 a_2327_22895# _0418_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2011 vssd1 cal_lut\[9\] a_13453_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2012 a_9167_21601# _0677_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2013 vccd1 _0720_ _0732_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2014 vccd1 cal_lut\[115\] a_22322_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2015 vccd1 net29 a_9687_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2017 a_27606_10205# a_27333_9839# a_27521_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2018 vccd1 cal_lut\[4\] a_10914_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2019 a_22059_1109# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2021 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2022 a_14523_16885# dbg_result[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2023 a_23719_12791# a_23815_12791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2024 vccd1 _0704_ _0705_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2025 a_1673_22351# ctr\[1\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2026 _0502_ a_18645_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X2027 cal_lut\[171\] a_28199_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2028 a_17411_29245# cal_lut\[43\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X2029 vssd1 a_20598_16885# a_20556_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2030 a_3695_23671# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.165 ps=1.33 w=1 l=0.15
X2031 a_9548_4399# _0495_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X2032 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2033 a_16481_21807# _0041_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2034 vssd1 net23 a_8951_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2035 a_7826_6941# a_7387_6575# a_7741_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2036 _0459_ a_19439_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2038 _0853_ a_17732_14441# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2039 vccd1 a_11366_28588# dbg_result[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X2040 a_1963_21365# _0414_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X2041 vccd1 a_17739_7815# cal_lut\[112\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2043 _0436_ a_1683_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2044 a_2313_15823# _0198_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2045 a_19421_10927# a_19255_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2046 vccd1 a_19681_12161# _0525_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2047 _0841_ a_13459_22359# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2048 vssd1 a_7072_15797# net41 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2049 a_20499_8439# _0441_ a_20733_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2050 a_4811_17705# clknet_1_0__leaf__0380_ _0384_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2052 vssd1 net47 a_21831_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2053 net38 a_16731_9813# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2054 a_19333_24135# cal_lut\[83\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X2055 _0063_ a_25787_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2056 temp1.capload\[1\].cap.Y net56 a_1677_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2057 _0389_ _0411_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2058 vssd1 a_9595_3311# net25 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2059 _0654_ a_11527_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X2060 vccd1 _0379_ a_2879_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2061 vccd1 _0390_ a_4981_28940# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X2062 vssd1 a_5227_26935# _0812_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2063 a_15541_9985# _0549_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2064 a_25295_21781# net43 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2065 _0676_ _0667_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2066 a_15494_19319# dbg_result[1] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X2067 a_15531_4564# _0365_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2068 a_10827_3677# a_9963_3311# a_10570_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2069 vccd1 net27 a_5915_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2070 a_9452_32375# net11 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2071 vssd1 _0681_ a_10784_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2073 a_18807_9673# a_18671_9513# a_18387_9527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2074 a_3848_27399# _0826_ a_3990_27574# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X2076 _0192_ ctr\[2\] a_5377_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2077 _0626_ _0609_ a_11895_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2078 vssd1 a_15963_28853# a_15921_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2079 a_19303_18695# dbg_result[1] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X2080 a_27123_15431# a_27219_15253# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2081 a_25345_4943# a_25007_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2082 vssd1 a_3399_10601# a_3406_10505# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2085 a_25218_19997# a_24971_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2086 a_6982_7093# a_6814_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2087 a_19308_17973# _0507_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2088 a_22875_9867# _0450_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2089 a_14733_15431# cal_lut\[35\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X2090 vssd1 a_23719_4087# cal_lut\[117\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2091 a_8251_29789# a_7387_29423# a_7994_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2092 vccd1 _0841_ a_12815_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X2093 vccd1 cal_lut\[120\] a_15991_8903# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2095 a_4484_30663# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2096 a_25839_14165# a_26130_14465# a_26081_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2097 vssd1 _0857_ a_23763_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2098 a_5451_3677# a_5271_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2099 vssd1 _0465_ a_18085_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2101 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2102 vccd1 clknet_1_0__leaf__0380_ a_5460_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2103 a_10178_10383# _0515_ a_9929_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X2104 a_15603_27791# a_14821_27797# a_15519_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2105 a_5503_27399# a_5599_27221# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2106 a_9372_24135# _0723_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X2107 cal_lut\[10\] a_14123_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2109 vssd1 a_9929_10357# _0516_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X2110 vssd1 _0444_ a_22269_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2112 io_out[0] a_2023_19319# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2113 ctr\[3\] a_3175_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 vccd1 a_11639_5755# a_11555_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2115 vccd1 _0805_ _0806_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2116 a_9542_4649# _0495_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X2118 a_12219_17130# _0845_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2119 a_13453_23983# a_13183_24349# a_13363_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2120 vccd1 _0467_ a_15023_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2121 vssd1 _0450_ a_22843_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2122 a_7749_28335# a_7557_28640# _0210_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2123 a_27931_7119# a_27149_7125# a_27847_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2124 a_11587_8725# net29 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2125 a_24235_12937# a_24106_12681# a_23815_12791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2126 cal_lut\[10\] a_14123_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2127 vccd1 _0330_ a_22291_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X2128 vssd1 ctr\[12\] a_8329_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2130 a_18669_22325# _0620_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2132 a_25106_15797# a_24938_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2133 vssd1 net24 a_6375_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2134 vccd1 a_8146_18796# dbg_result[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2135 vssd1 cal_lut\[124\] a_13592_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2136 a_15071_13268# _0852_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2137 a_9471_29097# clknet_1_1__leaf_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2138 vccd1 a_7716_22325# _0786_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2139 a_14331_3285# _0290_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2140 a_5157_28169# a_4167_27797# a_5031_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2141 a_5864_26819# _0811_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2142 a_15557_25071# a_15391_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2144 a_4068_32463# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2145 vccd1 a_12263_20495# _0481_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2146 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2147 vccd1 a_15207_18543# _0483_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2148 vccd1 _0294_ a_18887_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2149 a_13353_12559# _0191_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2150 a_26417_18231# cal_lut\[70\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X2151 vssd1 _0493_ a_13172_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X2152 a_13840_29257# a_13441_28885# a_13714_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2153 a_11020_21807# _0671_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X2156 a_16635_26324# _0215_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2157 a_23197_7663# _0109_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2158 cal_lut\[89\] a_18539_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2159 a_22235_22173# a_21537_21807# a_21978_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2160 a_27211_8513# _0341_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2161 a_3781_12565# a_3615_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2162 vssd1 a_18187_1679# a_18355_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2164 vssd1 cal_lut\[110\] a_19709_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2165 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_8951_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2166 vssd1 a_17381_15425# _0554_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X2169 vssd1 a_2419_12015# _0390_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2171 a_10773_14191# a_10607_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2172 vssd1 _0316_ a_5499_5249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2173 vccd1 a_6603_11777# a_6427_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2174 a_15097_28885# a_14931_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2175 a_6503_16733# a_5805_16367# a_6246_16503# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X2176 a_5391_29789# a_4609_29423# a_5307_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2178 vssd1 _0421_ _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2179 a_25375_12167# a_25471_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2180 vccd1 a_7895_11690# _0037_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2181 a_2504_17271# a_2317_16911# a_2417_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X2182 vccd1 dbg_result[3] a_13291_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2183 cal_lut\[6\] a_12927_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2184 vssd1 a_9005_24501# _0728_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2185 a_22435_27221# a_22719_27221# a_22654_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2186 a_8055_25321# dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2187 vssd1 a_19057_26935# _0227_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2189 a_15519_29789# a_14655_29423# a_15262_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2190 a_13291_18909# a_13508_18517# a_13466_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2191 vssd1 _0712_ a_10517_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2192 vssd1 a_17727_2589# a_17895_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2193 a_23009_7663# a_22843_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2194 a_15001_24905# a_14011_24533# a_14875_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2195 vccd1 a_13459_22359# _0841_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2196 vccd1 net44 a_19807_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2197 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2198 vccd1 _0025_ a_24469_17289# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2199 a_4461_25913# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2200 a_23355_23671# cal_lut\[56\] a_23481_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2201 a_27774_17567# a_27606_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2202 vccd1 cal_lut\[164\] a_24630_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2203 a_6377_26409# _0399_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2205 a_11605_16055# _0836_ a_11768_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2206 a_9033_13353# _0501_ a_9117_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2207 net8 a_10844_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2208 a_1743_18259# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2209 cal_lut\[183\] a_10995_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2210 a_8611_3855# a_7829_3861# a_8527_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2211 _0159_ a_24315_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2212 vssd1 a_15503_7093# a_15461_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2213 a_4406_9951# a_4238_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2214 a_15189_29789# a_14655_29423# a_15094_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2215 vssd1 a_7994_11039# a_7952_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2216 vssd1 net33 a_22843_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2217 a_7565_23983# _0752_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2218 vssd1 a_15370_19407# _0467_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2219 a_23815_4087# a_24099_4073# a_24034_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2220 vssd1 cal_lut\[128\] a_10280_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2221 a_4947_5249# _0316_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2223 a_4491_13879# _0808_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2224 _0661_ _0650_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0894 ps=0.925 w=0.65 l=0.15
X2225 _0873_ a_19756_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2226 vssd1 cal_lut\[161\] a_25873_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2229 a_12383_3677# a_11601_3311# a_12299_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2230 vccd1 net32 a_21187_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2231 a_7553_8751# a_7387_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2232 vssd1 a_27802_13924# a_27731_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2233 a_7952_6575# a_7553_6575# a_7826_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2234 a_10347_25321# _0720_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2235 a_14039_23439# a_13257_23445# a_13955_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2236 vssd1 ctr\[10\] a_7133_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2237 a_7289_25321# _0733_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2238 _0429_ a_3615_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2239 vccd1 cal_lut\[30\] a_20407_16519# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2240 vccd1 _0451_ a_12079_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X2241 cal_lut\[154\] a_21759_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2242 vccd1 a_20690_3423# a_20617_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2244 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2245 a_27731_14025# a_27602_13769# a_27311_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2246 vccd1 a_15979_12559# a_16147_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2247 cal_lut\[69\] a_25531_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2248 a_27774_15797# a_27606_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2249 _0564_ a_14287_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2250 a_19681_12161# _0524_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2251 vccd1 a_23811_27412# _0055_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2252 a_18274_15529# _0851_ a_18192_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2253 a_6607_9514# _0322_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2254 a_2939_23047# ctr\[1\] a_3113_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2255 a_4189_15279# _0411_ a_4091_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.111 ps=0.99 w=0.65 l=0.15
X2256 a_21591_25437# a_20727_25071# a_21334_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2258 a_4401_28918# _0801_ a_4187_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2259 a_4253_7663# a_3983_8029# a_4163_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2260 vssd1 a_15979_12559# a_16147_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2262 _0243_ a_23299_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2264 vccd1 net30 a_3707_9303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2266 _0283_ a_13459_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2267 vssd1 net38 a_16679_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2269 vccd1 net27 a_6375_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2271 a_8454_4917# a_8286_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2272 vssd1 net24 a_4259_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2273 a_6929_20719# a_6646_21041# a_6516_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2274 a_21717_2223# a_20727_2223# a_21591_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2275 _0862_ a_9131_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2276 vssd1 io_in[5] a_1407_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2278 a_5008_29423# a_4609_29423# a_4882_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2279 a_4811_25935# _0801_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X2280 vccd1 a_5843_13371# a_5759_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2281 a_12433_1679# _0183_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2282 a_7843_5487# cal_lut\[145\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X2283 a_22619_15253# net38 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2284 a_25295_21781# net43 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2285 vccd1 _0464_ a_15959_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2286 vccd1 clknet_1_0__leaf_io_in[0] a_7111_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2287 a_20756_12559# _0535_ a_20654_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2288 a_21261_25437# a_20727_25071# a_21166_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2289 a_25042_13077# a_24842_13377# a_25191_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2290 vssd1 a_14307_4917# a_14265_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2291 a_16771_23439# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2292 vccd1 a_6245_21781# _0820_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2293 a_17197_19777# _0579_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2295 vssd1 a_10995_1653# a_10953_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2296 a_17993_10955# _0445_ a_17907_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2297 a_22649_24233# _0468_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2298 vssd1 a_13111_1653# a_13069_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2299 a_21136_27497# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2300 a_4472_21807# _0757_ a_4381_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X2301 a_3299_19061# _0744_ a_3730_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X2303 vccd1 net81 a_16069_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2305 vccd1 a_2419_12015# _0390_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2306 vssd1 a_4495_21495# _0781_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2307 a_6800_5059# cal_lut\[135\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X2308 vssd1 net28 a_8951_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2309 a_27167_14557# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2310 a_23759_13469# a_23579_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2311 a_21997_27797# a_21831_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2312 a_2504_27023# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2313 a_13897_21641# a_12907_21269# a_13771_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2315 ctr\[0\] a_2439_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2316 vssd1 a_12299_3677# a_12467_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2317 a_15667_20719# cal_lut\[40\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2318 a_25253_22173# a_24915_21959# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2319 vccd1 _0411_ a_1773_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X2320 a_4066_7396# a_3866_7241# a_4215_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2321 vssd1 a_1945_15431# _0388_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2322 a_8987_14735# a_8123_14741# a_8730_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2323 a_28157_9839# a_27167_9839# a_28031_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2324 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2325 vccd1 cal_lut\[124\] a_13674_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2327 vssd1 a_14273_15431# _0880_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2328 a_7716_25589# _0734_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X2329 vccd1 a_25962_20452# a_25891_20553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2330 vssd1 _0033_ a_26309_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2331 vssd1 _0350_ a_25143_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2332 _0712_ a_11896_24233# a_12097_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2333 _0560_ a_18611_20288# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2334 a_17129_23145# _0500_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2335 a_26580_18115# cal_lut\[70\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X2337 vssd1 a_25271_7119# a_25439_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2338 a_10252_11849# a_9853_11477# a_10126_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2339 a_27931_17999# a_27149_18005# a_27847_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2340 vssd1 net32 a_17139_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2341 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2342 a_21428_7913# cal_lut\[111\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X2343 vccd1 a_16807_11293# a_16975_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2344 a_21169_11471# cal_lut\[158\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2346 vssd1 a_14243_16532# _0035_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2347 _0864_ a_11707_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2348 _0539_ _0534_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0894 ps=0.925 w=0.65 l=0.15
X2349 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6007_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2351 vccd1 a_16373_16341# _0625_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X2353 a_5775_19631# ctr\[2\] a_5412_19783# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2354 vssd1 a_9558_14303# a_9516_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2355 vccd1 cal_lut\[5\] a_12938_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2356 vssd1 _0721_ _0734_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X2357 a_8657_14735# a_8123_14741# a_8562_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2358 a_12079_5737# _0502_ a_12162_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X2359 vssd1 a_21978_16479# a_21936_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2360 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2361 a_27595_13865# net37 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2362 a_10827_3677# a_10129_3311# a_10570_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2363 vccd1 a_6637_5175# _0318_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X2364 vssd1 a_22863_8181# a_22821_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2365 vccd1 _0175_ a_26309_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2366 a_5724_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2367 cal_lut\[27\] a_24243_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2368 vccd1 a_24519_14709# a_24435_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2370 a_10692_30287# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2371 a_26325_18543# _0075_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2372 vssd1 net19 a_21029_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2373 vssd1 a_13219_27613# a_13387_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2374 vccd1 a_7239_7119# a_7407_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2375 temp1.capload\[3\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2376 vccd1 a_26099_17821# a_26267_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2377 a_23653_14741# a_23487_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2380 vssd1 cal_lut\[50\] a_14465_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2381 a_20256_12015# cal_lut\[162\] a_19681_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X2382 a_20525_16911# a_19991_16917# a_20430_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2383 _0229_ a_21136_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2384 vssd1 ctr\[3\] a_3852_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X2385 vccd1 net23 a_7663_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2386 vccd1 a_7975_14557# a_8143_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2387 vccd1 a_17711_9269# a_17627_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2388 a_24636_9839# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X2390 vssd1 _0412_ a_3339_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2391 a_10416_31599# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2392 vccd1 _0225_ a_14747_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2394 _0581_ a_15667_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2395 vssd1 a_5412_19783# _0738_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2396 a_2485_22351# clknet_1_1__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2397 cal_lut\[81\] a_11639_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2398 _0617_ a_16390_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X2399 vssd1 a_2099_18695# _0743_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.179 ps=1.85 w=0.65 l=0.15
X2400 a_18383_5175# _0514_ a_18617_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2401 a_10041_13103# _0020_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2402 a_23351_21959# _0531_ a_23585_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2403 a_12318_26677# a_12150_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2404 a_25769_9839# a_25603_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2405 net40 a_12723_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2406 a_18087_6941# a_17305_6575# a_18003_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2407 vssd1 a_18647_28879# a_18815_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R6 temp1.capload\[0\].cap_49.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2408 a_7553_29423# a_7387_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2409 a_12597_7809# _0570_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2410 vssd1 a_2377_28500# temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2411 a_25355_7119# a_24573_7125# a_25271_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2412 vssd1 _0660_ _0661_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X2415 a_20216_22057# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2416 a_19609_15279# _0023_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2417 vccd1 a_2939_23047# _0417_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X2418 a_5825_15823# _0381_ a_5460_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2420 vccd1 a_26394_6687# a_26321_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2421 a_10589_27247# a_10423_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2422 a_23039_3145# a_22903_2985# a_22619_2999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2423 _0279_ a_14375_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2424 a_19303_23047# _0454_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2425 a_12150_26703# a_11877_26709# a_12065_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2426 vssd1 _0439_ a_8491_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2427 a_24469_17289# a_23915_17129# a_24122_17188# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2428 a_7350_10357# a_7182_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2429 vssd1 a_7071_25045# _0735_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2430 vssd1 cal_lut\[20\] a_9221_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2431 vccd1 _0497_ a_10029_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2434 a_19694_11293# a_19421_10927# a_19609_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2435 a_25471_11989# a_25755_11989# a_25690_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2436 a_20713_19631# _0059_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2437 a_24051_17289# a_23922_17033# a_23631_17143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2439 vccd1 a_17415_7119# net34 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2440 vccd1 a_11896_24233# _0712_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2441 vssd1 net29 a_11067_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2442 a_13441_4949# a_13275_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2443 vccd1 cal_lut\[76\] a_17555_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2444 a_7168_4649# cal_lut\[133\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X2445 vssd1 _0862_ a_9595_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2446 a_12893_25071# _0008_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2447 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2448 vccd1 _0237_ a_23119_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X2449 vccd1 a_15703_2767# a_15871_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2451 a_9941_1135# a_8951_1135# a_9815_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2452 a_12245_1685# a_12079_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2453 a_16390_5487# _0615_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X2454 vssd1 _0664_ a_10677_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2458 vccd1 a_19583_2741# _0338_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X2459 vssd1 net32 a_19715_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2460 vccd1 _0784_ a_4401_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2462 a_4217_30006# _0801_ a_4003_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2463 a_23791_8029# a_23009_7663# a_23707_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2464 cal_lut\[75\] a_25623_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2465 a_2355_14735# a_1573_14741# a_2271_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2466 vssd1 _0492_ a_16116_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X2468 a_20441_20719# _0531_ a_20359_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2469 a_23823_20393# net43 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2470 a_4273_26159# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2471 _0752_ _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X2472 vccd1 _0454_ a_16127_20288# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2473 _0447_ a_14103_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2474 vccd1 _0500_ a_9117_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2475 vssd1 _0744_ a_3338_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X2476 a_12617_13103# _0021_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2477 a_21334_25183# a_21166_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2478 a_20010_12265# _0523_ a_19930_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2479 a_15262_23413# a_15094_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2480 vssd1 _0152_ a_23457_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2481 a_11279_28701# a_10497_28335# a_11195_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X2482 vssd1 _0097_ a_13245_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2484 vccd1 _0370_ a_11987_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2485 a_22779_27791# a_21997_27797# a_22695_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2486 vssd1 _0591_ a_9821_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2487 _0266_ a_12355_21271# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2489 vssd1 a_23763_4943# _0476_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2491 io_out[5] a_2564_25045# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2492 vssd1 cal_lut\[32\] a_24769_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2493 a_15623_15431# _0467_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2494 a_11881_7119# _0123_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2495 a_4211_27247# _0826_ a_3848_27399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2496 a_20154_9295# a_19881_9301# a_20069_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2497 a_27521_17455# _0073_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2498 _0028_ a_18611_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2499 a_16340_7913# _0515_ a_16238_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2500 vccd1 _0744_ a_3351_27569# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X2501 vccd1 a_21334_25183# a_21261_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2502 vccd1 a_10995_3579# a_10911_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2503 vccd1 a_24094_14709# a_24021_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2504 vssd1 cal_lut\[182\] a_9876_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X2505 vssd1 a_15531_24135# _0645_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2506 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2507 a_14465_28335# a_14195_28701# a_14375_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2508 vccd1 a_2722_20175# _0424_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2509 a_22235_16733# a_21371_16367# a_21978_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2510 vccd1 clknet_1_1__leaf_io_in[0] a_4167_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2511 cal_lut\[4\] a_10627_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2512 a_4528_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2513 _0475_ a_18369_18337# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X2514 _0861_ a_7751_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2515 vccd1 a_13019_2491# a_12935_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2517 _0883_ a_11891_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2518 a_15094_23439# a_14821_23445# a_15009_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2519 _0555_ _0554_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
X2520 a_19609_24527# _0083_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2521 _0241_ a_20216_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2523 a_25523_5321# a_25387_5161# a_25103_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2524 vccd1 ctr\[1\] a_3981_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2525 a_8454_4917# a_8286_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2526 a_18774_13647# a_18501_13653# a_18689_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2527 vssd1 a_22291_20175# net43 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2529 a_20482_15939# _0851_ a_20400_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2530 vssd1 _0294_ a_18887_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2531 a_7691_10383# a_6909_10389# a_7607_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2532 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_4811_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2533 a_19659_25615# a_18961_25621# a_19402_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2534 vccd1 a_5031_27791# a_5199_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2535 a_8093_22895# _0724_ a_8021_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2536 a_16373_16341# _0624_ a_16753_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X2539 a_1962_27791# a_1913_28023# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X2540 a_19234_25615# a_18795_25621# a_19149_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2541 vccd1 cal_lut\[88\] a_17135_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2543 vccd1 _0411_ a_4624_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2544 vccd1 a_10459_15823# a_10627_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2545 vccd1 _0335_ a_21463_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2546 vccd1 a_15715_5175# _0566_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2547 a_25743_14343# a_25839_14165# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2550 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2551 a_10746_10615# _0701_ a_11049_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X2552 a_14081_23817# a_13091_23445# a_13955_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2553 _0365_ a_15479_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2554 a_14523_6549# a_14699_6549# a_14651_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X2557 a_20390_14441# _0851_ a_20308_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2558 a_23811_4564# _0296_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2559 a_4413_7497# a_3859_7337# a_4066_7396# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2560 a_9411_8751# cal_lut\[139\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2561 a_8546_1653# a_8378_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2562 a_16904_25321# _0872_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2563 a_16845_14741# a_16679_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2564 vccd1 net26 a_10607_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2565 a_20525_19631# a_20359_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2567 a_8229_25071# dec1.i_ones _0734_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X2569 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2570 a_2933_14709# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X2571 _0571_ a_12539_6144# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2572 a_12705_25071# a_12539_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2573 a_13717_26709# a_13551_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2574 a_3525_20291# _0422_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2576 vccd1 a_13135_15253# a_12959_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2577 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2578 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2580 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2582 vssd1 a_18763_20871# _0486_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2583 a_13835_17277# _0447_ a_13751_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0567 ps=0.69 w=0.42 l=0.15
X2584 vccd1 a_20598_16885# a_20525_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2585 a_10787_4221# cal_lut\[132\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X2586 a_15588_19631# a_15189_19631# a_15462_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2587 a_7478_19453# ctr\[4\] a_6979_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X2588 a_7350_2335# a_7182_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2589 vssd1 net27 a_7387_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2590 vssd1 a_9673_23047# _0726_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2591 a_12429_13103# a_12263_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2592 vssd1 a_21265_7815# _0292_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2593 a_14449_27247# cal_lut\[50\] a_14103_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2594 cal_lut\[93\] a_14583_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2595 _0472_ _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2596 vssd1 a_23155_6031# a_23323_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2597 vccd1 _0442_ a_19715_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X2598 a_6449_3311# a_6283_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2599 a_24769_22717# a_24499_22351# a_24679_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2600 a_9773_25935# _0715_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2601 _0196_ _0385_ a_10423_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2602 vssd1 a_20119_15645# a_20287_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2603 a_7636_31849# a_7387_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2604 a_4003_30333# a_3749_30006# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X2605 _0411_ a_1651_14165# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2606 vssd1 a_20867_2986# _0153_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2608 a_26321_6941# a_25787_6575# a_26226_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2609 a_25539_17999# a_24757_18005# a_25455_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2611 vccd1 ctr\[8\] a_5661_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2612 vssd1 _0714_ a_8419_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2614 vssd1 _0676_ a_10975_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2615 vccd1 _0442_ a_15207_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.0588 ps=0.7 w=0.42 l=0.15
X2616 vssd1 a_4167_16367# _0839_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2617 vccd1 a_18187_25437# a_18355_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2618 a_13487_23261# a_12705_22895# a_13403_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2619 a_20119_5853# a_19255_5487# a_19862_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2621 vssd1 a_26651_6941# a_26819_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2622 vccd1 _0438_ a_13714_19407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X2623 vssd1 a_12223_2741# _0330_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2624 cal_lut\[111\] a_20747_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2625 _0637_ a_21923_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2626 a_8803_1679# a_8105_1685# a_8546_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2627 vssd1 _0299_ a_9765_6727# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2628 a_6081_29423# a_5915_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2629 _0265_ a_21872_25731# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2630 a_15094_23439# a_14655_23445# a_15009_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2631 a_15278_2767# a_15005_2773# a_15193_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2634 _0386_ a_9559_26481# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.178 ps=1.41 w=1 l=0.15
X2635 vssd1 clknet_0_net67 a_3685_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2636 a_18937_20747# _0485_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2637 a_26026_8181# a_25858_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2638 vssd1 a_15998_25183# a_15956_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2639 vccd1 _0838_ a_12355_21271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2640 vssd1 a_16635_26324# _0042_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2641 a_15484_18543# dbg_result[1] a_15378_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2642 vccd1 a_16757_7637# _0498_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2644 a_20201_18543# _0485_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2645 vssd1 cal_lut\[67\] a_23389_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2646 a_23239_6031# a_22457_6037# a_23155_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2647 vssd1 a_14156_11989# _0440_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2648 a_23849_13103# a_23579_13469# a_23759_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2649 vssd1 cal_lut\[19\] a_7841_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2650 a_21081_2223# _0153_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2651 cal_lut\[20\] a_8419_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2652 a_8309_19881# _0764_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2653 vccd1 a_18878_9572# a_18807_9673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2654 vccd1 net24 a_6743_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2655 _0101_ a_16035_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2656 a_10459_15823# a_9595_15829# a_10202_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2657 a_25014_24095# a_24846_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2659 vssd1 _0606_ a_17841_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2660 a_12623_30287# net13 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2662 vssd1 a_5199_27765# a_5157_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2663 a_15477_15823# _0546_ a_15371_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2664 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2666 _0003_ a_9595_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2667 a_13035_14557# a_12337_14191# a_12778_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2669 a_18243_19200# cal_lut\[70\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2670 vccd1 _0290_ a_10055_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X2671 _0769_ a_4892_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X2672 vssd1 _0327_ a_6375_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2673 vccd1 a_1963_21365# _0772_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2674 a_19609_4399# _0117_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2675 a_19961_14191# cal_lut\[12\] a_19889_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2676 a_5181_20719# _0768_ a_4771_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X2677 _0474_ a_13291_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.331 ps=1.71 w=1 l=0.15
X2678 _0069_ a_25327_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2679 vssd1 net35 a_18335_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2680 a_18255_7663# a_18126_7937# a_17835_7637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2681 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2682 _0299_ a_7439_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2683 vssd1 cal_lut\[114\] a_20676_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2685 a_17831_24746# _0220_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2686 a_18731_28879# a_17949_28885# a_18647_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2687 a_11277_19659# _0666_ a_11191_19659# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2688 a_11142_24233# _0707_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2689 a_18201_19659# _0467_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2690 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2691 a_11117_23777# _0679_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2692 vssd1 _0850_ a_24683_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2693 vccd1 a_14979_24148# _0094_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2695 a_2907_15823# a_2125_15829# a_2823_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2696 _0801_ _0800_ a_3171_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2698 vccd1 _0441_ a_12079_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2699 a_7839_32143# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X2700 a_14499_26703# a_13717_26709# a_14415_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2701 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2702 vccd1 net1 a_10699_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2703 vssd1 a_17739_7815# cal_lut\[112\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2704 a_17025_24847# cal_lut\[46\] a_16679_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2705 a_9677_16617# cal_lut\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2707 vccd1 a_9201_3829# _0700_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X2708 a_13714_19407# _0447_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X2709 net11 a_8543_30485# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2710 vccd1 _0507_ a_18243_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2711 vccd1 _0188_ a_5517_10761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2712 a_24648_17705# cal_lut\[74\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X2713 vssd1 a_14986_5599# a_14944_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2714 vssd1 _0105_ a_19225_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2715 a_24853_15823# _0068_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2716 a_17029_2223# a_16863_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2717 a_9558_1247# a_9390_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2719 a_18961_25621# a_18795_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2720 vccd1 cal_lut\[137\] a_17095_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2721 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9496_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2724 a_18497_26159# a_17507_26159# a_18371_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2725 net23 a_5324_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2726 vssd1 a_17107_4073# a_17114_3977# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2728 vssd1 a_3155_7663# net39 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2729 vccd1 _0839_ a_9779_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2731 a_23389_14191# a_23119_14557# a_23299_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2732 vccd1 _0319_ a_3983_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2733 a_9043_10089# _0700_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2734 a_6527_23439# _0755_ _0827_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X2735 a_15749_20719# _0464_ a_15667_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2736 _0462_ a_19255_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2737 vccd1 net51 temp1.capload\[11\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2739 vccd1 a_20947_3677# a_21115_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2740 a_13729_2223# a_13459_2589# a_13639_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2742 a_6538_5853# a_6265_5487# a_6453_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2745 a_16845_26703# cal_lut\[91\] a_16761_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2746 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2747 a_6182_22895# clknet_0_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
R7 temp1.capload\[13\].cap_53.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2749 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7636_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X2750 a_11371_27613# a_10589_27247# a_11287_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X2751 a_5687_4564# _0317_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2752 a_8197_3855# a_7663_3861# a_8102_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2754 a_11110_21807# _0665_ a_11020_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X2755 _0027_ a_25235_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2756 _0355_ a_25507_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2757 a_7888_32375# net10 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2758 a_17489_1685# a_17323_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2759 a_11711_10205# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2760 a_3171_26703# _0414_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2761 net21 a_4995_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2762 a_24861_6397# a_24591_6031# a_24771_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2763 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2764 _0415_ _0414_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2765 vccd1 net27 a_7387_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2766 a_18229_12559# _0017_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2768 a_10835_4161# _0290_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2769 a_27287_22173# a_26505_21807# a_27203_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2770 a_2497_14191# _0202_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2771 a_3817_7119# a_3479_7351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2772 a_1641_28500# _0825_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2774 vccd1 _0238_ a_24683_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2775 cal_lut\[18\] a_18907_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2777 _0312_ a_12535_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2779 a_20349_9839# _0505_ a_20267_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2780 a_6929_20719# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2781 _0603_ a_16035_6144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2782 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2783 a_12165_22671# _0664_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2784 a_14729_21269# a_14563_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2785 vssd1 a_8146_18796# dbg_result[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X2786 vccd1 a_8845_28023# _0408_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X2787 _0211_ a_9179_28309# a_8951_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2788 a_1951_26703# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X2789 a_2576_17271# net6 a_2504_17271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X2791 a_16889_22689# _0464_ a_16803_22689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2792 a_3885_21263# _0427_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X2793 vssd1 net32 a_21187_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2794 a_27774_12533# a_27606_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2795 cal_lut\[18\] a_18907_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R8 vssd1 net52 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2796 a_19820_15279# a_19421_15279# a_19694_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2797 a_23361_9985# _0658_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X2798 vccd1 a_15519_27791# a_15687_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2799 vssd1 _0221_ a_18519_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2800 vccd1 _0428_ a_1917_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2801 vccd1 a_13783_24148# _0009_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2802 _0360_ a_25875_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2803 a_17066_12559# _0602_ a_16986_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2804 _0497_ a_9126_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X2805 cal_lut\[62\] a_25439_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2806 cal_lut\[41\] a_15595_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2807 a_5583_14735# a_4885_14741# a_5326_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2808 vssd1 a_18291_9527# cal_lut\[106\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2809 a_14821_23445# a_14655_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2810 vccd1 a_22441_21237# _0639_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2811 cal_lut\[24\] a_20287_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2812 a_22270_1679# a_21997_1685# a_22185_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2813 vssd1 _0360_ a_26063_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2814 vssd1 a_6799_28853# a_6541_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X2815 vccd1 cal_lut\[57\] a_22891_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2816 a_26578_18655# a_26410_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2817 vccd1 cal_lut\[102\] a_18055_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2819 _0212_ a_6914_28111# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X2820 a_2931_17455# _0422_ a_2489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2821 vccd1 _0663_ _0669_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2822 vssd1 a_9907_6031# a_10075_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2823 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2824 vccd1 a_23355_23671# _0471_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X2825 _0047_ a_18519_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2826 a_7741_16367# _0001_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2827 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2828 a_7084_32143# a_6835_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2830 vssd1 a_25502_21781# a_25431_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X2831 a_8573_21263# _0434_ _0785_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2832 net30 a_3339_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2833 a_17677_23983# _0082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2834 vssd1 a_26835_18909# a_27003_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2835 a_16986_13647# _0599_ a_16737_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X2836 vccd1 cal_lut\[129\] a_11742_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2837 a_15541_9985# _0547_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X2839 a_14710_7775# a_14542_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2840 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2841 _0633_ a_21831_9408# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2843 a_8711_4943# a_7847_4949# a_8454_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2844 vssd1 a_5675_9295# a_5843_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2845 _0732_ _0715_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2846 vssd1 a_21759_2491# a_21717_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2847 vssd1 _0670_ a_9253_21601# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2848 a_17835_7637# a_18126_7937# a_18077_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2849 vccd1 cal_lut\[69\] a_25047_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2850 vssd1 cal_lut\[178\] a_15569_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2851 _0514_ a_17599_6039# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2852 vccd1 _0349_ a_24039_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2853 vssd1 a_24094_14709# a_24052_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2854 a_8532_31751# net11 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2855 vccd1 a_11581_21781# _0674_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2856 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2857 a_17257_5487# _0495_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2858 vssd1 dbg_result[2] a_14770_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2859 a_2000_26935# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2860 a_24846_23261# a_24407_22895# a_24761_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2861 vccd1 _0531_ a_20359_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2862 dbg_result[5] a_11366_28588# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2863 vssd1 _0544_ a_15909_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2864 vccd1 a_20322_9269# a_20249_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2866 _0223_ a_19664_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2867 vssd1 _0414_ _0746_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2869 _0296_ a_22240_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2870 vccd1 net33 a_21831_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2871 vccd1 _0435_ a_6646_21041# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X2872 a_25586_11293# a_25339_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X2873 vssd1 net46 a_19439_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2875 a_23481_23439# _0463_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X2876 _0024_ a_21095_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2877 vssd1 clknet_1_1__leaf_net67 net70 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2878 vccd1 cal_lut\[23\] a_18274_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2879 vssd1 a_7994_29535# a_7952_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2880 vssd1 clknet_1_0__leaf__0380_ a_5377_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2881 a_7741_6575# _0126_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2882 cal_lut\[111\] a_20747_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2883 a_17811_17999# a_17029_18005# a_17727_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2884 a_17536_10383# _0515_ a_17434_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2886 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2888 a_14611_11079# _0483_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2889 a_22291_7663# cal_lut\[159\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2890 vssd1 a_25295_21781# a_25302_22081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2891 a_7559_18909# a_7277_18543# a_7465_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X2893 a_25327_10383# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2894 a_23259_3133# a_23039_3145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2895 vccd1 _0266_ a_17691_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X2896 vssd1 a_28199_10107# a_28157_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2897 a_11705_10703# cal_lut\[39\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2898 a_19915_19087# dbg_result[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2899 vccd1 net25 a_11987_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2900 vccd1 _0514_ a_16127_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2901 a_26593_9839# a_25603_9839# a_26467_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2903 a_19694_4765# a_19255_4399# a_19609_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2904 vccd1 _0492_ a_11693_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2906 a_25962_11989# a_25755_11989# a_26138_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2907 vssd1 a_16069_22923# _0487_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X2908 a_20798_19997# a_20525_19631# a_20713_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2909 _0422_ a_1743_18259# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2910 vssd1 a_14151_11079# _0567_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2911 vccd1 a_5675_13469# a_5843_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2912 a_9638_4399# cal_lut\[134\] a_9548_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X2913 _0317_ a_5451_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2914 vssd1 a_23063_25437# a_23231_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2916 a_23189_4233# a_22199_3861# a_23063_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2918 vccd1 cal_lut\[32\] a_23201_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2919 vssd1 a_7410_17973# dbg_result[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2920 a_20345_16911# _0029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2921 _0539_ _0538_ a_19987_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.13 ps=1.26 w=1 l=0.15
X2922 vccd1 _0454_ a_18597_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2923 a_2805_30265# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2925 vssd1 a_2221_13255# _0412_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2926 _0150_ a_19439_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2927 vccd1 a_4647_12533# a_4563_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2928 vccd1 a_17930_24095# a_17857_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2929 a_16951_23439# a_16771_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2930 a_10562_19319# _0590_ a_10865_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X2931 a_9873_16617# _0702_ a_9749_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.235 ps=1.47 w=1 l=0.15
X2932 a_6458_20175# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2933 a_7111_10205# _0836_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2934 a_15519_27791# a_14655_27797# a_15262_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2935 vccd1 net42 a_26983_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2936 a_24551_5461# a_24835_5461# a_24770_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2937 a_18015_5639# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2938 vccd1 _0460_ a_22903_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2941 a_8504_16201# a_8105_15829# a_8378_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2942 vssd1 a_6429_28309# _0209_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2943 a_7652_18909# a_7111_18543# a_7559_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X2944 vssd1 temp_delay_last a_4027_16144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2945 vssd1 a_25439_7093# a_25397_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2946 a_13809_28879# a_13275_28885# a_13714_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2947 _0269_ a_17871_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X2949 a_4701_7663# a_4535_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2951 vccd1 a_5693_21781# _0758_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2952 vssd1 _0432_ _0779_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2954 a_10783_30511# net13 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2955 a_22270_23439# a_21831_23445# a_22185_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2956 dbg_result[2] a_8146_18796# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X2957 a_3005_17999# _0422_ a_2921_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2958 a_11597_14191# a_10607_14191# a_11471_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2959 a_3953_10761# a_3399_10601# a_3606_10660# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2960 vccd1 a_3848_24135# _0823_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2961 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd a_3056_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2962 a_26417_18231# _0246_ a_26580_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2963 a_10501_13879# cal_lut\[80\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X2964 a_6508_32375# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2965 vssd1 a_15262_29535# a_15220_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2966 a_15189_27791# a_14655_27797# a_15094_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2967 a_10129_3311# a_9963_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2969 a_18272_12265# _0605_ a_18170_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2970 a_10522_19631# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2971 vssd1 a_7407_12283# a_7365_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2972 vccd1 _0422_ a_3799_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2973 vccd1 clknet_1_0__leaf_io_in[0] a_1959_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2974 vssd1 a_22955_14709# a_22913_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2975 a_15737_14025# a_14747_13653# a_15611_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2976 a_11882_25321# _0730_ a_11579_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X2977 a_6823_14735# a_6375_14741# a_6729_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2978 a_6703_6549# a_6879_6549# a_6831_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X2979 a_3931_30006# a_3749_30006# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2980 vssd1 a_27774_15797# a_27732_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2981 a_6354_29789# a_6081_29423# a_6269_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2982 vccd1 net48 a_16219_25623# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2984 cal_lut\[165\] a_25439_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2985 vssd1 clknet_1_0__leaf_io_in[0] a_3615_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2986 vccd1 _0814_ a_5264_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X2987 a_2778_24527# temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2988 a_12160_18543# net16 a_11857_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X2989 a_27881_8751# a_26891_8751# a_27755_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2990 vssd1 _0773_ a_4224_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X2991 a_10589_27247# a_10423_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2992 a_9673_23047# _0717_ a_9836_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2995 a_2014_14709# a_1846_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2996 vccd1 a_23110_3044# a_23039_3145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2997 a_22247_9991# _0450_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2998 _0653_ a_10607_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2999 a_12502_17567# a_12334_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3001 vccd1 a_20303_26703# a_20471_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3002 a_3133_14191# a_2143_14191# a_3007_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3003 vccd1 net30 a_10607_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3004 vssd1 a_9551_2388# _0181_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3005 a_20889_2057# a_19899_1685# a_20763_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3006 a_5307_29789# a_4443_29423# a_5050_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3007 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3008 vccd1 a_20287_5755# a_20203_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3009 a_5779_8426# _0324_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3010 _0819_ _0557_ a_8853_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3012 vccd1 a_2823_15823# a_2991_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3013 vccd1 a_19977_14709# _0501_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3014 vssd1 a_25375_12167# cal_lut\[176\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3015 _0850_ a_10699_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3016 _0156_ a_19807_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3017 a_23377_8029# a_22843_7663# a_23282_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3018 vssd1 a_12759_17821# a_12927_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3019 _0025_ a_23763_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3020 vssd1 ctr\[1\] a_2221_13255# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3021 _0064_ a_19531_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3022 vccd1 a_24075_19087# a_24243_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3023 vccd1 a_15446_2741# a_15373_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3024 a_17746_6687# a_17578_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3025 vssd1 _0419_ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3026 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7084_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X3027 a_17669_15113# a_16679_14741# a_17543_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3028 vccd1 a_26107_8725# a_25931_8725# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X3030 vssd1 a_9687_29423# net9 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3031 vccd1 net44 a_21371_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3032 vssd1 _0812_ a_5573_29217# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3033 vssd1 a_23754_26980# a_23683_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3034 vccd1 a_20287_24501# a_20203_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3035 a_24099_12777# net36 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3036 a_20253_1679# _0150_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3037 a_17746_6687# a_17578_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3038 _0347_ a_26519_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X3039 _0460_ a_20451_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3040 a_20161_22351# _0064_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3041 vccd1 a_5751_14709# a_5667_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3042 a_16859_2045# cal_lut\[149\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X3043 a_8447_7338# _0308_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3044 a_9117_13353# cal_lut\[20\] a_9033_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3045 a_7188_19453# a_7157_19319# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X3046 vccd1 a_13459_17455# _0438_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3048 a_23723_25045# cal_lut\[86\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X3049 _0631_ _0630_ a_10247_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3050 a_5250_3855# a_4977_3861# a_5165_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3051 vccd1 a_21759_11195# a_21675_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3054 a_18291_16532# _0254_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3055 vccd1 a_23763_4943# _0476_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3057 net35 a_15812_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3058 _0467_ a_15370_19407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X3059 a_14637_1501# a_14103_1135# a_14542_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3060 a_23482_27069# a_23167_26935# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3062 a_4679_10615# a_4963_10601# a_4898_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3063 vccd1 _0231_ a_23395_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3064 vccd1 _0248_ a_27351_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3065 a_11601_3311# a_11435_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3067 a_25410_10901# a_25203_10901# a_25586_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3068 vssd1 a_8544_17429# _0433_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X3069 _0839_ a_4167_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3070 io_out[2] a_2511_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3071 a_22089_14741# a_21923_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3072 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3074 a_5099_10761# a_4970_10505# a_4679_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3075 a_14375_28701# a_14195_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3076 a_22937_23983# _0469_ a_22503_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3077 vccd1 cal_lut\[26\] a_23205_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X3078 a_4889_7663# _0142_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3079 a_24262_10383# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X3080 a_17007_29397# a_17298_29697# a_17249_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3083 a_13122_6147# _0299_ a_13040_6147# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3084 _0784_ ctr\[6\] a_4273_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X3085 vccd1 a_19303_18695# _0507_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3086 a_5346_10383# a_5099_10761# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3087 vssd1 _0358_ a_27351_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3088 a_21131_27791# a_20433_27797# a_20874_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3089 a_7273_3311# a_6283_3311# a_7147_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3090 a_9555_25847# _0720_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3091 vssd1 _0266_ a_15711_24833# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3094 _0145_ a_7571_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3095 a_15312_14025# a_14913_13653# a_15186_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3096 a_25339_10927# a_25203_10901# a_24919_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3097 vccd1 a_9559_26481# _0386_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3098 vccd1 _0775_ a_7853_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3099 vssd1 a_21970_18231# _0490_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X3101 a_24179_20541# a_23959_20553# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3102 a_21223_19997# a_20525_19631# a_20966_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3103 vccd1 net23 a_4811_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3104 vccd1 a_25439_24251# a_25355_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3105 _0711_ a_10915_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X3106 vccd1 a_19915_19087# _0443_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3109 a_16566_22173# a_16127_21807# a_16481_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3110 a_11705_8527# cal_lut\[123\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3111 _0631_ _0630_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X3112 a_20893_10927# a_20727_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3113 vssd1 _0850_ a_17875_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3114 _0498_ a_16757_7637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X3115 a_4714_23483# _0821_ a_4713_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X3117 a_7847_28992# ctr\[11\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3118 a_17417_22895# _0466_ a_16983_23047# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3119 vccd1 _0027_ a_25389_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3120 a_19421_5487# a_19255_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3121 vccd1 clknet_1_1__leaf_io_in[0] a_6927_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3123 a_8251_6941# a_7387_6575# a_7994_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3124 a_20296_13647# _0501_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X3125 a_19820_4399# a_19421_4399# a_19694_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3126 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_2504_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X3127 vccd1 a_25295_21781# a_25302_22081# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3129 a_19373_21835# _0454_ a_19287_21835# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3130 ctr\[0\] a_2439_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3131 vssd1 io_in[6] a_1407_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3132 vccd1 a_4663_10205# a_4831_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3133 vccd1 cal_lut\[24\] a_20482_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3134 _0014_ a_23671_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3135 a_13127_13469# a_12429_13103# a_12870_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3136 vssd1 _0264_ a_23763_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3137 a_20303_26703# a_19439_26709# a_20046_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3138 vssd1 _0728_ a_8093_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3139 vccd1 net25 a_14103_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3140 a_8377_8751# a_7387_8751# a_8251_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3141 a_3399_10601# clknet_1_0__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3142 _0222_ a_20963_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3143 vccd1 _0697_ a_9293_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3144 a_24770_13103# a_24455_13255# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3146 vssd1 a_14979_24148# _0094_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3147 a_23481_23439# _0466_ a_23683_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3149 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3150 vssd1 a_13847_9269# a_13805_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3151 a_24075_19087# a_23211_19093# a_23818_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3152 a_14825_7119# _0125_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3153 vssd1 a_9371_2741# _0367_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X3154 a_11943_8751# a_11723_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3155 vccd1 _0464_ a_15667_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3156 vccd1 a_2271_14735# a_2439_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3157 vccd1 cal_lut\[12\] a_20390_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3158 vccd1 cal_lut\[184\] a_13823_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3159 vccd1 cal_lut\[183\] a_11707_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3160 a_21675_10205# a_20893_9839# a_21591_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3162 vssd1 a_2209_25589# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X3163 vccd1 a_6706_5599# a_6633_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3164 a_22409_9839# _0452_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X3165 vssd1 _0280_ a_16035_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3166 vssd1 a_10746_10615# _0702_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X3168 a_4984_25615# _0801_ a_4893_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X3170 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3171 vssd1 _0532_ a_19865_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3173 a_6982_12533# a_6814_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3174 vssd1 a_2773_9991# _0837_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3177 vccd1 a_15193_15431# _0518_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X3178 a_19641_2589# a_19303_2375# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3179 a_1761_12559# _0200_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3180 a_10025_29257# a_9478_29001# a_9678_29156# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3181 a_12223_2741# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3183 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_5724_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X3184 vccd1 a_21155_26133# a_21162_26433# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3185 temp1.dac_vout_notouch_ net13 a_10692_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X3186 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3187 vccd1 _0269_ a_17875_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3188 a_21997_23445# a_21831_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3189 a_5639_23759# _0818_ a_5545_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3190 a_22373_23145# _0685_ a_22291_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3191 a_27847_17999# a_26983_18005# a_27590_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3192 vssd1 a_19303_17607# _0610_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X3193 vccd1 net27 a_6743_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3194 vccd1 _0364_ a_16955_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3195 a_15373_2767# a_14839_2773# a_15278_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3196 vssd1 _0160_ a_25941_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3197 a_9963_9001# cal_lut\[140\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X3198 _0795_ ctr\[7\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3199 a_20065_1685# a_19899_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3200 a_26210_9951# a_26042_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3201 a_14375_10205# a_14195_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3204 a_26283_8207# a_25419_8213# a_26026_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3205 a_3995_7497# a_3859_7337# a_3575_7351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3206 a_25339_10927# a_25210_11201# a_24919_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3207 a_27333_12565# a_27167_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3208 vccd1 _0681_ a_10229_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3209 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3211 a_27606_15823# a_27167_15829# a_27521_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3212 a_24731_6740# _0348_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3213 a_3607_25615# clknet_1_1__leaf_temp1.i_precharge_n temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X3214 vssd1 dbg_result[3] a_21997_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0619 ps=0.715 w=0.42 l=0.15
X3215 cal_lut\[5\] a_12099_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3216 vccd1 a_27595_13865# a_27602_13769# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3217 _0298_ a_19343_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X3218 a_26099_17821# a_25401_17455# a_25842_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3219 vccd1 a_8803_15823# a_8971_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3220 vccd1 a_7607_10383# a_7775_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3221 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3222 _0268_ a_18560_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X3223 a_10145_19203# _0628_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X3224 vssd1 _0594_ a_17565_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3225 a_17875_10383# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3227 vssd1 net37 a_23487_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3228 vccd1 _0815_ a_7840_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X3229 a_7691_6031# a_6909_6037# a_7607_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3231 vssd1 cal_lut\[45\] a_15569_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3232 vssd1 _0379_ a_2879_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3234 a_8377_13103# a_7387_13103# a_8251_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3235 a_16156_15823# _0540_ a_16054_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3236 vssd1 a_22431_7338# _0158_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3237 a_19439_7119# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3239 vssd1 a_23355_10615# _0696_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X3240 vssd1 a_7895_12778# _0019_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3241 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3242 _0336_ a_22471_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X3243 vssd1 a_8447_7338# _0126_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3244 vssd1 net44 a_21371_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3245 vssd1 net26 a_14379_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3246 vccd1 cal_lut\[38\] a_8947_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3247 vccd1 _0403_ a_6647_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3248 vssd1 a_9835_26703# _0385_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3249 vssd1 a_6674_16620# dbg_result[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X3250 a_9275_15444# _0256_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3252 cal_lut\[89\] a_18539_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3253 _0152_ a_22659_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3254 a_13913_2045# a_13643_1679# a_13823_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3255 a_11797_2045# a_11527_1679# a_11707_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3256 vssd1 a_20671_22351# a_20839_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3257 vssd1 clknet_1_1__leaf_io_in[0] a_7387_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3258 a_6729_17999# _0195_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3259 a_9390_14557# a_9117_14191# a_9305_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3260 vccd1 clknet_0_temp1.i_precharge_n a_3882_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3261 a_22770_21263# _0637_ a_22690_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3263 a_13241_5633# _0568_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X3264 vccd1 cal_lut\[150\] a_16340_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X3265 vccd1 cal_lut\[109\] a_23481_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X3266 a_15170_10357# a_15002_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3267 vssd1 a_6955_23671# _0753_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3268 vccd1 a_4032_25847# _0829_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3269 a_23535_17143# a_23631_17143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3270 a_9344_6575# cal_lut\[127\] a_9224_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3271 a_22659_8751# cal_lut\[153\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3272 a_24459_8181# a_24635_8513# a_24587_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3274 vccd1 cal_lut\[69\] a_23811_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3275 a_11609_21379# _0670_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3277 a_20114_13647# _0533_ a_19865_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3279 a_5555_24233# _0414_ _0773_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3280 a_7853_22351# _0434_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3281 cal_lut\[6\] a_12927_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3282 a_8887_1679# a_8105_1685# a_8803_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3284 a_20273_18543# cal_lut\[53\] a_20201_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3285 a_6722_3677# a_6449_3311# a_6637_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3286 _0334_ a_18975_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X3287 vssd1 _0488_ a_15391_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3288 a_19421_15279# a_19255_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3289 vccd1 _0174_ a_26861_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3290 vssd1 a_13783_24148# _0009_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3291 vssd1 cal_lut\[60\] a_21136_23145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3292 a_23303_18909# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3293 vccd1 a_22151_3073# a_21975_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X3294 a_5170_10660# a_4963_10601# a_5346_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3295 a_12219_17130# _0845_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3296 vssd1 cal_lut\[143\] a_6277_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3297 a_27498_8863# a_27330_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3298 a_21709_26159# a_21162_26433# a_21362_26133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3299 a_2366_25615# ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X3300 a_9831_24501# _0720_ a_10262_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X3301 a_6955_23671# _0752_ a_7101_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3302 vccd1 ctr\[12\] a_6737_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X3303 vccd1 net20 a_21831_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3305 a_10843_2197# a_11019_2197# a_10971_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3306 a_23481_10703# _0506_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X3307 vssd1 a_6674_16620# dbg_result[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X3309 vccd1 _0352_ a_26983_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3310 a_16297_10927# _0101_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3311 a_25014_23007# a_24846_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3312 vssd1 a_1407_15823# net7 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3313 temp1.capload\[7\].cap.Y net62 a_1493_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3314 vccd1 a_5897_28335# a_6003_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X3315 a_2973_19407# _0411_ a_2023_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3316 vccd1 _0588_ a_11765_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
X3317 vccd1 a_28031_17821# a_28199_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3318 a_2000_29111# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3319 vccd1 a_23823_20393# a_23830_20297# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3320 a_8491_18319# _0517_ a_8645_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3321 a_27422_17999# a_27149_18005# a_27337_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3322 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3323 a_2931_22325# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3324 _0670_ _0666_ a_10121_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X3325 vssd1 _0769_ a_5181_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X3326 a_19303_17607# _0454_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3327 a_17814_13647# _0595_ a_17565_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3328 _0354_ a_25783_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X3329 vssd1 a_15979_3855# a_16147_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3330 a_7239_12559# a_6541_12565# a_6982_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3331 a_4609_29423# a_4443_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3332 net31 a_16640_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3333 vssd1 _0349_ a_24039_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3334 a_16681_13353# _0600_ a_16585_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3336 _0070_ a_26063_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3337 a_7457_25071# _0724_ a_7373_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3338 a_11348_21807# _0672_ a_10857_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3339 vssd1 a_4663_10205# a_4831_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3341 vssd1 net12 a_10423_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3343 vccd1 a_10827_1679# a_10995_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3344 vssd1 a_22863_27765# a_22821_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3345 a_15569_25981# a_15299_25615# a_15479_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3346 _0424_ a_2722_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3347 vccd1 a_12943_1679# a_13111_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3348 vccd1 a_16179_29397# _0218_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3349 vssd1 a_10459_15823# a_10627_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3350 vssd1 a_27847_7119# a_28015_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3351 a_18907_19407# dbg_result[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X3352 vssd1 a_2010_24759# _0416_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0878 ps=0.92 w=0.65 l=0.15
X3353 a_23217_15279# cal_lut\[72\] a_23145_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3354 a_6633_5853# a_6099_5487# a_6538_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3355 vssd1 cal_lut\[113\] a_18605_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3356 a_9558_14303# a_9390_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3357 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3358 a_4897_27247# a_4705_27552# _0207_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3359 vccd1 a_25439_23163# a_25355_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3360 a_14269_7663# a_14103_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3361 a_20893_10927# a_20727_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3362 vssd1 _0359_ a_27903_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3363 a_17739_21959# _0452_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3364 vssd1 _0557_ a_10247_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3365 vssd1 cal_lut\[146\] a_10141_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3366 a_18100_17027# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3367 a_9749_16617# _0519_ a_9677_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X3368 vssd1 a_24099_4073# a_24106_3977# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3369 _0863_ a_13144_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3370 _0561_ a_19426_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X3371 a_27701_15823# a_27167_15829# a_27606_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3372 vccd1 net50 temp1.capload\[10\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3373 _0114_ a_20727_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3374 vccd1 ctr\[8\] a_5547_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3375 net43 a_22291_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X3376 a_27774_9951# a_27606_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3377 a_7607_10383# a_6743_10389# a_7350_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3378 vssd1 a_7534_27359# a_7492_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3379 vssd1 _0721_ _0748_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3380 a_6791_4074# _0315_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3381 a_16005_8573# cal_lut\[180\] a_15933_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3382 a_7618_26935# dec1.i_ones a_7921_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3383 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3384 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3385 a_13691_28500# _0224_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3386 vssd1 dec1.i_ones a_7618_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3387 vccd1 a_20046_26677# a_19973_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3388 a_12263_26525# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3390 vccd1 a_10385_23413# _0681_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3391 a_9201_3829# _0502_ a_9358_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3392 net36 a_24499_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3393 a_19084_17289# a_18685_16917# a_18958_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3394 a_27057_8751# a_26891_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3396 vccd1 a_21591_2589# a_21759_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3397 vccd1 net19 a_21003_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3398 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3399 vccd1 a_7607_2589# a_7775_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3401 a_2596_30511# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X3402 a_24653_12937# a_24106_12681# a_24306_12836# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3403 a_6890_3423# a_6722_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3404 vccd1 _0476_ a_21983_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3405 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3406 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3407 vssd1 a_17543_9295# a_17711_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3408 a_7277_10383# a_6743_10389# a_7182_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3409 a_21970_18231# _0489_ a_22273_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3410 a_13027_1679# a_12245_1685# a_12943_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3411 cal_lut\[93\] a_14583_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3412 vssd1 net48 a_12723_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3413 vccd1 _0839_ a_6467_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3415 a_3891_22057# _0737_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X3416 vccd1 _0057_ a_24377_20553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3417 vccd1 cal_lut\[27\] a_23903_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3418 a_5971_15253# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3420 a_17857_3311# a_17691_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3421 a_13091_9001# _0565_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3422 a_7921_11293# a_7387_10927# a_7826_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3423 a_21291_26159# a_21155_26133# a_20871_26133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3424 _0064_ a_19531_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3425 vssd1 _0421_ a_3525_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3426 vccd1 cal_lut\[84\] a_17739_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3428 vssd1 a_19865_13621# _0534_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X3429 vccd1 a_24306_12836# a_24235_12937# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3430 a_7389_23759# _0750_ a_6955_23671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3431 vccd1 a_15193_14343# _0852_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X3432 a_17094_20407# _0586_ a_17397_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3433 _0510_ a_22875_9867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3434 vssd1 a_25042_13077# a_24971_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3435 a_11120_28853# net14 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3436 vccd1 a_25003_24833# a_24827_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X3438 vccd1 a_6699_13268# _0018_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R9 vssd1 net59 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3439 a_25397_23983# a_24407_23983# a_25271_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3440 a_18341_8573# cal_lut\[113\] a_18269_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3441 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3442 vccd1 clknet_1_0__leaf_io_in[0] a_4811_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3443 vccd1 a_4831_10107# a_4747_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3444 a_9397_6031# _0127_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3447 vccd1 net48 a_17875_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3449 a_5547_26409# ctr\[9\] a_5801_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3450 a_8979_18543# _0517_ _0680_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3451 a_18774_13647# a_18335_13653# a_18689_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3452 a_24861_20719# a_24591_21085# a_24771_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3453 a_15009_27791# _0091_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3454 a_22151_3073# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3456 vccd1 a_9933_19061# _0630_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3457 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3458 a_14103_18793# _0447_ a_14353_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3460 a_16679_1501# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3462 a_7239_17999# a_6375_18005# a_6982_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3463 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3464 a_18187_25437# a_17489_25071# a_17930_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3465 a_5998_20495# _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X3466 _0194_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3467 vssd1 a_4066_7396# a_3995_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3469 a_13148_10499# cal_lut\[97\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X3470 _0414_ a_2419_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3471 a_11895_16367# _0609_ _0626_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3472 a_18873_16911# _0028_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3473 vssd1 clknet_0_temp1.i_precharge_n a_1753_26133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3475 a_19973_22357# a_19807_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3476 _0544_ a_15943_7232# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3477 vccd1 net52 temp1.capload\[12\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3478 a_25849_21807# a_25302_22081# a_25502_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3479 vccd1 _0058_ a_22813_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
R10 net51 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3482 vccd1 _0474_ a_22875_9867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3483 vssd1 cal_lut\[58\] a_21872_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3484 a_9447_8207# a_8749_8213# a_9190_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3485 cal_lut\[13\] a_21851_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3486 a_17314_4132# a_17107_4073# a_17490_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3487 a_18416_12015# cal_lut\[185\] a_17841_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3488 a_18709_19631# cal_lut\[28\] a_18637_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3490 vssd1 net8 a_12623_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X3491 a_7791_27613# a_6927_27247# a_7534_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3492 a_16209_20541# _0454_ a_16127_20288# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3493 _0495_ a_13714_19407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3494 vssd1 _0481_ a_12233_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3495 a_10126_13469# a_9687_13103# a_10041_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3496 vccd1 _0591_ a_8573_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3497 _0440_ a_14156_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3498 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3499 vccd1 _0354_ a_26155_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3501 vccd1 ctr\[12\] a_9563_28487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3502 vssd1 a_16737_12533# _0604_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X3503 vccd1 _0809_ a_4843_15307# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3504 cal_lut\[81\] a_11639_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3505 vssd1 net40 a_11711_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3506 a_21591_4765# a_20727_4399# a_21334_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3507 a_8711_4943# a_8013_4949# a_8454_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3508 cal_lut\[25\] a_22403_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3510 a_23075_27247# a_22855_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3511 cal_lut\[129\] a_11639_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3512 a_11151_29423# net13 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X3513 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3514 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3515 a_7461_27613# a_6927_27247# a_7366_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3516 cal_lut\[165\] a_25439_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3517 a_14611_11079# _0440_ a_14845_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3518 vccd1 cal_lut\[76\] a_17135_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3519 a_13445_23439# _0009_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3521 vccd1 _0433_ _0520_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3522 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3523 vssd1 a_23811_27412# _0055_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3524 a_21810_22173# a_21537_21807# a_21725_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3525 a_20798_19997# a_20359_19631# a_20713_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3526 vssd1 _0383_ _0194_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3527 vssd1 a_26417_18231# _0247_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3529 vssd1 a_15779_13621# a_15737_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3531 vccd1 _0413_ a_2419_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3532 a_12978_25437# a_12539_25071# a_12893_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3533 vssd1 _0432_ a_5996_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3535 a_5412_19783# _0736_ a_5554_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3536 vccd1 a_19862_24501# a_19789_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3537 vssd1 _0527_ a_20417_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3538 vccd1 a_27774_15797# a_27701_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3539 a_18647_28879# a_17783_28885# a_18390_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3540 a_15904_25589# net47 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3541 a_13969_18218# _0539_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3542 a_16718_17705# _0610_ a_16404_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X3543 a_12863_14954# _0275_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3544 a_19303_16519# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3545 _0305_ a_11247_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X3546 vssd1 a_13882_28853# a_13840_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3547 vccd1 _0287_ a_18519_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3548 a_6541_12565# a_6375_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3549 _0710_ _0674_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3550 a_17739_21959# _0531_ a_17973_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3551 net44 a_17875_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3552 a_21081_10927# _0103_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3553 vssd1 a_10380_19783# _0667_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3555 a_8378_1679# a_7939_1685# a_8293_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3556 a_5013_24825# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3557 a_7159_11092# _0374_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3558 a_12702_13469# a_12263_13103# a_12617_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3559 a_6914_28111# _0390_ a_6745_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X3561 vssd1 clknet_1_1__leaf__0380_ a_9319_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X3562 vccd1 a_15904_25589# net45 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3564 a_16484_7663# cal_lut\[150\] a_15909_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3565 a_6607_9514# _0322_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3566 a_23765_10703# _0509_ a_23355_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3567 a_11527_10383# _0496_ a_11705_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3569 vccd1 _0531_ a_21923_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3570 vccd1 a_14250_15797# a_14177_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3571 vssd1 a_4663_9117# a_4831_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3572 vssd1 a_17711_14709# a_17669_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3573 a_2071_11791# _0389_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X3575 _0344_ a_23943_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X3576 vccd1 a_12743_26677# a_12659_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3577 a_26203_6250# _0346_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3578 vccd1 _0263_ a_22291_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3579 vccd1 a_16187_23671# _0482_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3580 cal_lut\[79\] a_9155_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3582 a_20429_29257# a_19439_28885# a_20303_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3586 vccd1 a_7994_11039# a_7921_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3587 vssd1 net45 a_18795_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3588 vssd1 a_12815_20719# _0446_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3589 _0426_ _0421_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3590 a_21292_25071# a_20893_25071# a_21166_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3591 vssd1 _0299_ a_6637_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3592 a_6187_8029# a_6007_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3593 a_6779_29789# a_6081_29423# a_6522_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3594 vssd1 ctr\[4\] a_5643_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3595 vssd1 _0472_ a_16925_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3596 a_23124_11791# _0456_ a_22633_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3597 vssd1 cal_lut\[56\] a_22837_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3598 vccd1 a_8419_16635# a_8335_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3599 a_1769_8527# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3600 a_16933_10927# a_15943_10927# a_16807_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3601 a_19763_4074# _0298_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3602 a_6354_29789# a_5915_29423# a_6269_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3604 a_26318_16733# a_26045_16367# a_26233_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3606 vccd1 a_8971_22895# _0725_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X3607 vccd1 a_9319_26159# a_9671_26481# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.229 ps=1.36 w=0.64 l=0.15
X3609 a_27732_11849# a_27333_11477# a_27606_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3610 vccd1 a_15043_24501# a_14959_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3611 a_3759_21495# net21 a_4087_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3612 a_9305_1135# _0181_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3613 a_4897_20969# _0427_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X3614 a_20407_16519# net18 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3615 a_10055_8029# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3616 a_15189_19631# a_15023_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3617 _0162_ a_26799_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3619 a_23361_9985# _0656_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X3620 vccd1 _0445_ a_16771_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3621 a_15812_9269# net38 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3622 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3623 vssd1 a_14155_29397# _0224_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X3624 vccd1 _0838_ a_4167_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3625 vssd1 a_21334_11039# a_21292_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3626 a_9844_29967# a_9595_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X3627 vssd1 a_5179_14191# _0811_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3628 a_11287_27613# a_10423_27247# a_11030_27383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3629 vccd1 a_26451_8181# a_26367_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3630 a_23351_21959# _0531_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3631 a_22740_10703# cal_lut\[15\] a_22165_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3632 a_8767_11471# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3633 a_19329_25615# a_18795_25621# a_19234_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3634 a_24955_24893# cal_lut\[62\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X3635 _0568_ a_12539_5056# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3636 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3637 vccd1 a_15687_23413# a_15603_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3638 a_24573_22895# a_24407_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3639 vccd1 a_24823_15444# _0068_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3640 a_7465_18543# _0194_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X3641 vccd1 _0333_ a_16311_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3643 a_10294_11445# a_10126_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3644 a_21258_14557# a_20985_14191# a_21173_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3645 a_8096_31849# a_7847_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X3646 a_5993_16367# _0193_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3647 a_18140_13967# cal_lut\[77\] a_17565_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3648 a_27521_9839# _0170_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3649 _0400_ a_5864_26819# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X3650 vccd1 a_1407_4399# net1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3651 a_18222_28879# a_17949_28885# a_18137_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3652 vssd1 _0225_ a_14747_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3653 a_17117_27023# cal_lut\[43\] a_16679_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3654 vssd1 _0558_ a_19426_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X3655 a_17490_3855# a_17243_4233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3656 cal_lut\[146\] a_8879_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3657 vccd1 _0836_ a_12171_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3658 vccd1 a_18739_12559# a_18907_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3659 a_17470_2335# a_17302_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3660 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3661 dbg_result[2] a_8146_18796# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X3662 a_10046_9001# cal_lut\[122\] a_9963_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3663 vssd1 cal_lut\[17\] a_17088_12265# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3666 a_20963_15797# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3667 _0204_ a_4487_13077# a_4259_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3668 vssd1 a_18739_12559# a_18907_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3669 vccd1 net46 a_19255_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3670 a_23201_23145# _0468_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3671 a_23443_20407# a_23539_20407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3672 a_13882_4917# a_13714_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3673 a_11509_13353# cal_lut\[81\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3674 a_10402_1679# a_9963_1685# a_10317_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3675 vccd1 net23 a_7387_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3676 a_22109_17027# _0686_ a_22013_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3677 vccd1 _0290_ a_11067_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3678 a_16390_5487# _0616_ a_16636_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X3679 a_15023_22464# cal_lut\[93\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3680 a_2372_25935# _0801_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X3681 a_5179_8207# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3682 vssd1 net20 a_17993_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3683 vssd1 net10 a_7839_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X3684 a_25581_18377# a_24591_18005# a_25455_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3685 a_12337_14191# a_12171_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3687 vccd1 a_20119_15645# a_20287_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3688 vssd1 _0622_ a_17105_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X3689 vccd1 net40 a_13091_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3690 vccd1 a_6890_3423# a_6817_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3691 a_8397_24527# _0714_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X3692 a_8021_22895# _0748_ a_7939_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3693 a_9142_19631# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3694 _0867_ a_20400_15939# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3695 vssd1 a_22438_23413# a_22396_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3697 vccd1 a_7534_27359# a_7461_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3698 _0311_ a_11660_5059# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X3699 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3700 _0679_ _0678_ a_11422_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X3701 vccd1 _0411_ a_3575_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X3702 a_3990_27574# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3703 a_24793_5853# a_24455_5639# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3704 vccd1 a_14151_5652# _0118_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3705 vccd1 _0440_ a_14163_8903# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3706 vccd1 _0352_ a_24867_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3707 cal_lut\[31\] a_22403_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3708 vccd1 a_3995_18793# _0759_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3709 vssd1 clknet_1_1__leaf_io_in[0] a_6927_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3710 a_22339_27399# a_22435_27221# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3711 vssd1 cal_lut\[171\] a_27253_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3713 a_9034_6575# cal_lut\[145\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X3714 a_20900_12879# cal_lut\[114\] a_20325_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X3715 vssd1 net11 a_9779_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3716 vssd1 a_1464_23957# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.265 pd=1.47 as=0.091 ps=0.93 w=0.65 l=0.15
X3717 _0438_ a_13459_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3718 a_1673_16911# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3719 vssd1 dbg_result[3] a_12815_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3720 a_20937_15101# _0443_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X3721 a_13139_7351# net17 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3722 vccd1 a_20579_8029# a_20747_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3723 a_4733_16367# ctr\[3\] _0193_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3724 a_10853_8751# cal_lut\[141\] a_10781_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3725 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4988_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X3726 vccd1 _0483_ a_15023_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3727 vccd1 a_12815_20719# _0446_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3728 vssd1 _0370_ a_11987_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3729 vssd1 net25 a_14103_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3730 vssd1 _0472_ a_15637_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3732 a_6987_24233# _0751_ _0752_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X3733 a_15624_23145# _0645_ a_15522_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X3734 a_18637_18543# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X3735 vssd1 a_19862_5599# a_19820_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3736 a_21555_13469# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3737 vssd1 a_8419_9019# a_8377_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R11 net57 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3739 vccd1 net22 a_1917_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3740 _0383_ a_6979_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3741 _0452_ a_20690_18517# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X3743 a_3154_19881# a_3112_19783# a_3072_19637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3744 a_22523_5175# _0451_ a_22757_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3746 a_23539_20407# a_23823_20393# a_23758_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3747 vssd1 cal_lut\[24\] a_20400_15939# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3748 a_6244_25045# _0750_ a_6464_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3749 a_13403_25437# a_12539_25071# a_13146_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3751 vccd1 a_14153_20884# net17 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3753 a_26123_14165# net37 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3754 a_17727_17999# a_16863_18005# a_17470_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3755 a_26111_12015# a_25891_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3756 a_11195_28701# a_10497_28335# a_10938_28471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X3757 a_13882_4917# a_13714_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3759 a_8504_2057# a_8105_1685# a_8378_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3760 vccd1 _0514_ a_15483_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3761 a_2281_23983# _0414_ a_1464_23957# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3762 _0422_ a_1743_18259# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X3763 a_4951_7338# _0325_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3764 a_8299_32143# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X3765 a_3990_27247# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3766 a_17489_23983# a_17323_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3767 a_5142_7775# a_4974_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3769 a_15370_28879# a_14931_28885# a_15285_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3770 a_6632_16367# a_5639_16367# a_6503_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X3771 vssd1 _0491_ _0492_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3772 a_11895_16367# _0519_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3773 vssd1 _0418_ a_3327_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0894 ps=0.925 w=0.65 l=0.15
X3775 a_3730_19407# _0742_ a_3435_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X3776 vssd1 a_21155_26133# a_21162_26433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3778 vccd1 net1 a_13367_10391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
R12 vssd1 net58 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3780 a_13073_25437# a_12539_25071# a_12978_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3781 a_3115_10615# a_3399_10601# a_3334_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3782 _0259_ a_16951_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X3783 a_5841_19605# _0737_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3784 _0466_ a_17999_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X3785 vssd1 a_7239_7119# a_7407_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3786 vssd1 a_24823_11079# cal_lut\[177\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3788 a_4140_31849# a_3891_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X3789 a_17397_17999# a_16863_18005# a_17302_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3790 vssd1 a_24099_12777# a_24106_12681# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3791 vccd1 a_13403_23261# a_13571_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3792 a_20257_5309# _0441_ a_20175_5056# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3793 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3794 a_12134_7093# a_11966_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3795 a_16187_23671# _0481_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3796 vccd1 a_17739_21959# _0553_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3798 a_24846_24349# a_24573_23983# a_24761_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3800 a_7277_6031# a_6743_6037# a_7182_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3801 vccd1 _0863_ a_23579_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3802 cal_lut\[129\] a_11639_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3803 vssd1 net8 a_10783_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X3804 _0749_ _0732_ a_10883_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3805 temp1.dac_vout_notouch_ net14 a_9844_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X3806 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3808 a_27521_11471# _0171_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3809 a_22903_21959# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3810 vssd1 _0728_ a_8571_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X3811 a_5915_21263# ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X3812 a_8539_2986# _0367_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3813 vccd1 _0514_ a_15299_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3814 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3815 a_2741_24135# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X3816 _0673_ a_11191_19659# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3817 vssd1 a_5050_29535# a_5008_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3819 a_27253_10749# a_26983_10383# a_27163_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3820 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3821 vssd1 net26 a_11527_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3822 vssd1 a_13679_9295# a_13847_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3823 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8096_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X3824 vccd1 _0266_ a_16955_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X3826 a_8017_3855# _0132_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3827 a_13403_23261# a_12705_22895# a_13146_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3828 vssd1 _0423_ a_3057_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3829 a_3796_16189# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.104 ps=1 w=0.42 l=0.15
X3830 _0208_ a_4981_28940# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X3831 a_2447_19087# _0745_ a_2023_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3833 cal_lut\[21\] a_10719_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3834 vssd1 a_20303_26703# a_20471_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3835 cal_lut\[152\] a_22863_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3836 a_15903_3285# a_16079_3285# a_16031_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3837 a_12097_23983# _0708_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3838 vssd1 a_2823_15823# a_2991_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3839 vccd1 a_2750_14303# a_2677_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3840 cal_lut\[14\] a_23139_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3842 a_2695_20969# _0414_ _0419_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X3843 a_22642_19997# a_22395_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3844 a_16955_20719# cal_lut\[42\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3845 a_13415_20884# _0883_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3846 vccd1 _0850_ a_17875_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3848 a_9949_15823# _0003_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3849 a_4613_5487# _0136_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3850 vccd1 a_17187_18708# _0076_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3851 vccd1 a_22523_2999# cal_lut\[153\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3852 a_6716_31849# a_6467_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X3853 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3854 a_5938_22671# _0759_ a_5643_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X3855 _0069_ a_25327_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3856 vccd1 cal_lut\[20\] a_9131_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3858 a_20022_19881# _0222_ a_19940_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3859 a_17691_9117# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3860 a_6940_12015# a_6541_12015# a_6814_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3862 vccd1 cal_lut\[177\] a_22247_9991# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3864 _0429_ _0422_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3865 a_13905_26703# _0092_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3866 a_19421_15279# a_19255_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3867 a_20860_20969# _0872_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3868 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10028_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X3869 a_21166_2589# a_20893_2223# a_21081_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3871 a_20848_13353# _0526_ a_20746_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3872 cal_lut\[60\] a_21391_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3873 a_17187_18708# _0253_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3874 a_15093_7663# a_14103_7663# a_14967_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3875 vssd1 _0711_ _0730_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3876 a_24034_12925# a_23719_12791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3877 a_10037_19631# _0668_ a_9953_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3878 a_7182_2589# a_6909_2223# a_7097_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3879 a_10528_2057# a_10129_1685# a_10402_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3880 a_20154_8029# a_19715_7663# a_20069_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3881 vccd1 a_24683_14191# _0352_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3883 vccd1 a_13459_17455# _0438_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3885 a_9988_5487# cal_lut\[128\] a_9868_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3886 vssd1 _0590_ _0591_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3888 a_20499_8439# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3889 a_14729_10389# a_14563_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3890 a_16859_28879# a_16679_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3891 vccd1 a_21235_9514# _0104_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3892 _0748_ dec1.i_ones a_9235_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X3894 _0193_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3895 temp1.dac_vout_notouch_ net14 a_9864_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X3896 a_23305_16367# _0475_ a_22895_16519# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3898 a_25962_20452# a_25762_20297# a_26111_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3899 vssd1 a_10570_7093# a_10528_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3902 vccd1 a_5199_27765# a_5115_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3903 vccd1 _0206_ a_6437_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3904 _0802_ a_4984_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3905 vssd1 a_11674_15391# a_11632_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3906 cal_lut\[22\] a_13295_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3908 vssd1 temp1.i_precharge_n a_2778_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3910 vssd1 clknet_1_0__leaf_io_in[0] a_4719_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3911 a_9496_31375# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X3912 vssd1 a_18111_25589# net46 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3913 cal_lut\[116\] a_23231_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3914 a_24761_8751# _0164_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3915 a_20322_9269# a_20154_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3916 a_20039_18695# _0459_ a_20273_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3917 a_10677_20719# _0673_ a_10331_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3919 a_19435_3677# a_19255_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3920 vssd1 cal_lut\[46\] a_16904_25321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3921 a_7256_21237# _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3922 a_13375_18543# dbg_result[3] a_13291_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0567 ps=0.69 w=0.42 l=0.15
X3923 a_8108_25615# _0749_ a_7853_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3924 a_5545_23759# _0819_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X3925 a_18681_3311# a_17691_3311# a_18555_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3926 vssd1 _0444_ a_20256_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X3927 vccd1 cal_lut\[21\] a_11707_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3928 vssd1 ctr\[11\] a_7618_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3929 vccd1 a_25931_8725# _0350_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3930 a_21133_18543# dbg_result[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.213 ps=1.3 w=0.65 l=0.15
X3932 a_4818_25071# _0747_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3934 a_14776_9295# _0562_ a_14674_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3935 a_7826_16733# a_7387_16367# a_7741_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3936 a_9558_14303# a_9390_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3937 a_26203_6250# _0346_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3938 vccd1 a_14151_4564# _0131_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3939 a_9431_25071# _0714_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3940 a_11029_17429# a_11199_17607# a_11157_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3941 a_21978_16479# a_21810_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3942 a_17762_24349# a_17323_23983# a_17677_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3944 ctr\[10\] a_6947_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3945 a_6799_28853# ctr\[9\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3946 a_11324_28335# a_10331_28335# a_11195_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X3948 _0062_ a_24683_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3949 vccd1 cal_lut\[106\] a_15163_9527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3950 a_10443_25321# _0729_ a_10347_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X3951 a_13146_25183# a_12978_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3952 vccd1 a_14139_4943# a_14307_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3954 a_12407_10901# a_12698_11201# a_12649_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3955 vssd1 net9 a_11527_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3956 a_15299_3677# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3958 a_27755_9117# a_26891_8751# a_27498_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3959 vssd1 a_3606_10660# a_3535_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3960 vssd1 cal_lut\[172\] a_27161_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3961 vssd1 a_2287_22325# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3962 a_25389_19631# a_24835_19605# a_25042_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3964 a_10221_13469# a_9687_13103# a_10126_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3967 vssd1 a_28015_7093# a_27973_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3968 a_7741_10927# _0037_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3969 vssd1 net10 a_7387_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3970 vccd1 a_13146_25183# a_13073_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3971 a_16753_13353# _0604_ a_16681_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3972 vssd1 a_20775_14967# _0527_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X3973 a_25042_13077# a_24835_13077# a_25218_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3974 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4140_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X3976 a_25375_12167# a_25471_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3979 a_5508_24501# _0431_ a_5900_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3980 a_3794_7485# a_3479_7351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3981 vccd1 a_15623_26324# _0045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3982 a_5249_5487# a_4259_5487# a_5123_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3984 vssd1 net35 a_20727_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3985 a_15262_29535# a_15094_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3986 vssd1 a_15538_17567# a_15496_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3987 a_23926_14735# a_23487_14741# a_23841_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3988 vssd1 a_21591_2589# a_21759_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3989 a_8013_4949# a_7847_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3990 vssd1 a_4771_4917# _0320_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X3991 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_1775_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3992 a_23899_25045# _0237_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3993 a_3882_16911# net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3994 a_18029_16201# a_17482_15945# a_17682_16100# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3995 a_15078_7093# a_14910_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3996 a_24846_9117# a_24407_8751# a_24761_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3997 a_4222_12533# a_4054_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3998 vccd1 ctr\[10\] a_7847_28992# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4000 a_22983_15431# _0531_ a_23217_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4001 vssd1 _0529_ _0539_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.0878 ps=0.92 w=0.65 l=0.15
X4002 a_10761_24893# _0682_ a_10689_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4003 a_19672_20969# _0559_ a_19570_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X4004 vccd1 a_27203_22173# a_27371_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4005 a_23117_4943# _0476_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4007 a_10362_5059# _0299_ a_10280_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4008 a_3334_10749# a_2947_10615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4009 a_23079_17607# _0479_ a_23407_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4010 a_13564_12937# a_13165_12565# a_13438_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4011 vccd1 _0481_ a_10699_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4012 a_18475_18695# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4014 a_25139_15101# cal_lut\[68\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X4016 vssd1 a_17560_4917# _0441_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4017 vssd1 _0483_ a_15453_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4018 vssd1 _0319_ a_3983_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4019 vssd1 _0287_ a_18519_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4021 _0597_ a_15943_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4022 a_12075_18793# _0556_ a_11857_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4023 vccd1 a_14131_13879# _0575_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4024 vssd1 net24 a_6099_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4025 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4026 a_27530_14013# a_27215_13879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4027 vssd1 a_17711_9269# a_17669_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4028 a_7159_11092# _0374_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4029 vssd1 cal_lut\[40\] a_14604_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 _0111_ a_18519_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4032 a_14103_27497# _0487_ a_14185_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4034 vccd1 net7 a_1773_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X4035 a_24499_22351# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4037 a_11931_15645# a_11067_15279# a_11674_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4038 a_24846_23261# a_24573_22895# a_24761_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4039 a_22466_19605# a_22259_19605# a_22642_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4040 vssd1 a_20579_8029# a_20747_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4041 vccd1 net29 a_14563_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4042 vssd1 a_4584_24759# _0799_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4043 a_3075_24305# clknet_1_0__leaf_temp1.i_precharge_n a_2563_23957# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X4044 vccd1 net72 a_5460_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4046 a_19255_7663# cal_lut\[144\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4047 a_4889_7663# _0142_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4048 vccd1 a_7407_12283# a_7323_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4049 vssd1 a_28031_10205# a_28199_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4051 vccd1 a_10719_13371# a_10635_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4052 a_11142_23983# _0681_ _0708_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X4053 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6716_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X4054 vssd1 a_8803_15823# a_8971_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4055 vccd1 a_23063_25437# a_23231_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4056 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4057 vccd1 _0216_ a_23211_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4058 a_10871_27613# a_10423_27247# a_10777_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4060 a_18129_6575# a_17139_6575# a_18003_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4061 a_23833_7663# a_22843_7663# a_23707_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4062 a_18369_18337# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4063 vssd1 _0839_ _0193_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4064 a_17381_15425# _0553_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4065 a_16823_4087# a_17114_3977# a_17065_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4066 a_15335_7119# a_14637_7125# a_15078_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4067 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd a_1952_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X4068 a_5444_21807# ctr\[3\] a_5141_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X4069 a_13241_5633# _0566_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X4070 vccd1 a_20407_16519# _0540_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4071 a_21683_14557# a_20985_14191# a_21426_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4072 a_2972_14013# ctr\[3\] a_2866_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4073 vccd1 a_15427_10383# a_15595_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4074 vccd1 _0372_ a_17231_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4075 vccd1 _0505_ a_15023_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4076 a_23818_19061# a_23650_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4077 cal_lut\[135\] a_5843_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4078 vssd1 clknet_0_io_in[0] a_6182_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4079 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4080 a_7047_5853# a_6265_5487# a_6963_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4081 _0421_ a_3155_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4082 vccd1 _0243_ a_23671_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4083 vssd1 a_5841_19605# a_5775_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4084 vssd1 net37 a_27167_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4085 vccd1 net31 a_16863_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4086 a_20119_28701# a_19421_28335# a_19862_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4087 vccd1 a_4663_9117# a_4831_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4088 _0027_ a_25235_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4090 a_25198_17973# a_25030_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4091 vccd1 a_12391_7119# a_12559_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4092 a_20004_29257# a_19605_28885# a_19878_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4093 _0289_ a_23804_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X4094 a_23579_13469# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4095 vccd1 cal_lut\[122\] a_10235_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4096 a_20280_7663# a_19881_7663# a_20154_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4097 vssd1 a_14287_17999# net18 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4098 vssd1 _0791_ a_1464_23957# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X4099 a_5946_26819# _0811_ a_5864_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4100 a_17901_21807# _0452_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4101 a_24306_4132# a_24099_4073# a_24482_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4103 vccd1 a_20763_1679# a_20931_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4104 _0690_ a_14747_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4105 a_2287_22325# _0783_ a_2485_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X4106 a_15795_17821# a_14931_17455# a_15538_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4107 dbg_result[1] a_6674_16620# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X4108 cal_lut\[73\] a_26911_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4109 _0854_ a_20308_14441# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X4110 vccd1 a_18371_26525# a_18539_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4111 a_13525_20175# _0447_ a_13275_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4113 vssd1 a_13203_3829# a_13161_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4115 vssd1 a_20471_28853# a_20429_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4118 a_26479_14191# a_26259_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4121 a_18271_24349# a_17489_23983# a_18187_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4122 a_12258_20407# _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4123 vssd1 a_23535_17143# cal_lut\[26\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4124 a_24021_14735# a_23487_14741# a_23926_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4125 a_26443_13103# a_26314_13377# a_26023_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4126 a_26325_18543# _0075_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4128 a_1584_29423# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X4129 a_23281_6409# a_22291_6037# a_23155_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4130 a_24971_5487# a_24835_5461# a_24551_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4131 vssd1 a_6090_27221# a_6019_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4132 a_1753_26133# clknet_0_temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4133 _0773_ _0414_ a_5555_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.36 ps=2.72 w=1 l=0.15
X4134 vccd1 a_12759_17821# a_12927_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4135 _0395_ net75 a_4345_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4136 _0074_ a_24315_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4138 a_6537_19605# clknet_0__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4139 a_15465_17821# a_14931_17455# a_15370_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4140 a_21136_23145# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4141 vssd1 dbg_result[3] a_13942_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4142 vccd1 _0278_ a_12723_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4143 vssd1 a_20322_9269# a_20280_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4144 vccd1 a_19865_13621# _0534_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X4145 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4146 vssd1 a_18151_21271# _0464_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4148 vccd1 a_6947_29691# a_6863_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4149 a_14545_5487# a_14379_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4150 _0469_ a_19287_21835# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X4151 a_26042_10205# a_25769_9839# a_25957_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4152 vccd1 a_10294_13215# a_10221_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4154 _0501_ a_19977_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X4157 a_2023_19319# _0411_ a_2805_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4158 a_10971_2223# cal_lut\[186\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X4159 a_9779_27791# _0386_ _0197_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4160 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4161 vssd1 a_24122_17188# a_24051_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4162 vssd1 cal_lut\[182\] a_9681_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4163 _0647_ a_15378_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X4164 vccd1 _0627_ a_8025_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4165 a_8645_17999# _0520_ a_8491_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4166 a_6087_16733# a_5805_16367# a_5993_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X4167 a_15101_1679# _0184_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4168 _0024_ a_21095_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4169 vssd1 cal_lut\[88\] a_17225_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4170 a_17314_4132# a_17114_3977# a_17463_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4172 _0359_ a_27531_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4173 vccd1 _0352_ a_25603_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4174 a_7841_14013# a_7571_13647# a_7751_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4175 a_24757_18005# a_24591_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4176 a_6541_18005# a_6375_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4177 vssd1 _0242_ a_21739_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4179 a_4885_14741# a_4719_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4180 a_14082_3855# a_13809_3861# a_13997_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4181 vssd1 _0467_ a_9344_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X4182 a_14155_29397# cal_lut\[49\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X4184 a_9821_21583# _0627_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X4185 vssd1 a_4771_20871# _0770_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X4186 vccd1 net24 a_4535_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4187 vccd1 _0711_ a_11896_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4188 a_12212_30199# net9 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X4189 vssd1 _0817_ temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4190 a_10961_14191# _0080_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4191 a_23119_14557# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4192 a_24972_8751# a_24573_8751# a_24846_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4193 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4194 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4195 a_19609_5487# _0113_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4196 a_7715_5461# a_7891_5461# a_7843_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4197 vssd1 cal_lut\[188\] a_5541_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4198 _0066_ a_21739_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4199 a_1937_6549# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4200 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4201 a_19149_25615# _0047_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4202 vccd1 a_7147_3677# a_7315_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4203 vccd1 _0773_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 vssd1 cal_lut\[67\] a_23765_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X4205 vccd1 dbg_result[2] a_14770_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4207 vccd1 net35 a_20727_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4208 a_5555_24233# ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X4209 a_15998_25183# a_15830_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4210 a_3981_14441# _0411_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4211 a_18298_3423# a_18130_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4212 vssd1 _0292_ a_18519_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4213 a_22695_8207# a_21997_8213# a_22438_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4214 vccd1 a_14523_16885# _0442_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4215 a_9957_11177# _0504_ a_9861_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4216 a_15979_12559# a_15115_12565# a_15722_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4217 _0235_ a_21136_23145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4218 a_6645_21263# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X4219 vssd1 a_17727_17999# a_17895_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4220 a_6180_16733# a_5639_16367# a_6087_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X4221 _0232_ a_23391_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4222 vccd1 a_7239_17999# a_7410_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X4223 a_16309_5487# _0498_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X4224 a_9363_19631# _0447_ a_9000_19783# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4225 vssd1 dbg_result[3] a_15115_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X4226 vccd1 a_16737_12533# _0604_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X4227 a_4484_30663# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X4228 a_17999_22923# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4229 vssd1 cal_lut\[14\] a_23124_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X4230 vssd1 a_16731_1653# _0333_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X4231 vccd1 a_9184_20871# _0627_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X4232 vccd1 net25 a_13643_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4233 a_1944_28157# a_1913_28023# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X4234 a_2750_20407# _0421_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X4235 vccd1 net9 a_9135_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X4236 a_16727_4087# a_16823_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4237 a_15649_12559# a_15115_12565# a_15554_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4239 a_8484_20725# a_8297_20765# a_8397_20983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4240 a_12337_3861# a_12171_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4241 temp1.dac_vout_notouch_ net13 a_11152_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X4242 vssd1 net46 a_19255_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4243 a_7277_14191# a_7111_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4246 a_20871_26133# a_21162_26433# a_21113_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4247 a_14618_24501# a_14450_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4248 vssd1 a_9000_19783# _0704_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4249 vssd1 a_16147_3829# a_16105_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4250 vccd1 a_7251_1898# _0186_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4251 vssd1 net23 a_7387_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4252 a_19163_3855# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4254 _0340_ a_19435_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4255 _0432_ a_6375_19095# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4256 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4257 a_24482_3855# a_24235_4233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4258 a_23959_11177# cal_lut\[68\] a_23757_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4259 _0500_ a_16803_22689# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X4262 a_5165_9295# _0138_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4263 vssd1 _0389_ a_2224_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4265 a_17225_25981# a_16955_25615# a_17135_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4266 a_15971_19997# a_15189_19631# a_15887_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4267 a_20338_1679# a_20065_1685# a_20253_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4268 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4269 a_2366_25615# _0746_ a_2209_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4270 vssd1 _0646_ a_15378_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X4271 cal_lut\[42\] a_17159_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4272 a_6565_24527# _0750_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4273 _0680_ _0517_ a_8979_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4274 vssd1 _0363_ a_9547_3073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4275 a_14450_24527# a_14177_24533# a_14365_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4276 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4277 vccd1 a_21334_2335# a_21261_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4278 vssd1 net8 a_10239_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4279 vccd1 a_2564_25045# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X4280 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4281 vccd1 a_7350_2335# a_7277_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4282 vssd1 a_18878_9572# a_18807_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4283 _0705_ _0704_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4285 a_17286_14709# a_17118_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4286 temp1.capload\[15\].cap.Y net55 a_2137_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4287 vssd1 a_19862_28447# a_19820_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4288 _0522_ a_19807_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4289 a_22395_19631# a_22266_19905# a_21975_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4290 a_19709_7485# a_19439_7119# a_19619_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4291 a_2107_19631# _0418_ a_1917_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4292 vccd1 _0739_ _0740_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X4293 vssd1 a_24499_9295# net36 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4294 _0441_ a_17560_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4296 vssd1 clknet_0_temp1.i_precharge_n a_3882_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4297 a_15623_15431# _0531_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4298 vssd1 _0283_ a_21265_7815# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4299 vccd1 a_1857_21365# a_1963_21365# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4300 a_18107_7338# _0293_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4301 vssd1 net44 a_19807_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4302 vccd1 a_15538_17567# a_15465_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4304 a_6541_12015# a_6375_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4305 a_21426_14303# a_21258_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4306 _0499_ a_9678_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X4307 cal_lut\[5\] a_12099_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4310 _0325_ a_4163_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4311 vssd1 _0724_ a_7376_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4312 vssd1 net77 _0398_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4315 vssd1 a_3848_27399# _0830_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4316 a_3850_23759# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4317 vccd1 _0821_ a_4714_23483# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X4318 vccd1 net25 a_9963_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4319 a_8675_10383# _0496_ a_8758_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X4321 vccd1 a_13714_19407# _0495_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4322 a_9678_5487# cal_lut\[146\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X4323 _0272_ a_14283_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4324 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4325 vssd1 _0248_ a_27351_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4326 a_13997_15823# _0035_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4327 vccd1 cal_lut\[168\] a_21879_16055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4329 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4330 vssd1 _0442_ a_15484_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X4331 a_10740_29575# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4332 a_10049_24527# _0715_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4333 a_24683_19087# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4334 a_4843_15307# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4336 vccd1 a_2652_28487# _0832_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X4337 vssd1 ctr\[2\] a_4719_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4338 vccd1 a_11471_14557# a_11639_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4339 vssd1 a_6487_11195# a_6445_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4341 a_10317_7119# _0122_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4342 vccd1 cal_lut\[169\] a_25507_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4343 vccd1 a_7407_12533# a_7323_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4344 a_7994_16479# a_7826_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4346 vssd1 a_2327_22895# _0418_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4347 vssd1 clknet_0_net67 a_3869_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4348 vssd1 net7 a_2576_17271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
X4349 _0741_ a_2742_18082# a_3005_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X4350 vssd1 a_17314_4132# a_17243_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4352 a_17930_24095# a_17762_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4354 a_2739_30333# _0800_ a_2376_30199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4355 a_23547_26921# net47 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4356 a_10689_9839# _0450_ a_10607_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4357 _0231_ a_22747_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4358 a_17661_4233# a_17107_4073# a_17314_4132# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4359 a_25873_6397# a_25603_6031# a_25783_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4360 vccd1 a_27923_9019# a_27839_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4361 a_9586_19407# _0591_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X4363 vssd1 cal_lut\[106\] a_16168_9411# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4364 a_12391_7119# a_11527_7125# a_12134_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4365 vssd1 a_5503_27399# ctr\[7\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4366 a_9403_32463# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X4367 vccd1 a_11759_4564# _0129_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4368 vccd1 a_5170_10660# a_5099_10761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4369 a_24835_5461# net33 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4370 vssd1 a_15170_10357# a_15128_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4371 a_3991_26409# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X4372 vccd1 a_3851_25045# _0803_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X4374 a_2939_23047# _0410_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4375 a_13514_21237# a_13346_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4377 a_16382_11293# a_15943_10927# a_16297_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4378 a_4771_20871# net21 a_5099_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4381 vccd1 a_9983_14459# a_9899_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4382 vssd1 _0299_ a_7005_4551# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4383 a_15281_3861# a_15115_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4384 vccd1 a_18383_5175# _0541_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4385 a_14875_24527# a_14177_24533# a_14618_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4386 vssd1 net27 a_6375_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4387 vccd1 _0411_ _0428_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4388 vccd1 _0257_ a_10699_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4389 vccd1 a_5508_24501# _0796_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X4390 a_26961_18543# a_25971_18543# a_26835_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4392 _0414_ a_2419_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4393 _0561_ a_19426_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X4394 vssd1 a_12815_20719# _0446_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4395 cal_lut\[114\] a_20287_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4396 _0014_ a_23671_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4397 a_22971_13469# a_22273_13103# a_22714_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4398 a_9967_24847# _0718_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X4399 a_2931_17455# _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4400 a_13346_21263# a_13073_21269# a_13261_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4401 vssd1 a_7410_17973# dbg_result[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X4403 a_21810_16733# a_21537_16367# a_21725_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4404 a_13714_4943# a_13275_4949# a_13629_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4405 a_11522_8751# a_11207_8903# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4406 _0278_ a_12259_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4407 a_10570_7093# a_10402_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4409 _0080_ a_10699_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4410 a_9022_8207# a_8583_8213# a_8937_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4411 vssd1 a_23903_18695# _0642_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4412 vccd1 a_21371_17455# net42 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4413 vssd1 net11 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4414 a_23097_13103# a_22107_13103# a_22971_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4415 a_14710_1247# a_14542_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
R13 vssd1 net54 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4416 vccd1 cal_lut\[102\] a_15972_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4418 a_9037_28585# _0406_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.28 ps=2.56 w=1 l=0.15
X4419 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4421 vccd1 cal_lut\[8\] a_12995_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4422 a_2931_22325# _0773_ a_3149_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X4423 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4424 a_12737_18543# net15 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4425 a_6820_24527# _0751_ a_6565_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4426 a_20433_27797# a_20267_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4427 cal_lut\[71\] a_28015_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4429 _0686_ a_22291_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4432 a_19789_28701# a_19255_28335# a_19694_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4433 vccd1 a_9831_24501# _0727_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4434 a_23811_15431# _0460_ a_24045_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4435 a_24835_13077# net36 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4437 a_1477_10901# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4438 a_17717_19453# _0474_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4440 a_21261_2589# a_20727_2223# a_21166_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4441 vssd1 _0291_ a_19807_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4443 a_2043_31055# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X4444 vssd1 _0817_ temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4445 vssd1 _0269_ a_17875_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4446 vssd1 a_2511_21263# io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4448 a_15285_28879# _0044_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4449 _0811_ a_5179_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X4452 cal_lut\[37\] a_8143_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4453 vssd1 a_15538_28853# a_15496_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4454 a_24731_6740# _0348_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4455 vccd1 _0443_ a_18979_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4456 a_19789_4765# a_19255_4399# a_19694_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4457 cal_lut\[110\] a_23875_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4460 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4461 a_22185_23439# _0060_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4462 vccd1 net47 a_24407_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4463 a_10827_7119# a_10129_7125# a_10570_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4464 a_2839_27221# net70 a_3048_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X4465 vccd1 _0452_ a_15851_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4466 vssd1 a_4676_25223# _0828_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X4469 vssd1 a_2747_18517# net22 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4470 _0143_ a_6559_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4471 a_8758_10703# cal_lut\[37\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X4472 vssd1 a_23875_7931# a_23833_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4473 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4474 a_16949_1135# a_16679_1501# a_16859_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4475 _0263_ a_21872_24643# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X4476 vccd1 cal_lut\[34\] a_17628_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4477 a_16820_17705# _0611_ a_16718_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X4479 a_5278_12533# a_5404_12797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.186 ps=1.26 w=0.65 l=0.25
X4480 vccd1 cal_lut\[71\] a_26830_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4481 net41 a_7072_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4484 a_17088_12265# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4485 vccd1 _0266_ a_14103_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4486 _0671_ a_11715_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X4487 _0558_ a_18979_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4488 a_14705_17620# _0555_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4489 _0411_ a_1651_14165# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4490 vssd1 a_4811_30511# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4491 vccd1 a_1551_19605# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4492 vssd1 a_3615_17999# _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4494 _0152_ a_22659_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4495 a_21541_6575# _0157_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4496 vssd1 a_27035_8181# _0351_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X4497 vccd1 a_8419_9019# a_8335_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4498 vccd1 _0446_ a_3885_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X4499 vccd1 a_10083_24135# _0713_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4500 vssd1 cal_lut\[3\] a_9313_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4501 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4502 a_10041_13103# _0020_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4503 _0489_ a_15391_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4504 vssd1 _0763_ a_1959_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X4506 vccd1 a_7975_18909# a_8146_18796# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X4507 vssd1 cal_lut\[73\] a_23305_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X4508 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4509 _0847_ a_12443_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4511 a_2121_21623# _0414_ a_2049_21623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4512 vssd1 dbg_result[2] a_15662_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.107 ps=0.98 w=0.65 l=0.15
X4513 vssd1 a_20963_15797# _0222_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4515 a_13346_21263# a_12907_21269# a_13261_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4516 a_9096_27221# _0816_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4517 a_1761_14735# _0199_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4518 vssd1 a_21759_25339# a_21717_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4519 vssd1 a_26330_14165# a_26259_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4521 vccd1 a_16355_29397# a_16179_29397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X4522 a_2497_14191# _0202_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4523 vssd1 a_10699_4399# _0850_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4524 vssd1 a_1464_23957# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4527 _0364_ a_16859_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4528 a_27503_15253# net37 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4529 _0478_ a_22843_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4530 vccd1 cal_lut\[13\] a_21735_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4531 a_9043_10089# _0698_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4532 vccd1 a_12815_20719# _0446_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4533 _0430_ _0427_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4534 vssd1 a_5291_5755# a_5249_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4536 a_20713_19631# _0059_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4537 a_20947_3677# a_20249_3311# a_20690_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4538 a_15262_29535# a_15094_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4539 _0453_ dbg_result[4] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4540 cal_lut\[72\] a_28199_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4541 a_26651_6941# a_25787_6575# a_26394_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4542 a_4333_27797# a_4167_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4544 vssd1 _0641_ a_22625_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X4545 a_5883_27221# clknet_1_1__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4548 a_4606_27791# a_4333_27797# a_4521_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
R14 temp1.capload\[4\].cap_59.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4549 vccd1 cal_lut\[106\] a_16250_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4550 a_12885_17455# a_11895_17455# a_12759_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4551 a_23823_20393# net43 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4552 cal_lut\[13\] a_21851_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4553 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4554 _0125_ a_14195_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4555 vccd1 a_26307_13077# a_26314_13377# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4556 a_17498_29397# a_17298_29697# a_17647_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4557 vssd1 _0741_ a_4995_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X4559 vccd1 a_14250_3829# a_14177_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4560 vssd1 a_7716_25589# _0750_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X4561 _0859_ a_17088_12265# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4562 a_12617_13103# _0021_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4563 a_1917_19881# net22 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4564 vssd1 _0278_ a_12723_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4565 a_20069_9295# _0107_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4567 _0664_ a_10596_17705# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X4568 a_8263_15444# _0255_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4571 a_22677_27613# a_22339_27399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4572 vssd1 a_9385_4373# _0503_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X4574 vssd1 cal_lut\[156\] a_19525_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4575 _0657_ a_21003_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4576 cal_lut\[188\] a_7775_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4577 vssd1 _0406_ a_8845_28023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4578 cal_lut\[25\] a_22403_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4580 a_1551_19605# _0761_ a_1917_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.585 ps=2.17 w=1 l=0.15
X4581 a_1464_23957# _0414_ a_2121_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0747 ps=0.88 w=0.65 l=0.15
X4582 a_6637_5175# _0299_ a_6800_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4583 a_23477_8751# _0450_ a_23395_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4584 vssd1 _0519_ a_11895_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
X4586 vssd1 net31 a_20727_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4587 a_22925_4399# _0451_ a_22843_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4588 a_9493_8751# _0476_ a_9411_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4589 vssd1 _0335_ a_21463_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4590 vssd1 _0705_ a_10761_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4591 _0517_ _0516_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4592 a_13840_5321# a_13441_4949# a_13714_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4593 a_13691_28500# _0224_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4594 a_14321_19881# _0447_ a_14237_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4595 a_9313_16367# a_9043_16733# a_9223_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4596 a_9148_8585# a_8749_8213# a_9022_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4597 a_2489_8181# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4599 vssd1 a_18171_6843# a_18129_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4600 a_8246_8323# _0299_ a_8164_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4602 a_1953_7439# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4603 _0419_ ctr\[2\] a_2782_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X4604 vssd1 a_9647_14709# _0256_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X4605 a_23610_10089# _0658_ a_23361_9985# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4606 a_9678_29156# a_9478_29001# a_9827_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4607 a_2330_24887# _0412_ a_2249_24887# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X4610 vccd1 a_2092_31287# a_2043_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X4612 vssd1 a_7439_4373# _0299_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4614 a_9358_3855# cal_lut\[181\] a_9201_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4616 _0011_ a_18151_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4617 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4811_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X4618 a_17433_15823# a_17095_16055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4619 a_21913_9661# _0450_ a_21831_9408# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4620 a_3851_15253# _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.14 ps=1.08 w=0.65 l=0.15
X4621 vssd1 a_15703_2767# a_15871_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4622 a_15094_27791# a_14655_27797# a_15009_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4623 vccd1 _0836_ a_5271_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4624 a_27774_12533# a_27606_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4626 vccd1 a_16423_25339# a_16339_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4627 vssd1 _0785_ a_7716_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4628 a_5709_15113# a_4719_14741# a_5583_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4629 a_9991_6031# a_9209_6037# a_9907_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4631 vccd1 _0424_ a_3075_24305# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4632 a_26743_16733# a_26045_16367# a_26486_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4633 temp1.capload\[14\].cap.Y clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4634 vssd1 _0755_ a_6548_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4635 a_24945_17999# _0074_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4636 a_20556_17289# a_20157_16917# a_20430_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4637 _0128_ a_10331_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4638 a_8397_24527# dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4639 a_24653_4233# a_24106_3977# a_24306_4132# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4641 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4642 a_4381_21807# _0759_ a_4283_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X4643 a_23841_14735# _0067_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4645 a_22714_13215# a_22546_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4646 a_5722_28111# _0811_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X4647 a_3057_19407# _0418_ a_2973_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4649 a_2023_19319# _0745_ a_2447_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4650 vssd1 net79 _0402_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4651 vccd1 a_20506_1653# a_20433_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4652 a_22362_14735# a_21923_14741# a_22277_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4653 a_6706_5599# a_6538_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4654 vssd1 _0708_ a_12097_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4655 vssd1 a_23351_21959# _0638_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X4656 _0630_ a_9933_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.91 w=0.65 l=0.15
X4657 a_5165_13103# _0204_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4658 a_8675_10383# cal_lut\[187\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X4659 vssd1 a_12310_10615# _0660_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X4660 vssd1 a_11302_16519# _0629_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4661 vccd1 a_9823_15041# a_9647_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X4662 a_17007_29397# a_17291_29397# a_17226_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4663 a_8617_22351# _0775_ a_8533_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4664 vccd1 cal_lut\[176\] a_22790_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X4666 a_28115_15823# a_27333_15829# a_28031_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4667 a_25823_23439# a_24959_23445# a_25566_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4668 vccd1 _0462_ a_22843_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4669 a_6706_5599# a_6538_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4670 _0648_ a_22383_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4671 vccd1 a_26267_17723# a_26183_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4672 a_6920_15113# a_6541_14741# a_6823_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X4673 _0661_ _0515_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4674 cal_lut\[114\] a_20287_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4675 a_8749_8213# a_8583_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4677 vssd1 _0795_ a_5508_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4678 _0297_ a_23344_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X4679 vssd1 cal_lut\[85\] a_21872_24643# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4680 _0085_ a_22291_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4681 _0193_ _0382_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4682 vccd1 a_6244_25045# _0807_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X4683 vccd1 _0485_ a_20359_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4684 vccd1 cal_lut\[100\] a_14776_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4685 vssd1 a_4313_17429# _0790_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4687 vccd1 cal_lut\[167\] a_27347_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4688 a_14177_24533# a_14011_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4689 a_10247_21583# _0557_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4690 a_7749_28335# _0815_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4691 a_19862_24501# a_19694_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4692 a_17973_21807# cal_lut\[84\] a_17901_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4693 a_25493_23439# a_24959_23445# a_25398_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4694 _0591_ _0589_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4695 _0616_ a_16127_5056# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4696 a_10221_11471# a_9687_11477# a_10126_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4698 a_16158_7913# _0545_ a_15909_7809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4699 vssd1 net40 a_12539_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4700 a_5449_8573# a_5179_8207# a_5359_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4701 cal_lut\[62\] a_25439_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4702 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4703 a_15071_13268# _0852_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4705 a_25014_7093# a_24846_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4706 _0574_ a_13091_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X4707 a_14611_11079# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4708 vssd1 a_10827_1679# a_10995_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4709 a_22185_8207# _0108_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4710 vssd1 a_12943_1679# a_13111_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4711 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4712 vccd1 a_22619_15253# net37 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4713 a_22806_3829# a_22638_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4715 vccd1 _0259_ a_17323_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4716 _0291_ a_19619_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4717 a_9224_6575# _0476_ a_9034_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X4718 a_14139_4943# a_13441_4949# a_13882_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4719 a_10262_24847# _0726_ a_9967_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X4720 a_2563_23957# _0823_ a_2790_24305# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X4721 _0455_ a_12950_16988# a_13309_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.52 pd=3.04 as=0.135 ps=1.27 w=1 l=0.15
X4722 vssd1 cal_lut\[66\] a_21228_15529# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4723 vssd1 net40 a_14655_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4724 a_23903_18695# net18 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4725 a_6779_9117# a_6081_8751# a_6522_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4726 a_12097_23983# _0706_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4727 vccd1 a_22259_19605# a_22266_19905# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4728 a_11579_3829# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X4729 a_24455_5639# a_24551_5461# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4730 vssd1 _0261_ a_18979_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4732 a_15715_30186# _0218_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4733 a_7255_20871# ctr\[10\] a_7381_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4734 vccd1 a_22903_2985# a_22910_2889# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4735 a_24306_4132# a_24106_3977# a_24455_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4736 a_18475_5639# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4737 _0097_ a_12815_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4738 net81 a_15023_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4739 vssd1 _0514_ _0515_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4740 cal_lut\[52\] a_18815_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4741 vccd1 _0782_ a_2931_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4742 a_15299_25615# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4743 a_17739_21959# _0531_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4744 a_9209_6037# a_9043_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4745 vssd1 a_12743_26677# a_12701_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4747 _0535_ a_19255_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X4748 vccd1 a_2009_30676# io_out[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4750 a_4069_25071# net21 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4751 _0083_ a_18979_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4752 a_9452_32375# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4754 vccd1 a_6779_29789# a_6947_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4756 _0393_ _0808_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4758 vssd1 cal_lut\[116\] a_23344_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4759 a_19793_21959# _0222_ a_19956_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4760 a_9113_15113# a_8123_14741# a_8987_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4761 vssd1 a_5971_15253# a_5713_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X4762 a_12425_3311# a_11435_3311# a_12299_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4763 a_12079_5737# cal_lut\[129\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X4764 a_14651_6575# cal_lut\[125\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X4765 io_out[3] a_2287_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4766 a_25271_7119# a_24573_7125# a_25014_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4767 vccd1 a_10719_11445# a_10635_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4768 vccd1 net44 a_20359_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4769 vssd1 _0776_ a_5813_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X4770 vccd1 a_5779_8426# _0141_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4771 a_27606_12559# a_27167_12565# a_27521_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4773 a_21971_13879# _0474_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4774 _0532_ a_19807_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4775 a_22438_27765# a_22270_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4776 vccd1 net48 a_13551_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4777 a_11950_18319# _0574_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X4779 vccd1 a_25375_12167# cal_lut\[176\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4780 a_11243_30761# net13 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X4781 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4782 vccd1 _0237_ a_16955_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4783 vccd1 _0850_ a_25143_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4784 _0287_ a_17871_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X4786 vssd1 _0717_ a_10505_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4787 vccd1 a_1458_30199# a_1407_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4788 _0539_ _0525_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4789 a_20046_28853# a_19878_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4790 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4791 vccd1 _0517_ a_8769_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.117 ps=1.24 w=1 l=0.15
X4792 a_20407_16519# _0459_ a_20641_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4794 vccd1 net29 a_12263_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4795 a_4885_6037# a_4719_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4796 a_17302_2589# a_17029_2223# a_17217_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4797 a_15378_18543# _0438_ a_15289_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0619 ps=0.715 w=0.42 l=0.15
X4798 _0382_ clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4799 a_24761_8751# _0164_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4800 vccd1 _0201_ a_3953_10761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4801 a_23719_4087# a_23815_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4802 vssd1 a_8251_9117# a_8419_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4803 a_22270_27791# a_21997_27797# a_22185_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4804 a_7491_19087# _0439_ a_6979_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X4805 a_6955_23671# _0705_ a_7101_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4806 vccd1 _0453_ a_19439_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4807 a_20433_1679# a_19899_1685# a_20338_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4808 vccd1 a_3339_9295# net30 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4809 vssd1 net8 a_11243_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X4810 a_20572_6031# _0583_ a_20470_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4811 _0767_ _0432_ a_5915_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4813 a_4977_29789# a_4443_29423# a_4882_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4814 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4815 a_10975_20719# _0678_ a_10975_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4816 _0473_ a_22875_17249# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X4817 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4818 vssd1 a_21879_19783# cal_lut\[59\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4820 a_25363_15823# a_24665_15829# a_25106_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4821 a_6636_25321# _0751_ a_6381_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4822 _0162_ a_26799_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4823 a_19667_18517# dbg_result[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4824 a_14821_27797# a_14655_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4825 vccd1 a_5507_22325# _0789_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4826 vccd1 _0290_ a_14471_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X4827 a_15255_28500# _0270_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4828 a_8556_20725# dec1.i_ones a_8484_20725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4829 a_23063_25437# a_22365_25071# a_22806_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4831 vccd1 net53 temp1.capload\[13\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4832 a_27774_11445# a_27606_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4833 temp1.capload\[5\].cap.Y net60 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4834 a_20579_9295# a_19715_9301# a_20322_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4835 a_6541_12015# a_6375_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4836 a_20522_21263# a_20083_21269# a_20437_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4837 vssd1 a_10562_19319# _0666_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X4838 _0719_ _0718_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4839 a_5416_23413# _0737_ a_5639_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X4840 a_13146_23007# a_12978_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4841 a_17109_20719# cal_lut\[42\] a_17037_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4842 a_6265_5487# a_6099_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4843 vssd1 _0784_ a_3933_28918# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X4844 vccd1 _0267_ a_17231_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4845 a_7631_17171# dbg_result[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4848 vccd1 a_18291_9527# cal_lut\[106\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4851 _0195_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4852 vccd1 cal_lut\[85\] a_21954_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4853 vccd1 a_25566_23413# a_25493_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4854 vccd1 a_1959_21807# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4855 _0472_ _0447_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4856 a_27035_8181# cal_lut\[166\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X4857 _0102_ a_18335_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4858 vccd1 a_10294_11445# a_10221_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4859 vccd1 _0441_ a_12539_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4860 vssd1 _0341_ a_22887_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4861 a_6729_12015# _0190_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4862 vccd1 _0748_ a_8485_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4863 vssd1 _0447_ _0382_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4864 a_25941_5321# a_25394_5065# a_25594_5220# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4865 vccd1 cal_lut\[55\] a_21919_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4866 a_24101_27081# a_23554_26825# a_23754_26980# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4867 vccd1 a_15469_20407# _0878_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X4868 vccd1 a_21971_13879# _0533_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4869 a_16983_23047# cal_lut\[88\] a_17129_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4870 a_14729_21269# a_14563_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4871 a_10241_19203# _0629_ a_10145_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4872 a_20775_18231# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4873 a_21257_28169# a_20267_27797# a_21131_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4875 a_28149_14025# a_27602_13769# a_27802_13924# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4877 a_26693_21807# _0063_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4878 a_21923_21376# cal_lut\[87\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4880 a_26486_16479# a_26318_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4881 a_25198_17973# a_25030_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4882 a_15369_5487# a_14379_5487# a_15243_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4883 a_9963_9001# _0493_ a_10046_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X4884 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_1584_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X4885 _0332_ a_13639_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4886 vssd1 a_7791_27613# a_7959_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4887 cal_lut\[123\] a_10995_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4888 vssd1 a_24473_9813# _0511_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X4890 vccd1 _0631_ a_11869_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X4891 a_21349_19631# a_20359_19631# a_21223_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4892 cal_lut\[122\] a_9615_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4893 net69 clknet_1_1__leaf_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4894 vssd1 a_10851_11079# _0496_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X4895 io_out[5] a_2564_25045# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4896 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4897 a_5135_25398# _0827_ a_4676_25223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X4898 a_10924_31751# net65 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4899 vssd1 _0495_ a_10853_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4900 vssd1 a_5326_6005# a_5284_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4901 a_6982_12127# a_6814_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4902 a_18187_24349# a_17323_23983# a_17930_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4903 _0116_ a_23671_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4904 a_23125_20719# cal_lut\[57\] a_23053_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4905 vssd1 a_24306_4132# a_24235_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4906 vssd1 a_10943_23671# _0717_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X4907 vssd1 _0437_ a_8111_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X4908 vccd1 _0521_ _0764_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4909 a_25030_17999# a_24757_18005# a_24945_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4910 vssd1 a_14151_5652# _0118_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4911 a_15005_7119# a_14471_7125# a_14910_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4913 a_24653_4233# a_24099_4073# a_24306_4132# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4914 a_9375_29397# ctr\[11\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4915 a_20635_6941# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4916 vccd1 _0442_ a_18698_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4918 _0464_ a_18151_21271# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4919 vccd1 _0465_ a_21923_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X4920 cal_lut\[77\] a_17895_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4921 a_4128_20149# net21 a_4520_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X4922 a_24863_19087# a_24683_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4923 a_3091_14557# a_2309_14191# a_3007_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4924 a_12212_30199# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4926 vssd1 _0380_ a_7102_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4927 a_10247_21583# _0627_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X4928 vssd1 a_14655_18115# _0491_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X4930 a_14131_13879# cal_lut\[22\] a_14277_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4931 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd _0746_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4932 vccd1 a_11292_30663# a_11243_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X4933 a_12701_27081# a_11711_26709# a_12575_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4935 vccd1 _0837_ a_1867_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4936 a_19807_22895# cal_lut\[90\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4937 _0611_ a_16035_18112# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4938 a_15569_3311# a_15299_3677# a_15479_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X4939 vssd1 a_25271_25437# a_25439_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4940 a_5460_17999# _0384_ a_5825_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4941 a_23745_19087# a_23211_19093# a_23650_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4942 vccd1 a_18555_3677# a_18723_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4943 a_12621_6397# _0441_ a_12539_6144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4944 vccd1 net41 a_7939_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4946 vccd1 clknet_1_0__leaf_io_in[0] a_6375_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4947 vssd1 net42 a_24499_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4948 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4950 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4951 vssd1 _0502_ a_18416_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X4952 a_22270_27791# a_21831_27797# a_22185_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4953 a_12263_20495# a_12258_20407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=2.52 w=1 l=0.15
X4954 a_24377_20553# a_23830_20297# a_24030_20452# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4955 a_4921_10383# a_4583_10615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4956 vccd1 _0282_ a_20175_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4957 a_12545_19087# _0519_ _0556_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X4958 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4960 a_20154_8029# a_19881_7663# a_20069_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4961 _0524_ a_19071_11584# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4962 a_1972_12937# a_1573_12565# a_1846_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4963 a_7553_25071# _0728_ a_7457_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X4964 a_21029_12043# _0505_ a_20943_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4965 a_3981_14441# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X4966 _0397_ net72 a_3891_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4967 _0330_ a_12223_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4968 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd _0773_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4969 vccd1 a_22891_20871# _0636_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4970 a_25674_17821# a_25235_17455# a_25589_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4971 a_19409_7663# cal_lut\[144\] a_19337_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4972 vccd1 _0718_ _0719_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4973 a_7975_14557# a_7277_14191# a_7718_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4974 vccd1 a_24030_20452# a_23959_20553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4975 a_14158_26677# a_13990_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4976 vssd1 _0706_ _0729_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4977 a_22633_11445# _0451_ a_22886_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X4978 vccd1 a_13863_12559# a_14031_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4979 vssd1 net9 a_9135_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4981 vssd1 a_4678_26311# _0800_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0878 ps=0.92 w=0.65 l=0.15
X4982 vssd1 _0390_ a_6546_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X4983 a_25415_22351# a_25235_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4984 a_20985_14191# a_20819_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4986 a_18015_5639# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4988 a_13104_25071# a_12705_25071# a_12978_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4990 vssd1 a_13863_12559# a_14031_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4991 vccd1 net41 a_14563_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4992 a_4698_5853# a_4425_5487# a_4613_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4993 a_11030_27383# a_10871_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4994 cal_lut\[82\] a_13571_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4995 vssd1 a_8263_15444# _0078_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4996 a_26506_14557# a_26259_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4997 a_16640_4373# net34 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
R15 net66 vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4998 a_12042_3423# a_11874_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5000 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5001 a_15535_24501# cal_lut\[94\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X5002 a_5077_24233# _0429_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5003 vccd1 a_25531_15797# a_25447_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5004 a_17789_19453# cal_lut\[76\] a_17717_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5005 a_17762_1679# a_17489_1685# a_17677_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5006 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5007 vccd1 a_15427_21263# a_15595_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5008 vccd1 a_17919_3073# a_17743_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X5009 vccd1 cal_lut\[133\] a_9358_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X5010 vccd1 net33 a_25787_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5011 vssd1 a_23351_8439# _0640_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5012 a_9275_28023# ctr\[12\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5013 cal_lut\[148\] a_13019_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5014 a_2139_12265# _0390_ a_1921_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5015 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5016 vssd1 a_17187_18708# _0076_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5017 a_22051_6941# a_21353_6575# a_21794_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5018 cal_lut\[43\] a_17159_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5019 vssd1 a_15427_21263# a_15595_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5020 a_13074_11293# a_12827_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5021 vssd1 a_2563_23957# _0824_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5022 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5024 a_21831_9408# cal_lut\[105\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5025 a_9459_19958# _0703_ a_9000_19783# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5026 a_15887_19997# a_15023_19631# a_15630_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5027 vssd1 a_14703_21972# _0040_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5028 _0167_ a_27259_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5029 vssd1 _0838_ a_12355_21271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5030 vccd1 a_16991_22173# a_17159_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5032 _0784_ _0414_ a_3991_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.36 ps=2.72 w=1 l=0.15
X5033 a_18611_22895# cal_lut\[83\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5034 a_27503_15253# net37 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5035 a_17187_18708# _0253_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5036 a_24846_9117# a_24573_8751# a_24761_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5037 a_12705_14557# a_12171_14191# a_12610_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5038 vccd1 a_13035_3855# a_13203_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5039 a_12851_2589# a_12153_2223# a_12594_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5040 vccd1 net45 a_17323_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5041 a_22711_6549# cal_lut\[158\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X5043 vssd1 net45 a_17323_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5044 vccd1 a_21879_16055# _0551_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
R16 temp1.capload\[8\].cap_63.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5046 a_4584_23671# a_4714_23483# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X5047 a_15557_19997# a_15023_19631# a_15462_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5048 a_6814_12559# a_6375_12565# a_6729_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5049 a_1917_19631# _0418_ a_2107_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5050 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5051 vssd1 cal_lut\[11\] a_17732_14441# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5052 a_22270_8207# a_21831_8213# a_22185_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5053 vssd1 _0578_ a_17094_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5054 vccd1 net28 a_8123_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5057 a_5883_27221# clknet_1_1__leaf_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5058 vccd1 a_9372_24135# _0724_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5059 a_20245_4399# a_19255_4399# a_20119_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5060 vccd1 _0722_ a_7291_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5061 vssd1 _0498_ a_16484_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X5064 a_24099_12777# net36 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5065 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5066 vssd1 a_19333_24135# _0261_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X5069 vccd1 _0514_ a_15943_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5070 vccd1 a_4593_8439# a_4406_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5071 a_10401_9615# cal_lut\[97\] a_9963_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5072 vccd1 net28 a_6375_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5073 vssd1 a_20779_15253# _0851_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5074 vssd1 a_3695_23671# _0791_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5075 a_8803_15823# a_7939_15829# a_8546_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5076 a_11199_17607# _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.157 ps=1.17 w=0.42 l=0.15
X5077 a_14208_16201# a_13809_15829# a_14082_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5078 vssd1 _0676_ a_11508_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5079 a_26479_16042# _0249_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5080 a_6745_27791# _0826_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5081 vssd1 a_21235_9514# _0104_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5082 vssd1 clknet_0_net67 a_3869_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5084 a_2931_17455# _0422_ a_2489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5085 a_4140_32143# a_3891_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X5086 vccd1 _0452_ a_18611_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5087 vccd1 a_18519_21263# _0454_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5088 _0759_ a_3995_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X5089 net3 a_1407_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5090 vssd1 a_21975_2741# _0337_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5091 vssd1 cal_lut\[118\] a_13040_6147# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5092 cal_lut\[108\] a_20747_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5095 a_20671_22351# a_19807_22357# a_20414_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5096 vssd1 a_5751_14709# a_5709_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5097 a_23351_7338# _0289_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5098 cal_lut\[73\] a_26911_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5099 a_11046_14557# a_10607_14191# a_10961_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5100 vssd1 a_15611_13647# a_15779_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5101 vssd1 net11 a_9403_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X5102 vccd1 a_23818_19061# a_23745_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5103 a_15036_7497# a_14637_7125# a_14910_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5104 vssd1 a_6927_16911# net48 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5105 a_4726_24893# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X5106 a_8473_15823# a_7939_15829# a_8378_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5108 vccd1 _0670_ a_9167_21601# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5110 a_22240_4649# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5111 _0827_ _0435_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X5112 _0838_ a_2235_9303# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5113 vssd1 _0691_ a_21878_17143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X5114 vssd1 a_14733_15431# _0879_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X5116 vssd1 cal_lut\[2\] a_9135_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5117 a_18597_13077# net80 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5119 vssd1 _0087_ a_21709_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5120 a_6055_10602# _0375_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5121 vssd1 cal_lut\[57\] a_23481_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5122 a_22596_10383# _0456_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5123 a_5143_11445# ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5124 vccd1 _0338_ a_19439_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5126 a_20341_22351# a_19807_22357# a_20246_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5127 cal_lut\[138\] a_5751_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5128 a_22561_2223# a_22291_2589# a_22471_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5129 vssd1 a_9563_28487# _0406_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5130 a_14365_24527# _0093_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5131 a_9223_16733# a_9043_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5132 a_13169_9295# _0099_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5133 a_12895_18543# net16 _0557_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X5134 a_9577_6031# a_9043_6037# a_9482_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5136 vccd1 a_22719_27221# a_22726_27521# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5137 vccd1 a_19402_25589# a_19329_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5138 vccd1 a_15135_7931# a_15051_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5139 a_6729_12559# _0018_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5140 vccd1 _0871_ a_18611_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5141 _0746_ ctr\[3\] a_3169_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X5142 _0869_ a_23483_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X5143 a_9411_1679# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5144 vssd1 cal_lut\[138\] a_5404_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5145 a_21997_27797# a_21831_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5148 a_17349_13103# _0474_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X5149 vccd1 a_9558_1247# a_9485_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5150 cal_lut\[152\] a_22863_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5151 _0857_ a_23759_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X5152 vssd1 _0664_ a_11884_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5153 a_17118_14735# a_16679_14741# a_17033_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5154 vccd1 ctr\[1\] _0389_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5155 vccd1 _0704_ a_8971_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X5157 vccd1 a_17470_2335# a_17397_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5158 a_12162_5737# cal_lut\[183\] a_12079_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5159 a_9531_8207# a_8749_8213# a_9447_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5160 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5161 vssd1 _0779_ a_6929_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X5162 a_22695_1679# a_21831_1685# a_22438_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5163 a_16025_7485# _0514_ a_15943_7232# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5164 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5165 a_15727_21959# _0483_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5166 vssd1 _0421_ a_2931_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5167 vssd1 a_4951_7338# _0142_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5168 vssd1 _0506_ a_20900_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X5170 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5171 a_20245_24905# a_19255_24533# a_20119_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5172 a_26330_14165# a_26123_14165# a_26506_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5173 a_21173_14191# _0012_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5174 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5176 vssd1 a_25287_12533# _0361_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5177 a_6831_6575# cal_lut\[144\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X5179 net42 a_21371_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5180 vccd1 _0850_ a_24407_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5181 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5182 a_14637_7125# a_14471_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5183 a_3399_10601# clknet_1_0__leaf_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5184 vccd1 clknet_1_1__leaf_io_in[0] a_5915_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5185 a_4345_13353# _0809_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.28 ps=2.56 w=1 l=0.15
X5186 vccd1 a_26635_10107# a_26551_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5187 _0381_ _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5188 vccd1 cal_lut\[18\] a_20848_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5189 a_9761_15829# a_9595_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5191 a_8335_29789# a_7553_29423# a_8251_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5192 vccd1 net46 a_20267_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5193 vccd1 _0177_ a_17661_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5194 a_4180_12937# a_3781_12565# a_4054_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5196 a_9737_28363# _0815_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X5197 _0059_ a_20359_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5198 vssd1 _0276_ a_12815_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5199 a_10041_11471# _0038_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5201 a_26259_14191# a_26123_14165# a_25839_14165# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5202 a_27595_13865# net37 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5203 a_27071_11293# a_26891_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5204 a_12898_10901# a_12691_10901# a_13074_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5205 vssd1 a_24835_13077# a_24842_13377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5206 a_7557_28640# _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5207 a_11581_21781# _0673_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X5208 vssd1 _0724_ _0734_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5210 vssd1 a_22438_1653# a_22396_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5211 a_6737_16189# a_6467_15823# a_6647_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5212 vccd1 _0450_ a_21003_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5213 vssd1 net23 a_7663_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5214 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5215 vccd1 _0438_ a_4897_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5216 vccd1 a_20747_9269# a_20663_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5217 vccd1 a_21131_27791# a_21299_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5219 a_17243_4233# a_17114_3977# a_16823_4087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5220 vssd1 _0372_ a_17231_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5221 a_9033_13353# _0503_ a_8951_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5222 a_8565_28879# a_8329_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X5223 _0419_ _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5225 a_15611_13647# a_14747_13653# a_15354_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5226 vccd1 a_5675_9295# a_5843_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5227 vccd1 cal_lut\[172\] a_27071_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5228 vccd1 a_12778_14303# a_12705_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5229 vssd1 net27 a_6743_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5230 vssd1 a_2839_27221# _0831_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5232 a_5503_27399# a_5599_27221# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5233 vssd1 _0243_ a_23671_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5234 a_24105_10357# _0476_ a_24358_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X5235 vssd1 a_6062_11039# a_6020_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5236 vccd1 a_13969_18218# net16 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5237 a_4531_17705# _0427_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5238 a_7921_16733# a_7387_16367# a_7826_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5239 a_9929_10357# _0515_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X5240 a_22465_18793# _0647_ a_22383_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5241 vssd1 _0246_ a_26417_18231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5242 _0411_ a_1651_14165# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5243 vssd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5245 vccd1 a_7256_21237# _0778_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X5246 vssd1 _0443_ a_19133_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5247 a_15830_25437# a_15557_25071# a_15745_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5248 _0805_ a_3525_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X5249 net22 a_2747_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5250 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5251 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5252 net13 a_11120_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5253 vssd1 _0836_ a_11605_16055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5254 a_15281_13647# a_14747_13653# a_15186_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5255 _0447_ a_14103_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5256 vccd1 clknet_1_0__leaf_io_in[0] a_5639_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5257 a_22414_10383# _0634_ a_22165_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5258 vssd1 _0482_ a_17117_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5260 a_16734_21919# a_16566_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5261 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd _0784_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5262 a_5639_27791# ctr\[7\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X5263 a_22396_8585# a_21997_8213# a_22270_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5264 a_16382_11293# a_16109_10927# a_16297_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5265 a_22054_12559# _0452_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X5266 a_6729_7119# _0143_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5267 a_13441_4949# a_13275_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5268 a_14441_8573# cal_lut\[112\] a_14369_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5269 vccd1 _0438_ a_12263_20495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.22 ps=1.44 w=1 l=0.15
X5270 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4140_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X5272 a_1951_29199# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X5274 _0102_ a_18335_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5276 a_12245_1685# a_12079_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5277 vccd1 a_5123_5853# a_5291_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5278 a_6982_12533# a_6814_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5279 a_10915_22923# _0675_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5280 vssd1 a_25439_23163# a_25397_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5281 vssd1 a_22806_3829# a_22764_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5283 a_7465_18543# _0194_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5284 a_23237_10955# _0460_ a_23151_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5285 a_16737_12533# _0603_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X5286 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5287 vssd1 _0432_ _0787_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5288 vssd1 _0432_ a_4627_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5289 _0472_ a_14770_18517# a_14550_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5290 a_25674_17821# a_25401_17455# a_25589_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5291 cal_lut\[72\] a_28199_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5292 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5293 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd a_9687_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X5294 a_22277_14735# _0066_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5295 vssd1 a_12467_3579# a_12425_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5296 a_15186_1679# a_14913_1685# a_15101_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5297 a_7067_5162# _0318_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5298 a_8175_11445# cal_lut\[37\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X5299 vccd1 a_8546_15797# a_8473_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5300 a_17812_15529# _0551_ a_17710_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5301 a_17213_14735# a_16679_14741# a_17118_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5302 vssd1 a_22895_16519# _0689_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X5303 vssd1 a_10844_31029# net8 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5304 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5305 a_5050_29535# a_4882_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5306 a_11200_29575# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5307 vccd1 cal_lut\[118\] a_13122_6147# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5308 net20 a_14747_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5309 vssd1 a_22530_14709# a_22488_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5310 vccd1 a_27503_15253# a_27510_15553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5311 a_21085_8573# _0450_ a_21003_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5312 vssd1 clknet_0_io_in[0] a_5341_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5313 vccd1 cal_lut\[157\] a_20815_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5314 a_2887_25615# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X5315 a_3848_24135# _0411_ a_3990_24310# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5316 a_7060_31751# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5317 vccd1 a_20414_22325# a_20341_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5319 _0341_ a_25143_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X5320 a_9311_30511# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X5321 a_9763_26703# clknet_1_1__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X5322 a_24587_8573# cal_lut\[164\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X5323 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6007_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X5324 vccd1 _0814_ a_7847_28992# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5325 _0765_ _0722_ a_7565_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5326 _0100_ a_14287_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5327 a_12525_18231# _0836_ a_12688_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5328 a_9485_1501# a_8951_1135# a_9390_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5329 vssd1 clknet_1_1__leaf_io_in[0] a_4167_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5330 a_20440_13967# cal_lut\[24\] a_19865_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X5332 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5333 _0146_ a_9963_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5334 a_5073_6031# _0137_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5335 _0572_ a_12079_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5336 _0813_ a_5487_29217# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X5337 vssd1 a_7347_24501# _0751_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5338 a_11527_8207# _0493_ a_11705_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5339 a_24761_23983# _0061_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5340 vccd1 a_4128_20149# _0761_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X5341 a_5167_19631# ctr\[8\] _0739_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5342 a_9389_13103# cal_lut\[80\] a_8951_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5343 vssd1 a_15170_21237# a_15128_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5344 a_11794_8725# a_11587_8725# a_11970_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5345 vssd1 _0418_ a_2953_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X5346 vssd1 a_23823_20393# a_23830_20297# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5347 _0070_ a_26063_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5349 a_6277_7663# a_6007_8029# a_6187_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5350 a_4187_29245# a_3933_28918# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X5351 _0248_ a_26748_17705# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5352 vccd1 a_15595_10357# a_15511_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5353 a_24455_5639# a_24551_5461# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5354 a_21997_8213# a_21831_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5355 a_7369_28879# a_7133_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X5356 a_10876_28335# a_10497_28335# a_10779_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X5357 a_19862_4511# a_19694_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5358 vssd1 _0188_ a_5517_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5359 a_23021_16367# _0473_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X5360 vccd1 net26 a_14747_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5361 vccd1 a_18003_6941# a_18171_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5362 vccd1 a_20322_7775# a_20249_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5363 vssd1 a_13459_21807# _0216_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5364 vssd1 a_12597_7809# _0573_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X5366 a_21675_25437# a_20893_25071# a_21591_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5367 a_15554_3855# a_15281_3861# a_15469_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5368 a_20867_2986# _0337_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5370 vssd1 a_21299_27765# a_21257_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5371 vccd1 _0866_ a_18611_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5372 a_16300_16143# cal_lut\[96\] a_15725_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X5373 a_16845_14741# a_16679_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5374 cal_lut\[103\] a_20287_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5375 a_5617_15431# a_5713_15253# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X5376 a_19609_15279# _0023_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5378 a_11207_14954# _0844_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5379 a_21334_9951# a_21166_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5380 vccd1 a_23811_15431# _0656_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5381 a_8948_10703# _0476_ a_8758_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X5382 a_5675_3855# a_4811_3861# a_5418_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5383 vssd1 net24 a_4719_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5384 a_4981_28940# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5385 a_18605_6397# a_18335_6031# a_18515_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5386 a_7277_18543# a_7111_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5388 vssd1 a_11931_15645# a_12099_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5389 a_27859_15279# a_27639_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5390 a_7256_21237# _0669_ a_7476_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5391 vccd1 clknet_1_1__leaf__0380_ a_7491_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X5392 vccd1 a_4866_5599# a_4793_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5393 vssd1 a_9096_27221# _0817_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5394 a_5644_12533# ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.193 ps=1.41 w=1 l=0.15
X5395 a_9385_4373# _0451_ a_9638_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X5397 a_21085_11471# _0457_ a_21003_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5398 a_11660_5059# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5400 a_7648_21263# _0777_ a_7393_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5401 _0528_ a_20267_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5402 a_4381_21807# _0758_ a_4472_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5403 a_7888_32375# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5404 vssd1 net74 _0401_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5405 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5406 a_17187_13255# _0474_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X5407 a_23355_23671# _0470_ a_23683_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5408 a_22361_16367# a_21371_16367# a_22235_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5409 a_20522_3677# a_20083_3311# a_20437_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5410 vssd1 a_20763_1679# a_20931_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5411 a_7072_15797# net48 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5412 vccd1 a_17930_1653# a_17857_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5414 vccd1 a_25387_5161# a_25394_5065# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5415 vccd1 ctr\[4\] a_1679_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5416 _0385_ a_9835_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5417 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5418 a_24052_15113# a_23653_14741# a_23926_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5419 a_18130_3677# a_17857_3311# a_18045_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5420 a_22730_6031# a_22457_6037# a_22645_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5421 a_6081_8751# a_5915_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5422 vccd1 a_7994_16479# a_7921_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5423 a_3685_22325# clknet_0_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5424 a_6437_27247# a_5890_27521# a_6090_27221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5425 vssd1 a_5418_3829# a_5376_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5426 vssd1 a_15411_5755# a_15369_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5427 vccd1 a_7715_5461# _0328_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5428 vssd1 net45 a_19255_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5429 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5430 vssd1 a_27774_12533# a_27732_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5432 a_16757_7637# net17 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5433 a_15790_10089# _0549_ a_15541_9985# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5434 vccd1 a_15354_13621# a_15281_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5436 dbg_delay clknet_1_0__leaf_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5437 a_24823_11079# a_24919_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5438 a_18387_9527# a_18671_9513# a_18606_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5440 cal_lut\[51\] a_15687_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5441 a_5645_24527# _0793_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5442 a_22373_23145# _0466_ a_22457_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5443 cal_lut\[102\] a_16975_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5444 a_4893_25615# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X5445 vccd1 a_13939_21237# a_13855_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5446 _0063_ a_25787_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5447 a_15538_17567# a_15370_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5448 cal_lut\[76\] a_27003_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5449 _0734_ _0721_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X5451 vccd1 a_1641_28500# io_out[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5452 _0746_ _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=2.1 w=0.65 l=0.15
X5453 vssd1 a_15795_17821# a_15963_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5454 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5455 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5456 a_7936_25935# _0728_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X5457 a_4128_20149# _0447_ a_4348_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5458 vccd1 a_17286_14709# a_17213_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5460 vssd1 cal_lut\[68\] a_24041_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X5461 vssd1 a_19862_24501# a_19820_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5462 cal_lut\[37\] a_8143_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5463 vccd1 ctr\[2\] a_2695_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5464 a_23959_20553# a_23830_20297# a_23539_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5465 vssd1 a_14616_14709# _0872_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5466 a_12120_14851# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5467 vccd1 a_25271_24349# a_25439_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5468 _0494_ a_10046_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X5469 a_13028_7913# _0493_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5470 vccd1 a_12723_23439# net40 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5471 vccd1 a_4495_21495# _0781_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5472 vccd1 a_15494_19319# a_15370_19407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X5474 cal_lut\[50\] a_14307_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5475 vssd1 a_7631_17171# _0425_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5476 a_11717_16617# _0519_ a_11302_16519# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X5477 net37 a_22619_15253# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5478 a_11768_15939# cal_lut\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X5479 a_15531_4564# _0365_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5480 _0771_ net21 a_3241_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5481 a_18739_12559# a_17875_12565# a_18482_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5482 a_23505_26703# a_23167_26935# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5483 a_22891_20871# _0531_ a_23125_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5484 a_1945_15431# _0838_ a_2108_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5485 a_13309_16911# _0425_ a_13213_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X5486 a_21228_15529# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5487 a_15479_25615# a_15299_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5488 _0416_ a_2010_24759# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X5489 vccd1 _0233_ a_22659_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5490 vssd1 a_17159_22075# a_17117_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5491 a_27553_13647# a_27215_13879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5493 vssd1 a_8251_11293# a_8419_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5494 vccd1 _0744_ a_4984_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X5495 _0508_ a_19308_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5497 a_8491_18319# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5498 a_15391_27247# _0484_ a_15569_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5499 vssd1 _0425_ a_12577_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.213 pd=1.3 as=0.0878 ps=0.92 w=0.65 l=0.15
X5500 _0588_ a_10832_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X5501 a_10141_4221# a_9871_3855# a_10051_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5502 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5503 a_16281_5309# cal_lut\[179\] a_16209_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5504 vccd1 a_12870_13215# a_12797_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5505 vccd1 _0416_ a_1683_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5506 a_15452_19407# a_15115_19087# a_15370_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5507 vccd1 _0462_ a_20175_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5508 a_2582_14557# a_2143_14191# a_2497_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5509 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5510 a_4676_25223# _0827_ a_4818_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5511 a_6269_8751# _0139_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5514 a_13969_18218# _0539_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5516 a_21983_4943# _0687_ a_21889_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X5517 a_10961_5487# _0128_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5518 vccd1 cal_lut\[160\] a_20572_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5520 vssd1 io_in[7] a_1407_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X5521 _0699_ a_9034_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X5522 a_24761_22895# _0031_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5523 a_3017_27399# _0744_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5524 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5525 a_4793_5853# a_4259_5487# a_4698_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5526 a_6541_7125# a_6375_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5527 a_13529_22895# a_12539_22895# a_13403_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5528 _0834_ a_4003_30006# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X5529 _0547_ a_15483_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5530 vccd1 a_25042_19605# a_24971_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5531 vssd1 a_5123_5853# a_5291_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5532 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5533 a_1477_10901# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5534 vssd1 net32 a_19255_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5535 a_3017_27399# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X5536 vccd1 cal_lut\[45\] a_15531_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5537 vccd1 a_22863_1653# a_22779_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5538 a_24596_10703# _0510_ a_24105_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5539 vssd1 a_13139_7351# _0570_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5540 _0424_ a_2722_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5541 a_17861_26159# _0088_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5542 a_16991_27613# a_16293_27247# a_16734_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5543 vssd1 net33 a_25787_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5545 _0242_ a_21228_15529# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X5547 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5548 vccd1 cal_lut\[26\] a_23483_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5549 a_19759_3073# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X5550 a_15419_7119# a_14637_7125# a_15335_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5551 vssd1 a_8951_31599# net10 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5552 a_8383_22583# _0434_ a_8533_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5553 a_10839_15444# _0661_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5554 vccd1 _0792_ a_6381_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5555 a_12539_5056# cal_lut\[136\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5556 a_17117_27247# a_16127_27247# a_16991_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5558 a_7089_5487# a_6099_5487# a_6963_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5559 a_23781_20175# a_23443_20407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5560 a_16731_9813# net39 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5561 vssd1 _0077_ a_18029_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5562 temp1.capload\[6\].cap.Y clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5563 vssd1 _0773_ a_3749_30006# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X5564 vccd1 _0495_ a_16127_20288# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5565 a_19303_2375# a_19399_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5566 _0443_ a_19915_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5567 _0301_ a_14651_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X5568 vccd1 a_12898_10901# a_12827_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5569 a_6508_32375# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5570 a_9308_24847# dec1.i_ones a_9005_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5571 a_20648_3311# a_20249_3311# a_20522_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5572 a_18314_12559# a_18041_12565# a_18229_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5573 _0545_ a_15851_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5574 vssd1 _0352_ a_25463_12865# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5575 a_24941_9117# a_24407_8751# a_24846_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5576 vssd1 a_4931_24135# _0798_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5577 a_10294_13215# a_10126_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5578 vssd1 _0237_ a_23899_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5579 _0599_ a_16035_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5580 a_12955_25834# _0848_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5582 a_7716_25589# _0748_ a_7936_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5583 a_5583_6031# a_4885_6037# a_5326_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5585 a_20952_10499# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5586 _0206_ a_6546_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5587 _0031_ a_23763_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5588 vssd1 _0760_ a_4128_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X5589 a_9821_21263# _0557_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5590 vssd1 a_6055_10602# _0188_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5591 _0602_ a_16127_20288# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5592 vssd1 _0333_ a_16311_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5593 vssd1 a_22438_27765# a_22396_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5594 vssd1 a_11199_17607# a_11029_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X5595 a_20245_10927# a_19255_10927# a_20119_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5596 vssd1 _0747_ a_4713_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X5597 a_21872_20291# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5598 a_13700_15529# cal_lut\[78\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X5599 vssd1 a_20287_4667# a_20245_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5600 vssd1 a_18003_6941# a_18171_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5601 _0460_ a_20451_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5602 vccd1 a_17323_7663# _0505_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5603 vssd1 _0420_ a_3525_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5604 vssd1 net28 a_6375_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5605 vssd1 _0316_ a_4947_5249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5606 a_5083_11293# a_4903_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5607 a_11765_17973# net4 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X5608 a_2271_14735# a_1573_14741# a_2014_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5609 a_22185_1679# _0151_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5610 _0143_ a_6559_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5611 a_27701_12559# a_27167_12565# a_27606_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5612 vccd1 a_14123_23413# a_14039_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5613 vccd1 _0316_ a_9871_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5614 vccd1 a_17727_2589# a_17895_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5615 a_18142_28068# a_17935_28009# a_18318_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X5616 vssd1 _0446_ _0472_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5617 vssd1 _0563_ a_14345_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X5618 vccd1 _0395_ a_3335_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5619 vssd1 a_22235_16733# a_22403_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5620 a_16381_25071# a_15391_25071# a_16255_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5621 a_23056_17999# _0475_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5622 vssd1 a_15541_9985# _0550_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X5623 vssd1 a_6516_20871# _0736_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5624 a_14705_17620# _0555_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5625 _0706_ a_10607_24640# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5628 a_17129_23145# _0466_ a_16983_23047# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X5629 a_5250_13469# a_4811_13103# a_5165_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5630 _0856_ a_23207_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X5631 vssd1 a_15469_26935# _0270_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X5632 a_24971_19631# a_24842_19905# a_24551_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5633 vccd1 _0868_ a_23763_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5636 a_11896_24233# _0711_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5637 vccd1 net59 temp1.capload\[4\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5638 a_8477_14735# _0078_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5639 a_24473_9813# _0510_ a_24630_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5640 _0672_ a_10372_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5641 cal_lut\[47\] a_18355_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5642 a_11895_16367# _0625_ _0626_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X5643 vccd1 a_18298_3423# a_18225_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5644 vccd1 a_22898_6005# a_22825_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5645 a_18071_28169# a_17935_28009# a_17651_28023# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5646 vccd1 a_22695_8207# a_22863_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5648 vccd1 a_15354_1653# a_15281_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5649 a_16640_4373# net34 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5650 vccd1 a_13387_27515# a_13303_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5651 a_5359_22057# _0755_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5652 vccd1 _0363_ a_11527_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5653 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5654 a_22373_7663# _0505_ a_22291_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5655 vccd1 a_24459_8181# _0349_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5656 a_10607_9839# cal_lut\[189\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5657 vccd1 _0363_ a_13643_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5659 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5660 a_21970_18231# _0458_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X5661 vssd1 net40 a_13091_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5662 _0439_ _0438_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5663 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5664 vccd1 a_7060_31751# a_7011_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X5666 a_24971_13103# a_24835_13077# a_24551_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5667 vssd1 a_22719_27221# a_22726_27521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5668 vssd1 a_7073_25589# _0792_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5669 vssd1 a_18015_5639# _0598_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5671 vccd1 a_26514_13077# a_26443_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5672 _0764_ _0437_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5673 net45 a_15904_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5674 vssd1 net33 a_21831_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5675 vccd1 a_18291_16532# _0077_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5677 vssd1 a_23079_17607# _0480_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X5678 a_22961_17249# _0460_ a_22875_17249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5679 _0595_ a_17231_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5680 a_22553_3855# _0115_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5681 vssd1 cal_lut\[191\] a_12441_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5682 vssd1 net26 a_9963_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5683 vccd1 net44 a_19991_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5684 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5685 vccd1 _0514_ a_16771_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5686 a_20617_21263# a_20083_21269# a_20522_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5687 vssd1 a_11207_8903# cal_lut\[99\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5688 a_3656_25847# temp1.dac_vout_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5689 a_24473_9813# _0451_ a_24726_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X5690 vccd1 a_17543_9295# a_17711_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5691 a_23481_22717# a_23211_22351# a_23391_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5692 a_17543_9295# a_16845_9301# a_17286_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5693 vssd1 _0612_ a_16574_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X5694 vccd1 _0436_ a_7111_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5695 a_27521_15823# _0071_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5696 a_5359_22057# _0432_ a_5141_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5697 _0491_ a_14655_18115# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5698 a_11337_6575# a_11067_6941# a_11247_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5699 a_9503_19087# _0626_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X5700 a_9933_19061# _0590_ a_10313_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X5701 a_11891_11471# a_11711_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5702 a_19153_11837# _0505_ a_19071_11584# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5703 vccd1 a_20855_16911# a_21023_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5704 vccd1 _0459_ a_19807_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5705 vccd1 net27 a_4811_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5706 vccd1 _0841_ a_21555_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5707 a_15645_23817# a_14655_23445# a_15519_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5708 a_14287_22895# cal_lut\[9\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5711 vssd1 net1 a_13459_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5712 _0882_ a_8947_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X5713 a_19862_28447# a_19694_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5714 _0559_ a_18243_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5715 a_16105_12937# a_15115_12565# a_15979_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5716 a_19360_25993# a_18961_25621# a_19234_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5717 a_5365_23983# _0796_ a_4931_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5719 net32 a_17783_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5720 vccd1 a_1741_30199# a_1554_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5721 vccd1 a_15722_3829# a_15649_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5722 a_11471_5853# a_10607_5487# a_11214_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5724 vccd1 cal_lut\[39\] a_11891_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5726 _0225_ a_14375_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X5728 a_25011_21781# a_25295_21781# a_25230_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5729 a_21809_14191# a_20819_14191# a_21683_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5730 a_18027_19783# _0453_ a_18201_19659# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5732 vccd1 _0482_ a_16761_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5733 a_25455_17999# a_24757_18005# a_25198_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5734 vccd1 a_12299_3677# a_12467_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5735 _0530_ a_15299_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5736 vssd1 net9 a_11619_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5738 _0082_ a_17323_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5739 vssd1 _0422_ a_3072_19637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5740 vccd1 a_5843_3829# a_5759_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5741 a_7741_16367# _0001_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5742 _0485_ _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5743 a_2234_18793# _0420_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.148 ps=1.34 w=0.42 l=0.15
X5744 _0422_ a_1743_18259# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5745 vssd1 a_19308_17973# _0508_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5746 a_3171_26703# _0800_ _0801_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5747 vccd1 _0116_ a_24653_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5748 a_23355_10615# _0695_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X5749 a_6814_7119# a_6375_7125# a_6729_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5750 a_10688_23759# _0675_ a_10385_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5751 vccd1 a_5418_9269# a_5345_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5752 vccd1 a_22051_6941# a_22219_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5753 vssd1 temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5754 a_4725_14013# ctr\[4\] a_4653_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5755 vccd1 a_8543_30485# net11 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5756 vccd1 a_4584_23671# _0822_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5757 vccd1 ctr\[11\] a_6645_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5758 _0011_ a_18151_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5759 vccd1 a_7987_9514# _0120_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5760 vssd1 a_27710_15253# a_27639_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5761 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5762 vssd1 net81 a_14441_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5763 vssd1 a_12723_21807# _0237_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5765 vssd1 a_20690_3423# a_20648_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5766 a_14185_27497# cal_lut\[8\] a_14103_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5767 vssd1 a_15630_19743# a_15588_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5768 _0613_ a_16574_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X5769 a_5326_14709# a_5158_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5770 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6000_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X5771 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_1867_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5772 a_10961_14191# _0080_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5773 vccd1 io_in[0] a_6458_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5774 a_24235_4233# a_24106_3977# a_23815_4087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5777 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5778 a_20893_2223# a_20727_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5779 a_16853_8573# _0514_ a_16771_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5780 a_9779_27791# _0839_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5781 vssd1 clknet_1_0__leaf_io_in[0] a_5639_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5782 _0128_ a_10331_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5783 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5784 vssd1 a_17599_6039# _0514_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5785 a_9772_30287# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X5786 vccd1 a_27774_12533# a_27701_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5787 cal_lut\[63\] a_25991_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5788 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5789 vccd1 a_1919_20693# _0762_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5790 vccd1 a_15561_18231# _0274_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X5791 a_13035_3855# a_12337_3861# a_12778_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5792 vccd1 _0265_ a_21279_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5793 a_2505_10703# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5794 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5796 a_16737_13621# _0597_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5797 a_13254_9295# a_12815_9301# a_13169_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5798 vssd1 a_12525_18231# _0846_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X5799 a_17033_14735# _0022_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5800 a_25931_8725# cal_lut\[165\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X5801 a_16734_27359# a_16566_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5802 a_2959_25071# _0806_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X5803 a_26309_20553# a_25762_20297# a_25962_20452# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5805 a_10659_7637# net39 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5806 a_5158_14735# a_4885_14741# a_5073_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5807 a_7741_6575# _0126_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5808 _0321_ a_5404_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5809 vccd1 _0359_ a_27903_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5811 vccd1 dec1.i_ones a_9275_28023# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5812 cal_lut\[63\] a_25991_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5813 vccd1 a_6982_12127# a_6909_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5814 a_9496_31599# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X5815 _0542_ a_15023_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5816 a_4408_29245# _0800_ a_4187_28918# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5817 vccd1 cal_lut\[181\] a_9131_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5818 a_7079_24233# _0724_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5819 vssd1 a_17286_14709# a_17244_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5820 a_18225_3677# a_17691_3311# a_18130_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5821 a_22825_6031# a_22291_6037# a_22730_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5822 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5823 a_17283_28853# a_17459_29185# a_17411_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X5824 _0087_ a_21279_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5825 a_20690_18517# _0442_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X5826 a_19940_19881# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5827 a_15281_1679# a_14747_1685# a_15186_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5828 vssd1 a_13882_4917# a_13840_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5830 vccd1 _0713_ a_8951_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5831 a_15220_23817# a_14821_23445# a_15094_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5834 a_27606_17821# a_27167_17455# a_27521_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5835 vccd1 a_22235_22173# a_22403_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5836 vccd1 a_4995_17999# net21 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5837 a_5165_3855# _0134_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5838 vccd1 temp1.i_precharge_n a_2778_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5839 vccd1 a_17875_4399# _0290_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5841 vssd1 a_27503_15253# a_27510_15553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5842 vssd1 a_27755_9117# a_27923_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5843 a_27701_11471# a_27167_11477# a_27606_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5844 _0488_ a_14103_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5845 vccd1 a_22863_27765# a_22779_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5846 a_27333_9839# a_27167_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5847 a_10347_25071# _0732_ a_10197_25223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X5848 io_out[1] a_1551_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5849 a_12437_19407# cal_lut\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X5850 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_2044_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X5852 vccd1 a_8419_13371# a_8335_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5854 a_3488_9001# cal_lut\[140\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X5856 vssd1 a_12311_11079# cal_lut\[98\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5857 a_9607_29257# a_9471_29097# a_9187_29111# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5858 _0665_ _0631_ a_12165_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5859 vssd1 _0678_ a_11508_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X5860 _0279_ a_14375_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X5863 a_17094_20407# _0577_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X5864 a_23850_17277# a_23535_17143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5865 a_9275_28023# ctr\[12\] a_9509_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5866 vssd1 cal_lut\[48\] a_19664_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5867 vccd1 a_18671_9513# a_18678_9417# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5868 vssd1 a_15135_1403# a_15093_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5869 a_21878_17143# _0691_ a_22181_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X5870 vccd1 a_20287_15547# a_20203_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5871 a_8723_17130# _0842_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5872 vssd1 _0446_ _0384_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5873 _0851_ a_20779_15253# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5875 vccd1 cal_lut\[161\] a_25783_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5877 vssd1 a_13571_25339# a_13529_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5878 vccd1 a_10659_3829# _0314_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5879 a_26778_22173# a_26339_21807# a_26693_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5880 a_12926_7913# _0571_ a_12846_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X5881 net29 a_11527_9303# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5882 a_11508_20719# _0676_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5883 vccd1 a_11366_28588# dbg_result[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5884 vssd1 a_16255_25437# a_16423_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5885 a_22891_20871# _0531_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5886 a_25773_8207# _0165_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5887 _0492_ _0491_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5888 vccd1 _0808_ a_3891_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X5889 a_17401_24759# cal_lut\[42\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X5890 _0454_ a_18519_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X5891 a_24573_7125# a_24407_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5892 vssd1 a_16219_25623# net47 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5893 a_13261_21263# _0039_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5894 a_14818_5853# a_14545_5487# a_14733_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5895 a_17095_16055# a_17191_16055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5896 vssd1 net23 a_4811_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5897 vccd1 cal_lut\[176\] a_25047_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5898 a_9835_26703# _0460_ a_9763_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.0672 ps=0.85 w=0.64 l=0.15
X5899 a_23211_5263# cal_lut\[116\] a_23117_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5900 vssd1 a_2009_30676# io_out[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5901 _0715_ a_9167_21601# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X5902 vssd1 a_13512_13621# _0576_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5904 a_25927_13255# a_26023_13077# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5905 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5906 a_16534_5737# _0614_ a_16220_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X5907 vssd1 a_2805_30265# a_2739_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5908 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5909 a_23811_4564# _0296_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5910 cal_lut\[143\] a_5567_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5911 vccd1 net6 a_3155_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5912 a_5326_6005# a_5158_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5913 a_17674_29789# a_17427_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5914 vssd1 _0239_ a_25787_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5916 _0592_ dbg_result[5] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5917 vssd1 net22 a_2121_21623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0536 ps=0.675 w=0.42 l=0.15
X5918 vccd1 net9 a_11527_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X5919 a_8730_14709# a_8562_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5920 vccd1 _0363_ a_15299_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5921 vccd1 a_10827_7119# a_10995_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5922 a_5345_9295# a_4811_9301# a_5250_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5924 a_19889_14191# _0531_ a_19807_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5925 _0450_ a_17651_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5926 a_2552_31287# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5927 a_12426_2589# a_11987_2223# a_12341_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5928 a_19683_2197# net31 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5929 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5930 a_20671_22351# a_19973_22357# a_20414_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5931 a_12310_10615# _0655_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X5932 a_19605_26709# a_19439_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5933 vccd1 a_21115_3579# a_21031_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5934 cal_lut\[186\] a_18355_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5935 a_26026_8181# a_25858_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5937 vccd1 _0237_ a_20727_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5938 a_2563_23957# clknet_1_0__leaf_temp1.i_precharge_n a_2772_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X5939 _0031_ a_23763_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5940 a_21879_16055# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X5941 cal_lut\[132\] a_14675_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5942 vssd1 a_18597_13077# _0456_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5944 vssd1 a_18119_7637# a_18126_7937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5945 vccd1 a_25623_17973# a_25539_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5947 a_18182_17027# _0851_ a_18100_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5949 vssd1 _0464_ _0492_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5950 a_11895_16367# cal_lut\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5951 a_16031_3311# cal_lut\[179\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X5952 a_6940_7497# a_6541_7125# a_6814_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5953 vccd1 dbg_result[1] a_19915_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X5954 a_15002_10383# a_14729_10389# a_14917_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5956 vssd1 a_2271_12559# a_2439_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5957 a_23683_27081# a_23554_26825# a_23263_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5958 vccd1 a_13571_23163# a_13487_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5959 vssd1 a_6522_8863# a_6480_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5961 cal_lut\[116\] a_23231_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5962 ctr\[5\] a_5843_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5963 vccd1 a_11847_3073# a_11671_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X5964 vccd1 net8 a_10055_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X5965 a_2462_25935# _0418_ a_2372_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X5966 vccd1 a_14703_25236# _0093_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5967 a_11609_21379# _0670_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5968 _0403_ _0814_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5969 a_20065_1685# a_19899_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5970 cal_lut\[86\] a_23231_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5971 vccd1 a_12219_17130# _0005_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5972 vccd1 a_25463_12865# a_25287_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X5974 vssd1 _0362_ a_25419_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5975 a_9091_29111# a_9187_29111# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5976 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5977 a_13144_22325# _0838_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5978 vccd1 a_21223_19997# a_21391_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5979 vssd1 net41 a_9595_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5980 a_9678_24233# _0723_ a_9372_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5981 vccd1 cal_lut\[22\] a_14778_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5982 a_12935_2589# a_12153_2223# a_12851_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5983 a_15255_28500# _0270_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5984 a_12794_27613# a_12355_27247# a_12709_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5986 _0536_ a_20359_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5987 vssd1 a_27595_13865# a_27602_13769# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5988 vssd1 a_22441_21237# _0639_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X5989 a_27149_18005# a_26983_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5990 vccd1 a_26911_16635# a_26827_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5991 vssd1 net29 a_14563_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5992 vssd1 a_15071_13268# _0010_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5993 a_6828_28111# _0408_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5994 a_3785_17999# _0421_ a_4143_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5995 a_4091_15279# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X5996 a_13380_9673# a_12981_9301# a_13254_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5997 vccd1 _0422_ a_2371_18523# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5998 _0176_ a_25419_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5999 a_19746_27497# _0222_ a_19664_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6000 _0387_ a_4351_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X6001 vccd1 net20 a_19807_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6002 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6003 vssd1 a_6245_21781# _0820_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6004 vssd1 a_6246_16503# a_6184_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X6005 vssd1 a_14139_4943# a_14307_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6006 a_4606_27791# a_4167_27797# a_4521_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6007 vccd1 a_16635_26324# _0042_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6008 _0647_ a_15378_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X6009 vssd1 a_18698_19319# _0461_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X6010 a_18383_5175# _0514_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6011 vccd1 a_27774_11445# a_27701_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6012 vccd1 a_13127_13469# a_13295_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6013 a_22961_9867# _0450_ a_22875_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6014 _0831_ a_2839_27221# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6015 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X6016 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6375_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6017 a_5487_29217# ctr\[9\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6018 vccd1 a_5503_27399# ctr\[7\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6019 net46 a_18111_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6020 vssd1 _0032_ a_25849_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6021 a_6982_7093# a_6814_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6022 a_7741_13103# _0019_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6023 _0447_ a_14103_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X6024 a_15281_12565# a_15115_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6025 vssd1 _0246_ a_10501_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6026 a_12455_18793# net15 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X6027 a_8929_2057# a_7939_1685# a_8803_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6029 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X6032 a_25585_8213# a_25419_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6033 vssd1 net36 a_24407_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6034 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6035 _0003_ a_9595_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6037 a_11605_16055# cal_lut\[4\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X6038 _0374_ a_7291_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X6039 a_9033_12879# cal_lut\[19\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6040 a_4521_27791# _0207_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6041 a_5841_27613# a_5503_27399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6042 _0429_ _0422_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6043 vccd1 a_19303_16519# _0606_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6045 vccd1 _0841_ a_23579_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6046 a_3056_28111# temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X6047 vssd1 a_20039_18695# _0612_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6048 cal_lut\[53\] a_20471_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6049 a_8293_1679# _0180_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6050 _0684_ a_21831_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X6051 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6052 a_2376_30199# _0800_ a_2518_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X6054 vccd1 cal_lut\[182\] a_9591_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6055 a_5547_21263# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X6056 vccd1 _0495_ a_10699_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6057 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6058 vccd1 a_2991_15797# a_2907_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6059 cal_lut\[27\] a_24243_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6060 _0192_ _0839_ a_5825_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6063 _0374_ a_7291_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6064 vccd1 a_14583_26677# a_14499_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6066 _0074_ a_24315_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6068 a_15479_3677# a_15299_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6069 _0116_ a_23671_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6070 a_16153_8751# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6071 vssd1 net10 a_9311_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X6072 a_14550_18793# _0425_ a_14353_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6073 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6074 vccd1 cal_lut\[163\] a_24035_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6075 a_12981_9301# a_12815_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6076 a_22895_16519# _0688_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X6077 vccd1 cal_lut\[5\] a_11717_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6078 a_2271_12559# a_1407_12565# a_2014_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6079 vccd1 net33 a_22291_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6081 a_24972_22895# a_24573_22895# a_24846_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6083 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6084 a_17564_24643# cal_lut\[42\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X6085 a_7239_7119# a_6541_7125# a_6982_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6086 a_6552_31375# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X6087 vccd1 net27 a_3799_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6088 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6089 _0250_ a_27024_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6090 vssd1 a_22898_6005# a_22856_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6091 temp1.capload\[0\].cap.Y clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6092 a_14163_8903# _0472_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6093 a_14103_25437# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6094 a_3859_7337# net24 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6095 a_17498_29397# a_17291_29397# a_17674_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6096 a_10664_13763# cal_lut\[80\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X6098 vccd1 clknet_1_1__leaf__0380_ a_9595_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.173 ps=1.82 w=0.64 l=0.15
X6099 a_2782_20719# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X6100 vccd1 _0817_ _0826_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6101 a_2866_14013# ctr\[1\] a_2777_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0619 ps=0.715 w=0.42 l=0.15
X6103 a_7465_14191# _0036_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6104 vssd1 _0483_ a_16189_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6105 cal_lut\[135\] a_5843_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6106 vssd1 net1 a_13367_10391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6108 vccd1 a_3117_12533# _0203_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6109 vccd1 a_6982_12533# a_6909_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6110 a_6823_17999# a_6541_18005# a_6729_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X6111 a_5377_16143# ctr\[2\] _0192_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6112 _0198_ a_3851_15253# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6113 _0694_ a_9963_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X6115 _0819_ _0437_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6118 a_2413_23759# net22 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6119 a_7553_13103# a_7387_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6120 a_17427_29423# a_17291_29397# a_17007_29397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6121 vccd1 a_20775_18231# _0526_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6122 a_25137_16367# a_24867_16733# a_25047_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X6123 a_17560_4917# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6125 vssd1 a_7131_5755# a_7089_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6126 cal_lut\[164\] a_25439_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6127 vccd1 a_13679_9295# a_13847_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6128 a_24057_12559# a_23719_12791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6129 vssd1 a_17555_19319# _0580_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6130 vccd1 a_7523_24833# a_7347_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6132 a_12552_2223# a_12153_2223# a_12426_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6133 vccd1 cal_lut\[128\] a_10362_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6134 a_22638_25437# a_22365_25071# a_22553_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6135 vccd1 a_6062_11039# a_5989_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6136 a_7607_2589# a_6743_2223# a_7350_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
R17 vssd1 net63 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6137 vssd1 a_8251_29789# a_8419_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6139 a_19437_18543# dbg_result[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X6140 vssd1 a_25531_15797# a_25489_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6141 vssd1 _0431_ a_6363_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X6142 a_15851_8320# cal_lut\[180\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6144 vssd1 cal_lut\[169\] a_24596_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X6145 vccd1 a_27371_22075# a_27287_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6146 vssd1 clknet_0__0380_ a_6537_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6147 vssd1 a_20579_9295# a_20747_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6148 a_6062_11039# a_5894_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6149 vccd1 a_20119_11293# a_20287_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6150 a_19973_28879# a_19439_28885# a_19878_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6151 a_7101_23759# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6152 vssd1 a_26026_8181# a_25984_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6153 vccd1 _0437_ a_7393_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6154 vccd1 ctr\[4\] a_4491_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6155 a_26023_13077# a_26307_13077# a_26242_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6156 a_10317_1679# _0182_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6157 _0165_ a_25143_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6158 a_4238_10205# a_3965_9839# a_4153_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6160 vccd1 a_11019_2197# a_10843_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6161 a_20775_5639# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6162 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6164 vssd1 _0443_ a_19373_21835# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6165 a_22396_23817# a_21997_23445# a_22270_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6166 vccd1 cal_lut\[89\] a_18642_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6167 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6168 cal_lut\[1\] a_4831_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6169 _0817_ a_9096_27221# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X6170 vccd1 a_15243_5853# a_15411_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6171 a_2092_31287# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X6172 a_20387_26703# a_19605_26709# a_20303_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6173 vccd1 _0771_ a_2605_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6174 _0723_ a_8397_20983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6175 vccd1 net44 a_18519_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6176 a_3685_22325# clknet_0_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6177 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6178 a_20775_27412# _0228_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6179 vssd1 a_7251_1898# _0186_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6182 a_1464_23957# _0791_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.265 ps=1.47 w=0.65 l=0.15
X6183 a_26479_16042# _0249_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6184 a_23683_23439# cal_lut\[86\] a_23481_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6185 vccd1 a_18751_23671# _0620_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6186 a_24159_19087# a_23377_19093# a_24075_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6187 a_11547_24847# _0706_ _0714_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6188 a_20775_18231# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6189 a_24761_23983# _0061_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6190 cal_lut\[143\] a_5567_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6191 _0609_ a_16373_13077# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X6193 a_8102_3855# a_7829_3861# a_8017_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6194 a_4435_32463# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X6195 a_13275_20175# _0438_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6197 vccd1 a_19383_16911# a_19551_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6198 vssd1 a_21883_1109# _0335_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X6199 a_8105_1685# a_7939_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6200 vssd1 a_23723_25045# _0264_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X6201 a_22729_22895# cal_lut\[55\] a_22291_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6202 a_20437_3311# _0156_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6203 a_5207_5853# a_4425_5487# a_5123_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6205 ctr\[9\] a_5475_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6206 a_4733_16367# clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6207 a_3575_7351# a_3859_7337# a_3794_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6208 _0741_ _0420_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X6209 vccd1 _0307_ a_14195_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6210 a_8268_24501# _0721_ a_8397_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6212 a_15439_17130# _0274_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6213 vssd1 net10 a_7663_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6214 a_13537_15431# _0246_ a_13700_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6216 vccd1 _0746_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6217 vccd1 a_22438_8181# a_22365_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6218 vccd1 a_24823_11079# cal_lut\[177\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6219 vccd1 a_11458_27500# dbg_result[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X6220 vssd1 a_15687_23413# a_15645_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6221 vccd1 _0839_ a_7557_28640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X6222 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6223 vssd1 a_13751_16911# _0477_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6224 a_8105_15829# a_7939_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6225 vssd1 a_15519_29789# a_15687_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6226 a_18291_28157# a_18071_28169# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6228 a_22457_23145# cal_lut\[85\] a_22373_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6229 a_18271_1679# a_17489_1685# a_18187_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6230 a_6909_10389# a_6743_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6231 a_4345_11791# _0808_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6232 a_22165_10357# _0632_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X6233 vccd1 _0483_ a_8675_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X6234 vssd1 a_16147_12533# a_16105_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6235 a_13629_28879# _0049_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6238 a_10202_15797# a_10034_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6239 vssd1 cal_lut\[185\] a_16949_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6241 a_8383_22583# _0776_ a_8617_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X6242 a_20437_21263# _0065_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6243 a_13698_23413# a_13530_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6244 vccd1 _0418_ a_2695_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X6245 vccd1 _0427_ a_4265_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6246 vccd1 _0390_ a_4245_14796# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X6247 vssd1 a_18475_19783# _0579_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6248 vccd1 net8 a_10239_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6249 cal_lut\[3\] a_8971_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6250 vccd1 _0841_ a_12263_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6251 a_19426_20719# cal_lut\[52\] a_19345_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X6252 _0195_ net72 a_5377_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6253 vccd1 cal_lut\[77\] a_17538_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6254 cal_lut\[50\] a_14307_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6255 vssd1 cal_lut\[55\] a_22009_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6256 vssd1 _0237_ a_9823_15041# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6257 vssd1 a_26123_14165# a_26130_14465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6258 _0197_ _0386_ a_9779_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6259 vccd1 a_22530_14709# a_22457_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6260 vccd1 a_20119_4765# a_20287_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6261 vssd1 a_9815_1501# a_9983_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6262 vssd1 _0425_ a_8556_20725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
X6263 vccd1 _0453_ a_18763_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6264 vssd1 a_8419_16635# a_8377_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6265 vccd1 a_18539_26427# a_18455_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6266 a_24867_11471# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6267 vssd1 a_18355_24251# a_18313_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6268 vssd1 _0472_ a_14287_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X6269 a_10953_2057# a_9963_1685# a_10827_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6270 a_2564_25045# _0807_ a_2959_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6271 cal_lut\[65\] a_20839_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6272 a_25355_9117# a_24573_8751# a_25271_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6273 a_14920_9615# cal_lut\[100\] a_14345_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X6274 _0872_ a_14616_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X6276 a_13530_23439# a_13257_23445# a_13445_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6277 a_25858_8207# a_25419_8213# a_25773_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6278 a_20893_25071# a_20727_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6279 a_26946_21919# a_26778_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6280 vssd1 a_22523_2999# cal_lut\[153\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6281 vssd1 net39 a_3339_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X6282 a_10607_24640# _0682_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6283 cal_lut\[125\] a_15135_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6284 a_11776_29673# a_11527_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X6285 vccd1 a_14139_28879# a_14307_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6286 cal_lut\[65\] a_20839_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6287 _0234_ a_19940_19881# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6289 a_22471_2589# a_22291_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6290 vccd1 a_2014_12533# a_1941_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6291 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6292 vccd1 net7 a_1683_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6293 vccd1 a_14986_5599# a_14913_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6294 a_20775_18231# _0459_ a_21009_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6297 _0034_ a_14747_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6299 a_23631_17143# a_23915_17129# a_23850_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6300 a_5541_9839# a_5271_10205# a_5451_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X6301 vssd1 _0644_ a_15378_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X6302 vccd1 a_4679_19319# _0742_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6303 vssd1 cal_lut\[102\] a_18145_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6304 a_10740_29575# net8 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X6305 vssd1 _0627_ a_10247_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6307 a_14277_13967# _0501_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6308 a_12577_20495# _0447_ a_12463_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.137 ps=1.07 w=0.65 l=0.15
X6309 vssd1 net35 a_19715_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6310 a_13763_9295# a_12981_9301# a_13679_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6311 io_out[4] a_1464_23957# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6313 a_16692_21807# a_16293_21807# a_16566_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6314 a_12794_27613# a_12521_27247# a_12709_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6315 a_7849_26819# ctr\[11\] a_7753_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6316 a_17677_25071# _0046_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6317 vccd1 a_15595_21237# a_15511_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6318 a_13119_14557# a_12337_14191# a_13035_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6319 vccd1 a_26203_6250# _0161_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6320 _0236_ a_23299_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X6321 vccd1 a_25927_13255# cal_lut\[175\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6323 vccd1 a_14699_6549# a_14523_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6324 vccd1 net43 a_25971_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6325 a_10129_1685# a_9963_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6326 _0871_ a_18100_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X6327 a_1651_14165# ctr\[0\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X6328 cal_lut\[8\] a_13387_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6329 vccd1 _0363_ a_16679_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6330 vccd1 a_27755_9117# a_27923_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6331 vccd1 a_16975_11195# a_16891_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6332 vssd1 a_12594_2335# a_12552_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6333 net27 a_3707_9303# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X6335 vssd1 a_13291_18909# _0474_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6336 vssd1 _0871_ a_18611_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6337 a_2317_16911# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6338 a_13968_17218# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X6339 vccd1 a_10551_13469# a_10719_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6340 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6341 a_4443_18793# _0420_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6342 a_26869_16367# a_25879_16367# a_26743_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6343 vssd1 a_20046_28853# a_20004_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6344 vccd1 _0330_ a_18795_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6345 a_20705_7663# a_19715_7663# a_20579_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6346 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6347 a_21975_19605# a_22259_19605# a_22194_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6348 a_19383_16911# a_18519_16917# a_19126_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6349 a_26058_14191# a_25743_14343# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6350 vccd1 a_19862_15391# a_19789_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6351 cal_lut\[159\] a_23323_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6352 vssd1 dbg_result[2] a_13459_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6353 vccd1 a_5617_15431# net77 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6354 a_5813_22895# _0750_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X6356 _0515_ _0491_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6357 a_4003_30006# _0801_ a_4003_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6358 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6360 _0483_ a_15207_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.175 ps=1.26 w=0.65 l=0.15
X6361 vccd1 net31 a_20083_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6362 vssd1 a_23055_23047# _0470_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6363 a_22843_4399# cal_lut\[152\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6364 a_17427_29423# a_17298_29697# a_17007_29397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6365 a_10423_17455# _0662_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X6366 a_20775_14967# _0443_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6367 vssd1 a_23361_9985# _0659_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X6369 a_11693_8207# cal_lut\[123\] a_11609_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6370 a_23757_11177# _0509_ a_23959_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6371 _0304_ a_10235_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6372 a_19053_16911# a_18519_16917# a_18958_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6373 a_16761_24527# cal_lut\[94\] a_16679_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6374 vssd1 a_21327_24746# _0084_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6375 vssd1 a_10627_15797# a_10585_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6376 a_14591_15823# a_13809_15829# a_14507_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6379 vssd1 cal_lut\[28\] a_18100_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6380 a_9853_13103# a_9687_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6381 net10 a_8951_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6382 vssd1 a_13144_22325# _0863_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6383 a_19333_9991# cal_lut\[105\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X6384 a_6269_29423# _0209_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6385 a_8251_6941# a_7553_6575# a_7994_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6386 a_4491_13879# ctr\[5\] a_4725_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6387 a_24770_5487# a_24455_5639# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6388 a_10857_21781# _0672_ a_11014_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X6389 a_12437_19407# net4 _0556_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6391 a_13955_23439# a_13257_23445# a_13698_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6392 a_22365_8207# a_21831_8213# a_22270_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6393 vssd1 net35 a_20727_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6394 a_7755_25321# _0724_ _0734_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X6395 a_7067_5162# _0318_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6396 _0504_ a_8951_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6397 a_4477_22057# _0757_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X6398 cal_lut\[11\] a_15779_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6399 net33 a_23211_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6400 a_21327_24746# _0262_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6401 vccd1 _0453_ a_18151_21271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X6402 a_6611_22583# _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X6403 a_27732_16201# a_27333_15829# a_27606_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6404 vccd1 _0393_ a_3151_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X6405 vccd1 _0505_ a_19255_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6407 a_1919_20693# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6408 vccd1 cal_lut\[36\] a_15623_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6409 vssd1 _0872_ a_19333_25223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6410 cal_lut\[11\] a_15779_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6412 a_6269_8751# _0139_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6413 a_17927_4917# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6414 a_1913_28023# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X6416 a_9773_25935# _0720_ a_9555_25847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6417 vccd1 net47 a_22199_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6418 a_12959_15253# cal_lut\[96\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X6420 vssd1 a_11579_25045# _0731_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6421 a_14139_28879# a_13275_28885# a_13882_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6422 vccd1 net1 a_13459_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X6423 vccd1 _0352_ a_26983_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6424 _0059_ a_20359_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6425 a_11029_17429# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X6426 a_6729_14735# _0192_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6427 cal_lut\[115\] a_21759_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6428 a_23903_18695# _0460_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6429 vccd1 _0838_ a_13459_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X6430 a_14507_3855# a_13643_3861# a_14250_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6431 a_19881_7663# a_19715_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6432 _0405_ ctr\[10\] a_7194_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X6434 a_8951_2589# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6435 a_4461_25913# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6437 vssd1 _0820_ a_5416_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6438 vssd1 a_7775_10357# a_7733_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6439 a_10715_21263# _0591_ a_10521_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6440 a_26835_18909# a_26137_18543# a_26578_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6441 a_4977_13103# a_4811_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6442 a_23282_8029# a_23009_7663# a_23197_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6443 a_19667_18517# dbg_result[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6444 vccd1 cal_lut\[75\] a_23056_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6445 vccd1 net64 temp1.capload\[9\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6446 a_1937_6549# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6447 vssd1 a_16983_23047# _0578_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6448 a_3882_16911# net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6450 temp1.capload\[14\].cap.Y net54 a_1677_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6452 a_14913_5853# a_14379_5487# a_14818_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6453 a_16550_11039# a_16382_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6454 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_3056_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X6455 net80 a_16311_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6457 temp1.dac_vout_notouch_ net14 a_11776_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X6459 vccd1 net34 a_24407_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6460 _0698_ a_8951_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6461 vssd1 a_14250_3829# a_14208_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6463 vssd1 a_15243_5853# a_15411_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6464 cal_lut\[138\] a_5751_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6466 vssd1 cal_lut\[141\] a_5449_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6467 vccd1 net10 a_7203_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6468 a_25103_5175# a_25387_5161# a_25322_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6469 vssd1 net27 a_5915_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6470 a_2107_19631# _0428_ a_1551_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6471 a_24201_19465# a_23211_19093# a_24075_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6472 _0626_ _0625_ a_11895_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6474 a_16859_1501# a_16679_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6475 a_25984_8585# a_25585_8213# a_25858_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6477 vssd1 _0056_ a_24101_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6478 a_5583_6031# a_4719_6037# a_5326_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6479 vccd1 _0450_ a_10607_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6480 a_27337_17999# _0070_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6481 a_4600_31849# a_4351_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X6482 a_1867_23759# clknet_1_1__leaf_io_in[0] _0415_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6483 vssd1 _0411_ a_1932_22711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
X6484 cal_lut\[35\] a_16055_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6485 a_20848_13353# _0456_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6486 vccd1 a_15535_24501# _0273_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X6487 vccd1 a_12355_21271# _0266_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6488 vssd1 _0649_ a_11527_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6489 vccd1 a_15795_17821# a_15963_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6491 a_14542_1501# a_14269_1135# a_14457_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6492 a_24551_13077# a_24842_13377# a_24793_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6493 vccd1 _0841_ a_13183_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6495 a_9008_27907# dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X6496 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6497 vccd1 a_21879_19783# cal_lut\[59\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6498 a_5043_24566# _0798_ a_4584_24759# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X6499 vccd1 a_15812_9269# net35 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6500 vccd1 _0280_ a_16035_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6501 a_7875_27613# a_7093_27247# a_7791_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6502 vccd1 a_13714_19407# _0495_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6503 a_5158_6031# a_4719_6037# a_5073_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6504 vssd1 a_20855_16911# a_21023_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6505 vssd1 _0843_ a_9595_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6506 vccd1 clknet_0_io_in[0] a_5341_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6507 a_11877_26709# a_11711_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6509 a_5105_25045# _0747_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6510 vssd1 a_4222_12533# a_4180_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6511 a_6375_8207# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6512 a_11587_8725# net29 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6513 vssd1 a_22165_10357# _0635_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X6514 a_5993_16367# _0193_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X6515 _0502_ a_18645_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X6516 vccd1 a_21299_27765# a_21215_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6517 _0678_ a_10331_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6519 vccd1 _0245_ a_25327_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6521 a_22645_6031# _0158_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6525 vssd1 a_17831_24746# _0046_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6526 a_25489_16201# a_24499_15829# a_25363_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6527 vssd1 a_7005_4551# _0315_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X6528 a_23395_8751# cal_lut\[165\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6529 vccd1 a_21759_2491# a_21675_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6530 vccd1 a_9929_10357# _0516_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6531 a_7380_31375# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X6532 vssd1 a_11366_28588# dbg_result[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X6533 a_18475_5639# _0443_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6534 a_11014_22057# _0674_ a_10857_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6535 vccd1 a_7775_2491# a_7691_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6536 vccd1 _0460_ a_14287_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6537 vssd1 a_2750_20407# a_2722_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6539 a_23189_25071# a_22199_25071# a_23063_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6540 vccd1 a_19126_16885# a_19053_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6541 vssd1 a_20119_4765# a_20287_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6542 vccd1 _0707_ a_10699_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X6543 vssd1 _0232_ a_23579_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6544 a_21334_2335# a_21166_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6546 _0422_ a_1743_18259# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6547 a_2685_13103# _0411_ _0389_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6549 a_3151_14735# _0394_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6550 a_7350_2335# a_7182_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6552 a_17507_5487# cal_lut\[131\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6553 a_27517_7119# a_26983_7125# a_27422_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6554 vssd1 a_1743_18259# _0422_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X6556 a_4528_14735# _0398_ _0205_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X6557 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10488_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X6558 a_2564_25045# _0807_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X6559 vssd1 a_11581_21781# _0674_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6560 a_19525_3311# a_19255_3677# a_19435_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X6561 vssd1 _0015_ a_25389_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6562 a_21334_2335# a_21166_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6563 vssd1 a_17875_16367# net44 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6565 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_2879_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6566 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6567 _0057_ a_23579_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6569 a_9487_26159# clknet_1_1__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0567 ps=0.69 w=0.42 l=0.15
X6570 a_1625_19087# _0421_ a_1541_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6571 vccd1 cal_lut\[28\] a_18182_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6572 vccd1 a_18369_18337# _0475_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X6573 a_11421_15279# _0004_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6574 vccd1 _0710_ a_10915_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6576 a_7102_21807# _0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6577 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6578 vssd1 a_9983_14459# a_9941_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6579 a_16063_3855# a_15281_3861# a_15979_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6580 vccd1 cal_lut\[114\] a_20758_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6582 vssd1 a_6427_11445# _0377_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X6583 temp1.dac_vout_notouch_ net14 a_9772_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X6584 a_10809_19605# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6586 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6587 vccd1 net57 temp1.capload\[2\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6588 a_23211_21263# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6589 a_14967_8029# a_14269_7663# a_14710_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6590 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6591 _0370_ a_11707_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X6592 _0322_ a_6555_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6593 a_17946_26525# a_17507_26159# a_17861_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6594 vssd1 a_13459_17455# _0438_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6596 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6597 vccd1 net11 a_9779_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6598 vccd1 a_23754_26980# a_23683_27081# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6599 temp1.i_precharge_n a_1683_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6600 a_7239_14735# a_6375_14741# a_6982_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6601 vccd1 _0422_ _0426_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6602 a_2695_14013# ctr\[0\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.109 ps=1.36 w=0.42 l=0.15
X6603 vssd1 a_17094_20407# _0587_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X6604 cal_lut\[128\] a_10075_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6605 vssd1 cal_lut\[74\] a_23489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X6606 vccd1 a_27802_13924# a_27731_14025# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6607 vccd1 a_8270_3829# a_8197_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6609 a_9275_15444# _0256_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6610 a_7291_25615# _0733_ a_7073_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6611 a_18900_14025# a_18501_13653# a_18774_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6612 a_12759_17821# a_12061_17455# a_12502_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6613 a_26138_12381# a_25891_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6614 a_20322_7775# a_20154_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6615 a_5871_10004# _0321_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6616 a_13211_13469# a_12429_13103# a_13127_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6617 a_6619_23439# _0434_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6618 _0105_ a_18795_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6619 a_17118_9295# a_16679_9301# a_17033_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6623 a_14436_15529# cal_lut\[36\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X6624 a_14795_5162# _0301_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6625 vccd1 _0870_ a_25235_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6626 a_12334_17821# a_11895_17455# a_12249_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6627 vssd1 a_8146_18796# dbg_result[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X6628 a_4531_17705# _0741_ a_4313_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6629 _0839_ a_4167_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6630 a_26012_15939# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6631 vccd1 a_12042_3423# a_11969_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6632 a_7553_8751# a_7387_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6633 vssd1 a_15207_18543# _0483_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X6634 a_11425_13353# _0651_ a_11343_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6635 a_17857_24349# a_17323_23983# a_17762_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6636 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_1951_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X6637 a_5165_13103# _0204_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6638 vssd1 a_1641_28500# io_out[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6640 a_19618_2223# a_19303_2375# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6641 vccd1 a_26467_10205# a_26635_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6642 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6643 a_8951_25321# dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.41 ps=1.82 w=1 l=0.15
X6645 a_1753_26133# clknet_0_temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6646 vccd1 net29 a_12815_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6647 a_16727_4087# a_16823_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6650 _0021_ a_11987_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6651 vssd1 clknet_1_0__leaf_io_in[0] a_2143_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6652 a_2137_8751# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6653 vssd1 net10 a_7847_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6654 _0720_ dec1.i_ones vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6655 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4600_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X6656 net1 a_1407_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6657 vssd1 net34 a_25419_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6658 a_10252_13103# a_9853_13103# a_10126_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6659 vssd1 a_5693_21781# _0758_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6660 a_2511_21263# _0772_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X6661 a_8171_3476# _0314_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6662 vccd1 _0443_ a_20943_6369# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6669 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5823_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6671 a_9429_19605# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6672 vssd1 a_26203_6250# _0161_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6673 vccd1 net25 a_14839_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6675 a_22926_27221# a_22726_27521# a_23075_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6676 vccd1 a_1551_19605# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6677 vssd1 a_6979_19061# _0383_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6678 a_15469_12559# _0016_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6679 a_21997_11471# cal_lut\[157\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6681 _0262_ a_20907_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6682 a_18055_10383# a_17875_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6683 a_2741_24135# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6684 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6685 _0384_ _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6686 a_8951_13103# _0501_ a_9129_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X6687 vccd1 a_22235_16733# a_22403_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6688 vccd1 a_16079_3285# a_15903_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6689 _0594_ a_17507_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6690 vssd1 cal_lut\[38\] a_9037_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6691 vssd1 _0237_ a_25003_24833# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6693 vccd1 a_12723_21807# _0237_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6694 _0434_ net7 a_2489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X6695 a_4747_9117# a_3965_8751# a_4663_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6696 vssd1 a_4774_27765# a_4732_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6697 a_17401_24759# _0872_ a_17564_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6698 a_20924_19631# a_20525_19631# a_20798_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6699 a_6863_9117# a_6081_8751# a_6779_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6700 vccd1 net19 a_20943_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6701 dbg_result[5] a_11366_28588# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X6702 a_13257_23445# a_13091_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6703 a_5158_14735# a_4719_14741# a_5073_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6704 a_5284_6409# a_4885_6037# a_5158_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6705 net4 a_1407_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X6706 cal_lut\[115\] a_21759_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6708 net47 a_16219_25623# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6709 a_25047_16733# a_24867_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6710 a_16373_13077# _0596_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X6711 a_10501_13879# _0246_ a_10664_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6712 vccd1 a_15439_2388# _0179_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6713 a_20046_26677# a_19878_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6714 vssd1 a_8383_22583# _0777_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X6715 vssd1 cal_lut\[168\] a_25873_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6716 a_20756_12559# _0506_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6718 a_9235_25071# dec1.i_ones _0748_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.117 ps=1.01 w=0.65 l=0.15
X6719 a_6428_24501# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X6720 a_13990_26703# a_13717_26709# a_13905_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6721 a_4584_24759# _0798_ a_4726_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6722 vssd1 _0233_ a_22659_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6723 a_9117_14191# a_8951_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6724 a_12828_13103# a_12429_13103# a_12702_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6725 _0286_ a_16168_9411# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X6726 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6727 a_16168_9411# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6728 a_21591_4765# a_20893_4399# a_21334_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6729 a_9135_18319# _0519_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X6730 vssd1 a_12959_15253# _0275_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X6731 a_23549_8751# cal_lut\[165\] a_23477_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6732 vccd1 a_10108_4373# _0316_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6733 a_6000_31375# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X6734 vccd1 _0867_ a_21095_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6735 a_22997_4399# cal_lut\[152\] a_22925_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6736 a_9565_8751# cal_lut\[139\] a_9493_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6737 _0708_ a_10784_23983# a_11142_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6738 _0495_ a_13714_19407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X6739 vccd1 _0341_ a_23763_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6740 temp1.dac.vdac_single.en_pupd _0801_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6741 vccd1 a_20690_18517# _0452_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6742 temp1.capload\[11\].cap.Y net51 a_2505_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6743 a_3238_19881# _0421_ a_3154_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6744 vssd1 _0654_ a_12310_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6745 a_10585_16201# a_9595_15829# a_10459_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6747 vccd1 a_11579_25045# _0731_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X6748 vssd1 a_21334_25183# a_21292_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6750 a_13629_4943# _0118_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6752 vssd1 _0536_ a_20325_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6753 a_13487_25437# a_12705_25071# a_13403_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6754 a_6722_3677# a_6283_3311# a_6637_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6755 a_1551_19605# _0762_ a_1917_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6756 a_6480_29423# a_6081_29423# a_6354_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6757 a_12341_2223# _0147_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6758 vssd1 net8 a_10055_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6759 a_2489_17455# net7 _0434_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6760 dbg_result[0] a_7410_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X6762 _0051_ a_17415_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6763 vssd1 net22 a_2281_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6764 vccd1 _0361_ a_25051_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6765 a_2695_20969# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6766 vccd1 a_6879_6549# a_6703_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6767 vccd1 net38 a_24499_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6768 vccd1 a_8175_11445# _0881_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X6769 a_25271_25437# a_24573_25071# a_25014_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6770 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6771 a_21985_9661# cal_lut\[105\] a_21913_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6772 _0492_ _0464_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6773 vssd1 cal_lut\[5\] a_11895_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6774 vccd1 a_15623_15431# _0549_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6776 temp1.dac_vout_notouch_ net13 a_10488_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X6777 a_8533_22351# _0774_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X6778 vssd1 net42 a_24591_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6779 vssd1 a_13241_5633# _0569_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X6780 a_28031_15823# a_27167_15829# a_27774_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6781 cal_lut\[173\] a_28199_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6782 vccd1 _0713_ a_8055_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6783 _0707_ _0665_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6784 a_22806_25183# a_22638_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6786 a_24105_10357# _0510_ a_24262_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X6788 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd a_2879_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6790 a_24823_11079# a_24919_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6791 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6792 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_2327_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6793 a_21872_24643# _0260_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6794 cal_lut\[173\] a_28199_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6795 cal_lut\[82\] a_13571_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6798 a_2010_24759# _0415_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.151 ps=1.35 w=0.42 l=0.15
X6799 vccd1 a_25014_7093# a_24941_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6800 vccd1 _0464_ a_16187_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6801 a_19303_16519# _0459_ a_19537_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6802 vccd1 a_23351_7338# _0109_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6803 vssd1 net26 a_10607_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6804 a_18137_28879# _0051_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6805 _0523_ a_19623_23552# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6806 a_23117_4943# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X6807 vssd1 _0405_ a_7749_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6808 a_10235_8029# a_10055_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6809 a_10875_31849# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X6810 a_17244_9673# a_16845_9301# a_17118_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6811 a_25873_15101# a_25603_14735# a_25783_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X6812 a_4866_5599# a_4698_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6814 _0353_ a_27347_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6815 vccd1 a_14675_3829# a_14591_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6816 a_15299_12015# cal_lut\[192\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6817 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X6818 vssd1 _0484_ a_16300_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X6819 a_21173_14191# _0012_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6820 vccd1 cal_lut\[190\] a_14611_11079# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6821 a_8251_11293# a_7387_10927# a_7994_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6822 a_13863_12559# a_12999_12565# a_13606_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6825 vccd1 net10 a_7387_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6827 vccd1 a_5416_23413# _0821_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X6828 vccd1 net40 a_14655_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6829 a_5507_22325# _0788_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X6830 vssd1 a_21591_11293# a_21759_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6831 cal_lut\[53\] a_20471_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6832 vccd1 a_23450_7775# a_23377_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6833 vccd1 net29 a_15115_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6835 a_27149_7125# a_26983_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6836 a_3535_10761# a_3406_10505# a_3115_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6837 a_18489_28169# a_17935_28009# a_18142_28068# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6838 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_1775_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X6839 a_21725_16367# _0024_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6840 _0775_ _0724_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6841 a_20574_12559# _0537_ a_20325_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6842 a_18071_28169# a_17942_27913# a_17651_28023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6843 a_3990_24310# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X6844 a_19308_17973# _0507_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6845 vccd1 _0332_ a_14103_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6846 a_13533_12559# a_12999_12565# a_13438_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6848 a_22561_18793# _0643_ a_22465_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6850 a_13732_13967# _0487_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6852 a_22135_6941# a_21353_6575# a_22051_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6853 a_13349_9295# a_12815_9301# a_13254_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6855 vssd1 _0868_ a_23763_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6856 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6857 _0487_ a_16069_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X6858 vccd1 _0838_ a_2419_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6859 a_12672_30199# net8 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X6860 vccd1 _0240_ a_19531_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6862 _0300_ a_13040_6147# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6863 vssd1 _0422_ _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6864 a_20716_6351# cal_lut\[160\] a_20141_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X6865 _0284_ a_20952_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X6866 a_17743_2741# a_17919_3073# a_17871_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X6868 a_3882_22895# clknet_0_temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6869 _0581_ a_15667_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6870 vssd1 _0872_ a_15469_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6873 vccd1 cal_lut\[175\] a_22054_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6874 vccd1 a_5751_6005# a_5667_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6875 a_22009_11791# cal_lut\[103\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6876 _0865_ a_14696_14441# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6878 vccd1 a_13508_18517# a_13291_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.0672 ps=0.74 w=0.42 l=0.15
X6879 a_8837_5321# a_7847_4949# a_8711_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6880 vccd1 _0341_ a_24591_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6881 a_5809_10927# _0189_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6882 vccd1 cal_lut\[134\] a_5451_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6885 vccd1 a_14710_1247# a_14637_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6886 a_8372_31055# a_8123_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X6887 _0618_ a_18611_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6888 a_16845_9301# a_16679_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6890 a_4627_19631# _0738_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X6891 vssd1 a_18291_16532# _0077_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6892 vccd1 a_26283_8207# a_26451_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6893 vssd1 a_20747_7931# a_20705_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6895 a_1573_14741# a_1407_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6896 _0825_ a_1735_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6897 a_4885_14741# a_4719_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6899 vssd1 a_14123_23413# a_14081_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6900 a_23201_23145# _0469_ a_23055_23047# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6901 vssd1 net27 a_5455_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6902 vssd1 _0402_ a_5173_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6903 vssd1 a_9815_14557# a_9983_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6904 vccd1 a_6963_5853# a_7131_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6905 a_28115_12559# a_27333_12565# a_28031_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6907 vccd1 a_3155_16911# _0421_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X6910 vssd1 cal_lut\[104\] a_20952_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6911 a_9375_29397# ctr\[11\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6912 a_17946_26525# a_17673_26159# a_17861_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6914 _0826_ _0817_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6916 a_25962_11989# a_25762_12289# a_26111_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6918 a_15921_17455# a_14931_17455# a_15795_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6919 a_7147_3677# a_6283_3311# a_6890_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6920 a_17305_6575# a_17139_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6921 vccd1 cal_lut\[61\] a_23299_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6922 a_7323_12381# a_6541_12015# a_7239_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6923 a_15496_29257# a_15097_28885# a_15370_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6925 vssd1 a_19890_2197# a_19819_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6926 vssd1 _0679_ a_10233_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6927 vssd1 a_14967_1501# a_15135_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6928 _0160_ a_25879_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6929 _0226_ a_16859_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X6930 a_17661_5487# cal_lut\[131\] a_17589_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6932 vssd1 _0500_ a_9389_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X6933 vccd1 a_16255_25437# a_16423_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6934 _0233_ a_21872_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6935 a_12334_17821# a_12061_17455# a_12249_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6936 vccd1 net28 a_7387_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6937 a_9765_6727# _0299_ a_9928_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6938 vssd1 _0523_ a_19681_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6940 a_9947_26703# ctr\[6\] a_9835_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.131 ps=1.05 w=0.64 l=0.15
X6941 a_2249_24887# _0415_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.13 ps=1.11 w=0.42 l=0.15
X6942 _0730_ _0711_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6943 vccd1 cal_lut\[113\] a_18515_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6944 a_4187_28918# _0801_ a_4187_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6945 vccd1 net31 a_20727_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6946 _0310_ a_10280_5059# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X6947 vccd1 _0472_ a_16771_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6948 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9568_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X6949 vssd1 a_6611_22583# _0788_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X6951 vccd1 net23 a_6743_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6952 a_2121_23983# net22 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.101 ps=0.96 w=0.65 l=0.15
X6953 a_12827_10927# a_12691_10901# a_12407_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6954 a_7840_28585# _0405_ _0210_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X6955 vssd1 _0838_ a_3325_8903# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6956 a_2485_22671# net22 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6957 a_19705_23805# _0459_ a_19623_23552# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6958 _0613_ a_16574_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X6959 a_6848_3311# a_6449_3311# a_6722_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6961 vssd1 io_in[0] a_6458_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6962 a_13052_15797# _0518_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6963 _0363_ a_11579_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6964 vssd1 net25 a_13643_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6965 vssd1 cal_lut\[98\] a_11981_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6966 vssd1 cal_lut\[61\] a_22937_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6968 a_15002_21263# a_14729_21269# a_14917_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6970 vccd1 _0856_ a_23671_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6971 _0451_ a_22843_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6973 a_12337_3861# a_12171_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6974 a_6909_7119# a_6375_7125# a_6814_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6975 vccd1 a_11794_8725# a_11723_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X6976 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_4811_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6978 cal_lut\[64\] a_27371_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6980 vccd1 a_10924_31751# a_10875_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X6981 vssd1 a_12318_26677# a_12276_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6982 dbg_result[4] a_11458_27500# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X6983 _0382_ _0447_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6984 a_8723_17130# _0842_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6985 a_18114_26271# a_17946_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6986 vssd1 a_19383_16911# a_19551_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6987 _0655_ a_12162_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X6988 vccd1 a_23139_13371# a_23055_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6990 _0418_ a_2327_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6992 cal_lut\[172\] a_28199_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6993 a_2605_21263# _0770_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6994 vssd1 net41 a_14563_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6995 a_20779_15253# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6996 _0365_ a_15479_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X6997 a_11881_7119# _0123_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6998 a_4283_22057# _0758_ a_4477_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X6999 vssd1 _0467_ a_9988_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X7000 a_5081_19881# _0429_ _0739_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7001 vssd1 net18 a_22961_17249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7002 a_12679_28010# _0847_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7005 vssd1 a_22695_8207# a_22863_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7006 cal_lut\[172\] a_28199_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7008 vccd1 a_15991_8903# _0548_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7009 vssd1 a_7987_9514# _0120_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7010 _0714_ _0706_ a_11547_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7011 a_17217_17999# _0076_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7012 a_13904_13647# _0515_ a_13649_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X7014 vccd1 a_11671_2741# _0331_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X7015 _0246_ a_24407_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7017 a_2060_30199# _0833_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X7018 a_12575_26703# a_11877_26709# a_12318_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7019 vccd1 _0438_ a_13275_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7020 a_4425_5487# a_4259_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7021 cal_lut\[36\] a_14675_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7022 a_22431_7338# _0343_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7024 vssd1 a_5307_29789# a_5475_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7025 vccd1 a_9155_14709# a_9071_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7026 vccd1 a_13606_12533# a_13533_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7028 a_25014_25183# a_24846_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7029 vssd1 net43 a_26339_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7030 vccd1 net41 a_13643_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7032 vssd1 _0707_ a_11142_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7033 cal_lut\[3\] a_8971_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7034 a_11471_14557# a_10607_14191# a_11214_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7035 vccd1 _0803_ a_3418_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X7036 cal_lut\[86\] a_23231_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7038 vssd1 cal_lut\[163\] a_24125_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7039 dbg_result[4] a_11458_27500# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7040 vccd1 _0098_ a_12141_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7041 a_8297_20765# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7042 vccd1 _0474_ a_18369_18337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7043 a_19609_5487# _0113_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7044 vssd1 clknet_1_0__leaf__0380_ a_5377_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7045 _0477_ a_13751_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7047 vccd1 _0216_ a_22567_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7048 a_18475_18695# _0454_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7049 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7050 a_17871_9117# a_17691_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7051 _0105_ a_18795_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7052 a_6445_29111# a_6541_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X7053 vccd1 a_3299_19061# _0745_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7054 vccd1 a_14103_17455# _0447_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7055 vccd1 a_14507_15823# a_14675_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7056 vccd1 net40 a_12539_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7057 _0192_ _0381_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7058 a_25858_8207# a_25585_8213# a_25773_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7059 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8372_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X7060 _0757_ _0737_ a_3974_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X7061 a_10413_20969# _0677_ a_10331_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7062 vccd1 a_17727_17999# a_17895_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7063 a_11141_14557# a_10607_14191# a_11046_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7064 vccd1 a_8803_1679# a_8971_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7065 a_17475_16041# net44 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7066 a_17727_2589# a_16863_2223# a_17470_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7068 a_7826_13469# a_7387_13103# a_7741_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7069 a_8845_28023# dec1.i_ones vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X7070 vssd1 a_2564_25045# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7071 vssd1 a_14139_28879# a_14307_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7072 a_26505_18909# a_25971_18543# a_26410_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7073 vssd1 a_19402_25589# a_19360_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7074 vssd1 a_9275_15444# _0079_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7075 vssd1 cal_lut\[150\] a_19065_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7077 a_24573_23983# a_24407_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7079 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7081 a_4310_8439# a_4406_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7082 cal_lut\[163\] a_28015_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7083 a_1861_8751# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7084 a_24573_22895# a_24407_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7086 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7087 vccd1 a_20671_22351# a_20839_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7088 _0806_ _0805_ a_3339_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7089 a_11527_12559# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7090 a_7952_16367# a_7553_16367# a_7826_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7091 a_15879_17821# a_15097_17455# a_15795_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7092 _0593_ a_16771_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7093 vssd1 net45 a_20727_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7094 vccd1 _0681_ a_10607_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7095 a_23915_17129# net42 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7096 a_17888_23983# a_17489_23983# a_17762_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7097 vccd1 a_5141_21781# _0756_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7098 a_13275_20175# _0447_ a_13525_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7099 vccd1 _0467_ a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X7100 a_3351_27569# net70 a_2839_27221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X7103 io_out[4] a_1464_23957# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X7104 vccd1 a_13459_4399# _0283_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7105 temp1.dac_vout_notouch_ net13 a_11868_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X7107 vssd1 a_12219_17130# _0005_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7109 vssd1 net11 a_9319_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
R18 temp1.capload\[14\].cap_54.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7110 a_18821_10749# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7111 vccd1 _0720_ a_11317_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7112 a_12693_6397# cal_lut\[130\] a_12621_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7113 vssd1 _0338_ a_19439_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7114 a_8478_19631# _0764_ a_8392_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X7115 a_15281_3861# a_15115_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7116 a_16907_1985# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7117 vccd1 _0836_ a_7111_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7118 a_26891_11293# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7119 vccd1 net27 a_5455_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7120 a_23351_8439# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7121 a_2503_31055# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X7123 vssd1 a_6428_24501# _0793_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X7124 a_28115_11471# a_27333_11477# a_28031_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7125 a_8390_23439# clknet_0__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7126 a_24726_9839# cal_lut\[164\] a_24636_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X7127 a_23758_20541# a_23443_20407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7128 a_4974_8029# a_4535_7663# a_4889_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7129 a_9005_24501# _0727_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X7130 a_15327_5853# a_14545_5487# a_15243_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7131 vccd1 a_13219_27613# a_13387_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7132 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X7133 _0254_ a_17456_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X7135 _0474_ a_13291_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7136 vccd1 _0247_ a_26063_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7137 vccd1 _0446_ a_11199_17607# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.118 ps=1.4 w=0.42 l=0.15
X7138 vccd1 a_8251_6941# a_8419_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7139 vccd1 cal_lut\[162\] a_20112_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7140 a_25313_23439# _0062_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7141 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7143 vssd1 a_13035_3855# a_13203_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7144 vssd1 a_22633_11445# _0457_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X7145 a_12441_12015# a_12171_12381# a_12351_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X7146 vccd1 _0420_ a_4443_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7147 a_5341_17429# clknet_0_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7148 a_10402_3677# a_9963_3311# a_10317_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7149 vssd1 a_6890_3423# a_6848_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7150 a_11693_7125# a_11527_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7153 a_10832_16617# _0519_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7155 a_26107_8725# _0341_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7156 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7157 vssd1 _0500_ a_9297_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X7158 a_20433_27797# a_20267_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7159 vssd1 cal_lut\[167\] a_27437_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7162 vssd1 cal_lut\[33\] a_24861_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7163 a_22461_13103# _0013_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7164 vssd1 a_15262_23413# a_15220_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7165 a_6982_17973# a_6823_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X7168 a_20706_27791# a_20433_27797# a_20621_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7169 a_27701_17821# a_27167_17455# a_27606_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7170 vccd1 a_15795_28879# a_15963_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7171 _0848_ a_12995_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X7172 vccd1 a_13691_28500# _0049_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R19 vssd1 net64 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7175 a_14507_15823# a_13643_15829# a_14250_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7176 a_17739_7815# a_17835_7637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7177 a_10689_24893# _0681_ a_10607_24640# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7178 net11 a_8543_30485# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7179 vssd1 a_14703_25236# _0093_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7180 a_7182_6031# a_6909_6037# a_7097_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7181 vssd1 net29 a_9687_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7182 vssd1 _0413_ a_2419_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X7183 _0384_ clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7185 a_19789_24527# a_19255_24533# a_19694_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7186 vccd1 a_14163_8903# _0493_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7187 a_17066_13647# _0598_ a_16986_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7188 vssd1 a_6963_5853# a_7131_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7189 vssd1 a_16731_9813# net38 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X7190 vccd1 a_14611_11079# _0563_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7191 vccd1 a_22695_23439# a_22863_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7193 a_19399_2197# a_19683_2197# a_19618_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X7194 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7196 vssd1 net35 a_15943_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7198 vccd1 _0720_ a_6277_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X7199 vssd1 a_22695_23439# a_22863_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7202 vssd1 a_17401_24759# _0215_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X7203 vccd1 _0465_ a_17999_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7204 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7205 a_14177_15823# a_13643_15829# a_14082_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7206 vssd1 _0240_ a_19531_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7207 a_22431_13866# _0855_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7208 a_21897_12533# _0476_ a_22150_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X7209 vccd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7210 a_19333_25223# cal_lut\[47\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X7211 vccd1 _0744_ a_2247_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X7213 vssd1 net10 a_8123_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X7214 vssd1 a_13969_18218# net16 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7215 a_11214_14303# a_11046_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7216 vssd1 a_10501_13879# _0257_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X7217 vccd1 ctr\[1\] a_4744_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7218 a_8378_1679# a_8105_1685# a_8293_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7219 a_7323_12559# a_6541_12565# a_7239_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7221 _0850_ a_10699_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7222 _0308_ a_7980_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X7223 vssd1 a_15595_10357# a_15553_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7224 a_6699_13268# _0860_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7225 _0438_ a_13459_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X7226 a_23719_4087# a_23815_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7227 a_15991_8903# _0514_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7229 a_7011_31849# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X7230 vccd1 a_11214_14303# a_11141_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7231 a_12355_4765# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7232 vssd1 cal_lut\[112\] a_16996_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7233 a_6449_9117# a_5915_8751# a_6354_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7234 a_6647_28585# _0404_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7235 a_10045_9295# _0693_ a_9963_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7236 vccd1 net43 a_26339_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7237 vccd1 _0266_ a_12079_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7238 a_24846_24349# a_24407_23983# a_24761_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7239 vssd1 a_6375_19095# _0432_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X7240 vccd1 a_17159_22075# a_17075_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7241 vccd1 a_26578_18655# a_26505_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7242 a_20579_8029# a_19715_7663# a_20322_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7243 vccd1 a_5323_4917# _0319_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X7244 a_23631_11079# _0511_ a_23959_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7245 _0776_ _0728_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7246 _0433_ a_8544_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7247 a_17095_10004# _0286_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7248 a_10521_21263# _0591_ a_10715_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7249 vssd1 a_6503_16733# a_6674_16620# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7250 a_26330_14165# a_26130_14465# a_26479_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7251 _0658_ a_23395_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7253 _0693_ a_9411_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7255 vccd1 _0418_ a_3991_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7256 _0295_ a_20676_5059# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X7257 a_20119_24527# a_19421_24533# a_19862_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7258 a_6645_20719# _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X7259 a_22273_13103# a_22107_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7260 vccd1 _0331_ a_11711_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7261 vssd1 a_12134_7093# a_12092_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7262 a_27973_18377# a_26983_18005# a_27847_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7263 a_19111_19407# a_19057_19319# a_19011_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X7264 vssd1 a_10827_7119# a_10995_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7265 _0814_ a_5915_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7266 vccd1 temp1.dac.vdac_single.en_pupd a_3247_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X7267 a_1551_19605# _0428_ a_2107_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7270 a_19694_5853# a_19255_5487# a_19609_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7271 a_15630_19743# a_15462_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7272 a_4816_16617# ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7273 vccd1 a_12099_15547# a_12015_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7274 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X7275 vssd1 _0781_ a_4169_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X7276 vccd1 a_2552_31287# a_2503_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X7277 _0415_ clknet_1_1__leaf_io_in[0] a_1867_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7278 vssd1 a_15887_19997# a_16055_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7279 a_17536_10383# _0449_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7280 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_10239_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7281 vssd1 _0784_ a_3850_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7282 a_22523_5175# _0451_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7284 a_16293_21807# a_16127_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7285 a_2614_19631# _0761_ a_1551_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.0878 ps=0.92 w=0.65 l=0.15
X7286 vccd1 _0628_ _0668_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X7287 _0146_ a_9963_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7289 a_8971_22895# _0712_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X7290 a_11200_29575# net8 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X7291 vccd1 a_17930_25183# a_17857_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7292 vssd1 net40 a_14011_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7293 a_2125_15829# a_1959_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7296 a_2931_17455# _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7297 vccd1 a_7315_3579# a_7231_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7299 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7380_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X7300 a_21879_16055# _0505_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7301 a_10385_23413# _0680_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X7303 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6459_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X7304 a_4719_20495# _0747_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X7305 vssd1 a_26267_17723# a_26225_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7307 _0043_ a_17047_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7308 _0754_ a_2417_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7310 vccd1 a_7239_14735# a_7410_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X7311 vccd1 a_23211_6575# net33 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7312 vssd1 _0469_ a_19244_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X7313 vccd1 cal_lut\[58\] a_21954_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7314 a_6890_3423# a_6722_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7316 vccd1 cal_lut\[1\] a_6647_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7317 vssd1 _0419_ a_3435_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7318 vccd1 _0433_ _0662_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X7320 _0166_ a_26615_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7321 a_15439_17130# _0274_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7323 a_12518_1679# a_12245_1685# a_12433_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7324 dbg_result[5] a_11366_28588# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X7326 a_20203_4765# a_19421_4399# a_20119_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7327 a_20867_2986# _0337_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7328 a_18107_8439# net19 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7330 vccd1 clknet_0_io_in[0] a_6182_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7331 vccd1 a_27774_17567# a_27701_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7332 vssd1 a_17930_1653# a_17888_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7334 vssd1 _0424_ a_3067_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7335 vccd1 net26 a_9595_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7336 a_10528_3311# a_10129_3311# a_10402_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7337 vccd1 _0441_ a_20175_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7338 vssd1 a_12863_14954# _0096_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7339 a_17727_2589# a_17029_2223# a_17470_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7340 a_23009_7663# a_22843_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7341 a_8251_11293# a_7553_10927# a_7994_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7342 a_10911_1679# a_10129_1685# a_10827_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7343 vssd1 _0201_ a_3953_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7344 a_13345_27247# a_12355_27247# a_13219_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7345 vssd1 net67 a_3882_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7346 a_18041_12565# a_17875_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7347 vccd1 a_7159_11092# _0187_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7348 vccd1 ctr\[1\] a_2939_23047# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7349 vssd1 _0453_ a_19439_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X7350 _0650_ a_11527_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7351 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X7352 vssd1 _0422_ _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X7353 a_5073_14735# _0205_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7355 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7356 a_7102_21807# _0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7359 a_2397_15113# a_1407_14741# a_2271_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7360 vssd1 _0173_ a_28149_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7361 vssd1 a_10197_25223# _0733_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7362 vssd1 a_8695_3829# a_8653_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7363 net26 a_10659_7637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7364 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X7365 vssd1 a_6982_17973# a_6920_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X7366 vssd1 a_5326_14709# a_5284_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7367 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7368 vssd1 _0477_ a_16189_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7370 net73 a_7475_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7371 vssd1 a_13459_17455# _0438_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7372 a_13183_24349# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7373 a_2099_18695# a_2371_18523# a_2329_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7374 a_11966_7119# a_11527_7125# a_11881_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7375 a_12259_9295# a_12079_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7376 vssd1 a_3877_11703# _0396_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X7377 _0766_ a_8478_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7378 vccd1 a_14345_9269# _0565_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X7379 vccd1 a_15370_19407# _0467_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7380 vccd1 cal_lut\[155\] a_18015_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X7382 a_5801_9673# a_4811_9301# a_5675_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7384 a_21223_19997# a_20359_19631# a_20966_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7386 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7387 a_7994_8863# a_7826_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7388 a_20775_27412# _0228_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7390 vssd1 _0538_ _0539_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X7391 cal_lut\[20\] a_8419_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7392 _0326_ a_6187_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X7393 vccd1 _0390_ a_4705_27552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7394 vssd1 a_9375_29397# a_9117_29397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X7396 a_15972_10089# _0492_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7397 vssd1 a_24105_10357# _0695_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X7398 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X7399 _0381_ clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7401 a_27163_9295# a_26983_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7402 vccd1 _0459_ a_20451_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7403 a_26233_16367# _0072_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7406 vccd1 a_11366_28588# a_11279_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X7408 a_23565_19087# _0026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7409 vccd1 net23 a_7847_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7410 a_25957_9839# _0169_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7411 vccd1 net35 a_15943_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7413 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4435_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X7414 a_13127_13469# a_12263_13103# a_12870_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7415 a_14457_7663# _0124_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7417 a_17354_10383# _0623_ a_17105_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7419 _0697_ a_8758_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X7420 vssd1 a_28031_15823# a_28199_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7421 cal_lut\[108\] a_20747_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7422 dbg_result[2] a_8146_18796# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X7423 vccd1 cal_lut\[112\] a_17078_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7424 a_22813_8751# cal_lut\[153\] a_22741_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7425 a_9358_3855# _0476_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X7426 cal_lut\[162\] a_26819_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7428 vssd1 a_17739_21959# _0553_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X7429 a_17841_12161# _0605_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7431 _0155_ a_17415_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7432 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X7433 a_15553_10761# a_14563_10389# a_15427_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7434 vssd1 _0784_ a_4408_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X7435 vccd1 _0692_ a_9873_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.117 ps=1.24 w=1 l=0.15
X7436 a_3007_14557# a_2143_14191# a_2750_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7437 a_13570_5737# _0567_ a_13490_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7438 vccd1 net34 a_17783_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7439 a_27351_13469# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7440 _0519_ a_13052_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7441 a_4931_24135# _0797_ a_5077_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7442 vssd1 clknet_1_0__leaf_io_in[0] a_7111_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7443 a_21794_6687# a_21626_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7445 vccd1 cal_lut\[77\] a_17996_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7446 a_5399_8029# a_4701_7663# a_5142_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7447 vccd1 _0305_ a_11527_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7448 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7449 _0033_ a_25235_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7450 a_22633_18793# _0639_ a_22561_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7451 vccd1 a_17895_2491# a_17811_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7452 vssd1 _0266_ a_13135_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7453 a_7994_13215# a_7826_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7454 a_10746_10615# _0515_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X7455 a_10137_22895# _0680_ _0682_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7456 a_21794_6687# a_21626_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7457 vccd1 a_25439_25339# a_25355_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7458 a_19878_26703# a_19605_26709# a_19793_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7459 vccd1 dbg_result[1] a_19057_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X7461 a_3848_27399# _0829_ a_3990_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7462 a_17628_19881# _0468_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7464 a_14773_10927# _0483_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7465 vccd1 a_7072_15797# net41 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7466 a_2677_14557# a_2143_14191# a_2582_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7467 cal_lut\[164\] a_25439_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7468 vssd1 a_22903_2985# a_22910_2889# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7469 a_17305_6575# a_17139_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7470 _0625_ a_16373_16341# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.91 w=0.65 l=0.15
X7471 a_8293_15823# _0002_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7472 vccd1 _0242_ a_21739_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7473 a_18003_6941# a_17139_6575# a_17746_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7474 a_19820_5487# a_19421_5487# a_19694_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7475 a_21157_8573# cal_lut\[111\] a_21085_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7476 a_5336_31849# a_5087_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X7477 io_out[1] a_1551_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7478 vccd1 _0722_ a_7289_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7479 a_6062_11039# a_5894_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7480 vssd1 a_24306_12836# a_24235_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7481 vccd1 a_5227_26935# _0812_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7482 vccd1 a_21591_4765# a_21759_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7483 a_14542_8029# a_14103_7663# a_14457_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7484 vssd1 _0424_ a_3062_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X7485 a_22235_16733# a_21537_16367# a_21978_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7486 a_13069_2057# a_12079_1685# a_12943_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7487 vccd1 a_3799_19631# _0737_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7488 a_22654_27247# a_22339_27399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7489 _0034_ a_14747_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7491 a_22874_17999# _0642_ a_22625_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7492 a_9779_11177# _0512_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X7493 _0066_ a_21739_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7494 a_22619_2999# a_22910_2889# a_22861_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7495 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7496 a_5460_15823# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7497 a_24351_14735# a_23487_14741# a_24094_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7498 a_24455_19783# a_24551_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7499 _0253_ a_17135_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X7500 a_18090_12265# _0607_ a_17841_12161# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7501 vssd1 a_2695_14013# _0808_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X7502 a_7921_13469# a_7387_13103# a_7826_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7503 vccd1 a_9547_3073# a_9371_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X7504 vccd1 _0438_ a_13551_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X7505 a_16293_21807# a_16127_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7506 vssd1 cal_lut\[8\] a_13085_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7508 a_16508_10927# a_16109_10927# a_16382_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7509 a_7553_16367# a_7387_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7510 a_15623_15431# _0531_ a_15857_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7511 vccd1 cal_lut\[114\] a_20756_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7513 a_17555_28023# a_17651_28023# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7515 _0357_ a_27163_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X7516 a_22625_17973# _0640_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7517 a_15094_29789# a_14821_29423# a_15009_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7518 vssd1 cal_lut\[123\] a_11337_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7519 vccd1 dbg_result[4] _0453_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7520 vssd1 _0491_ a_15193_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7521 vccd1 a_7410_17973# a_7323_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X7522 a_1857_21365# clknet_1_1__leaf_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7523 vccd1 a_15903_3285# _0366_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X7525 vssd1 a_5751_6005# a_5709_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7526 vssd1 _0836_ a_12525_18231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7527 vssd1 _0290_ a_14699_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7528 vssd1 _0422_ a_2371_18523# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7529 vssd1 a_19303_18695# _0507_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7530 vssd1 a_10570_3423# a_10528_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7531 _0421_ a_3155_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7532 a_4903_11293# _0836_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7533 a_21913_11471# _0683_ a_21831_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7534 a_26307_13077# net37 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7535 vccd1 _0216_ a_16679_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7536 vssd1 a_25014_23007# a_24972_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7537 vccd1 _0492_ a_10129_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7538 _0390_ a_2419_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7539 a_20245_15279# a_19255_15279# a_20119_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7541 a_8297_20175# _0434_ _0435_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7543 a_19777_23805# cal_lut\[48\] a_19705_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7544 vssd1 a_1458_30199# a_1407_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7545 cal_lut\[180\] a_15871_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7547 a_22113_16189# cal_lut\[168\] a_22041_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7548 vssd1 a_10719_13371# a_10677_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7549 a_13291_18909# a_13091_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X7550 a_1917_19881# _0761_ a_1551_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7551 vccd1 _0442_ a_21555_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7553 a_18077_8029# a_17739_7815# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7555 _0258_ a_12120_14851# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X7556 vssd1 a_25007_5175# cal_lut\[161\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7557 _0644_ a_15023_22464# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7558 a_6979_19061# ctr\[4\] a_7206_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X7559 vccd1 net42 a_23211_19093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7560 vccd1 a_7350_6005# a_7277_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7561 vccd1 a_13367_10391# _0260_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7562 _0391_ a_2071_11791# a_2309_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X7563 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7564 vccd1 io_in[2] a_1407_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7565 _0646_ a_14287_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7566 a_11900_22351# _0679_ _0710_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X7567 a_26265_13469# a_25927_13255# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7568 a_20855_16911# a_19991_16917# a_20598_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7569 a_6637_3311# _0133_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7570 a_2750_20407# _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X7571 vssd1 _0490_ _0517_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7574 a_18773_29257# a_17783_28885# a_18647_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7575 vccd1 a_26835_18909# a_27003_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7577 _0456_ a_18597_13077# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X7578 a_6458_20175# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7579 a_25218_13469# a_24971_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7580 a_15711_24833# _0266_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7583 a_10304_29967# a_10055_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X7585 a_9836_23145# _0716_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X7586 a_17446_19881# _0581_ a_17197_19777# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7587 vccd1 a_19057_26935# _0227_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X7588 _0303_ a_8164_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X7589 a_17168_12559# _0601_ a_17066_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X7590 vccd1 _0446_ a_13459_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.109 ps=1.36 w=0.42 l=0.15
X7591 a_21085_11471# _0449_ a_21169_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7592 a_1736_18517# _0743_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X7593 a_16156_15823# _0484_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7594 net76 a_6739_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7595 _0164_ a_24039_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7596 a_25953_8207# a_25419_8213# a_25858_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7597 _0632_ a_22291_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7598 a_13085_26159# a_12815_26525# a_12995_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X7600 vccd1 a_8546_1653# a_8473_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7601 vccd1 a_5971_15253# a_5713_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X7602 vccd1 net15 a_12455_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7603 a_24469_17289# a_23922_17033# a_24122_17188# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7604 a_21166_4765# a_20727_4399# a_21081_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7606 a_25927_13255# a_26023_13077# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7607 vssd1 a_13415_20884# _0039_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7608 a_2750_14303# a_2582_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7610 a_17555_28023# a_17651_28023# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7611 a_19763_28010# _0223_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7612 a_3241_21583# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7614 a_3112_19783# _0420_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7615 vccd1 a_20747_7931# a_20663_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7616 a_22546_13469# a_22273_13103# a_22461_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7617 a_25014_24095# a_24846_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7618 a_27590_17973# a_27422_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7619 vssd1 _0245_ a_25327_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7620 a_12672_30199# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7621 a_8730_14709# a_8562_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7623 a_6624_31055# a_6375_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X7624 a_25891_20553# a_25755_20393# a_25471_20407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7625 a_15979_3855# a_15115_3861# a_15722_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7626 cal_lut\[190\] a_6487_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7627 a_27438_15279# a_27123_15431# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7628 a_13472_21641# a_13073_21269# a_13346_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7629 vccd1 a_24122_17188# a_24051_17289# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7630 vssd1 net39 a_17415_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X7631 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_5336_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X7632 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7633 _0268_ a_18560_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X7634 a_25907_23439# a_25125_23445# a_25823_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7635 vccd1 cal_lut\[177\] a_16859_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7636 a_6427_11445# a_6603_11777# a_6555_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X7637 vssd1 _0648_ _0661_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.0878 ps=0.92 w=0.65 l=0.15
X7638 vssd1 dbg_result[3] a_14655_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7639 vssd1 a_6947_29691# a_6905_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7640 a_3246_25321# _0803_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X7641 _0216_ a_13459_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X7642 vssd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7643 a_15645_28169# a_14655_27797# a_15519_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7645 a_8562_14735# a_8289_14741# a_8477_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7646 vssd1 a_18519_21263# _0454_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7647 vssd1 a_7994_6687# a_7952_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7648 a_5818_27247# a_5503_27399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7649 vccd1 _0462_ a_22659_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7650 a_6732_28335# _0403_ a_6429_28309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X7652 a_20797_22729# a_19807_22357# a_20671_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7653 a_22553_25071# _0085_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7654 a_20525_19631# a_20359_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7655 a_14668_7663# a_14269_7663# a_14542_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7656 a_2695_14013# ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X7657 vccd1 a_7994_13215# a_7921_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7658 cal_lut\[159\] a_23323_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7659 vssd1 a_15722_3829# a_15680_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7660 _0876_ a_24679_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X7661 _0054_ a_21463_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7662 a_12705_25071# a_12539_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7663 _0390_ a_2419_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7664 vssd1 net10 a_10239_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X7665 vccd1 a_3155_16911# _0421_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7666 vssd1 _0452_ a_16281_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7668 a_18555_3677# a_17691_3311# a_18298_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7670 a_17845_29423# a_17291_29397# a_17498_29397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7671 a_5143_11445# ctr\[4\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7672 vccd1 _0495_ a_16955_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7673 a_27057_8751# a_26891_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7674 vccd1 clknet_1_0__leaf_io_in[0] a_1407_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7675 a_11707_12559# a_11527_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7676 a_20119_11293# a_19421_10927# a_19862_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7677 a_12429_13103# a_12263_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7678 cal_lut\[162\] a_26819_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7679 a_4153_9839# _0000_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7680 a_18893_10749# cal_lut\[167\] a_18821_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7681 _0774_ a_7939_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7682 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7683 net68 clknet_1_0__leaf_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7684 a_22259_19605# net43 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7685 a_7718_18679# a_7559_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X7686 a_20775_14967# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7687 vccd1 net23 a_6283_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7688 a_15051_1501# a_14269_1135# a_14967_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7689 a_22730_6031# a_22291_6037# a_22645_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7690 vccd1 _0290_ a_19439_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7691 a_10844_31029# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7692 a_5013_24825# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X7693 vssd1 _0238_ a_24683_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7694 a_25106_15797# a_24938_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7695 a_14795_5162# _0301_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7696 a_20943_6369# _0441_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7697 vccd1 _0635_ a_22633_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7699 vccd1 a_12686_1653# a_12613_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7700 a_14195_28701# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7701 a_22887_6549# _0341_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7702 a_25690_12015# a_25375_12167# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7703 a_16255_25437# a_15557_25071# a_15998_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7704 vccd1 _0176_ a_25757_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7705 a_10229_24233# _0682_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X7706 a_16731_9813# net39 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X7707 vssd1 ctr\[2\] a_2972_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X7708 a_26651_6941# a_25953_6575# a_26394_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7709 _0703_ a_9749_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7710 vssd1 _0851_ a_15193_14343# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7711 a_5825_17999# _0839_ _0195_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7712 vccd1 _0808_ _0393_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7713 a_6081_29423# a_5915_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7714 a_10025_29257# a_9471_29097# a_9678_29156# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7715 a_24551_19605# a_24835_19605# a_24770_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X7716 a_22217_19997# a_21879_19783# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7717 _0282_ a_20032_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X7718 a_12075_18793# net15 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7719 vccd1 a_5278_12533# net72 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.273 pd=1.61 as=0.495 ps=2.99 w=1 l=0.15
X7720 a_25589_17455# _0069_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7721 a_9022_8207# a_8749_8213# a_8937_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7723 vssd1 a_7111_17455# _0437_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7724 a_6909_6037# a_6743_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7725 a_11247_6941# a_11067_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7727 a_6555_11837# cal_lut\[190\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X7729 vssd1 _0576_ a_11950_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X7730 _0166_ a_26615_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7731 vssd1 a_16179_29397# _0218_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X7732 a_7465_14191# _0036_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7734 a_10924_31751# net65 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X7736 temp1.dac_vout_notouch_ net13 a_10304_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X7737 a_15220_28169# a_14821_27797# a_15094_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7738 a_5998_21583# _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X7739 a_5418_13215# a_5250_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7740 a_17677_1679# _0185_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7741 a_11981_9839# a_11711_10205# a_11891_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X7742 a_21810_22173# a_21371_21807# a_21725_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7744 a_25375_20407# a_25471_20407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7745 a_10041_11471# _0038_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7746 a_8473_1679# a_7939_1685# a_8378_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7747 vccd1 a_8711_4943# a_8879_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7748 vccd1 net9 a_11619_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X7749 a_5081_19881# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X7750 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7752 vccd1 a_23631_11079# _0512_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X7753 vssd1 a_7159_11092# _0187_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7755 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7757 a_22441_21237# _0638_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X7758 vssd1 clknet_1_0__leaf__0380_ _0382_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7759 vccd1 _0341_ a_20635_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X7760 vssd1 _0492_ a_14920_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X7762 a_2060_30199# _0833_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7763 a_7013_26159# _0811_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7764 a_22488_15113# a_22089_14741# a_22362_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7765 vccd1 a_3155_9839# _0836_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7766 vccd1 _0417_ a_2327_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7767 vccd1 a_14523_6549# _0307_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X7768 a_2149_28585# _0817_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7769 a_1736_18517# _0743_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7770 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_1867_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X7773 _0371_ a_13823_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X7774 a_12079_7663# cal_lut\[142\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7775 vssd1 a_17197_19777# _0582_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7776 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6624_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X7777 a_21879_19783# a_21975_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7778 vssd1 a_16737_13621# _0600_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7779 a_17739_7815# a_17835_7637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7780 a_18751_23671# _0481_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7781 a_21292_4399# a_20893_4399# a_21166_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7782 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7783 a_7826_29789# a_7553_29423# a_7741_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7784 a_15519_23439# a_14821_23445# a_15262_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7785 _0481_ a_12263_20495# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.213 ps=1.3 w=0.65 l=0.15
X7786 vssd1 a_14507_15823# a_14675_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7789 a_9043_11177# cal_lut\[188\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X7790 a_19694_4765# a_19421_4399# a_19609_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7791 vssd1 cal_lut\[157\] a_20905_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7792 vssd1 _0463_ a_22729_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7793 a_7165_23983# _0722_ _0752_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7794 a_11149_19087# _0589_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7795 vssd1 net28 a_8123_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7797 a_1941_12559# a_1407_12565# a_1846_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7798 a_13751_16911# _0425_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X7799 vssd1 a_6982_12533# a_6940_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7802 vccd1 a_5324_4373# net23 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7803 vssd1 a_22983_15431# _0537_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X7804 a_27973_7497# a_26983_7125# a_27847_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7805 vssd1 _0870_ a_25235_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7806 a_16035_18112# cal_lut\[95\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7807 vccd1 a_28015_17973# a_27931_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7809 vssd1 a_2564_25045# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7810 vccd1 cal_lut\[59\] a_18475_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X7811 a_12065_26703# _0006_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7812 vccd1 _0444_ a_21169_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7813 a_21258_14557# a_20819_14191# a_21173_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7814 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7816 vssd1 a_22863_1653# a_22821_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7817 a_24033_6397# a_23763_6031# a_23943_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X7818 cal_lut\[157\] a_21115_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7819 a_22445_7663# cal_lut\[159\] a_22373_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7820 a_25927_10602# _0355_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7821 a_19609_10927# _0102_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7822 a_5039_25071# ctr\[7\] a_4676_25223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7823 _0874_ a_20860_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X7824 a_8171_3476# _0314_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7825 vccd1 net79 a_5353_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7826 a_11287_27613# a_10589_27247# a_11030_27383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X7827 a_22435_27221# a_22726_27521# a_22677_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7828 vssd1 _0447_ _0472_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7829 vssd1 a_10995_7093# a_10953_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7830 a_19619_7119# a_19439_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7831 vccd1 a_17475_16041# a_17482_15945# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7832 vssd1 a_2439_14709# a_2397_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7833 vssd1 a_3175_14459# a_3133_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7834 vccd1 net11 a_9779_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X7835 vccd1 net47 a_24407_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7836 vssd1 a_7350_6005# a_7308_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7837 a_13341_9001# _0565_ a_13269_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7838 a_12525_3855# _0130_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7839 vssd1 a_14710_7775# a_14668_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7840 vssd1 net35 a_19255_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7841 vssd1 net47 a_24407_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7842 vssd1 cal_lut\[41\] a_16076_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7843 vssd1 _0330_ a_11847_3073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7844 a_16566_22173# a_16293_21807# a_16481_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7845 vssd1 a_25042_5461# a_24971_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7848 a_3339_23983# _0804_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X7849 a_20414_22325# a_20246_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7851 a_10497_1679# a_9963_1685# a_10402_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7852 vssd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_2961_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7853 dec1.i_ones a_7959_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7854 a_12613_1679# a_12079_1685# a_12518_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7855 vssd1 a_23915_17129# a_23922_17033# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7856 vccd1 a_7891_5461# a_7715_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X7857 vccd1 _0440_ a_17323_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X7858 vccd1 _0251_ a_24315_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7859 a_15289_15823# _0554_ _0555_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7860 net25 a_9595_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7861 vccd1 a_2010_24759# _0416_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X7862 a_21970_18231# _0480_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X7864 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7865 _0458_ a_21003_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7866 vssd1 a_15439_2388# _0179_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7867 a_5007_19087# _0740_ a_4805_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7868 a_1769_9615# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7870 a_8390_23439# clknet_0__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7871 vccd1 cal_lut\[22\] a_14277_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X7872 vccd1 a_18659_10615# _0623_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7874 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_1407_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X7875 a_23145_15279# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7876 a_11317_25321# _0729_ a_11189_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X7878 a_4307_27574# _0829_ a_3848_27399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X7879 a_21709_26159# a_21155_26133# a_21362_26133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7880 a_22856_6409# a_22457_6037# a_22730_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7881 a_27732_12937# a_27333_12565# a_27606_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7884 a_15170_21237# a_15002_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7885 a_18689_13647# _0011_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7886 vssd1 a_19862_11039# a_19820_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7887 vccd1 net46 a_17783_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7888 a_21291_26159# a_21162_26433# a_20871_26133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7889 a_11506_15645# a_11233_15279# a_11421_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7890 vssd1 io_in[2] a_1407_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7891 _0622_ a_16771_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7892 vssd1 _0098_ a_12141_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7893 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7894 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7895 vssd1 _0867_ a_21095_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7896 a_19865_13621# _0530_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7897 a_13415_20884# _0883_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7899 vssd1 a_18942_13621# a_18900_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7900 a_15381_12015# _0514_ a_15299_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7901 a_7381_9839# a_7111_10205# a_7291_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X7902 a_20683_21972# _0241_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7903 a_3151_14735# _0390_ a_2933_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7904 a_10202_15797# a_10034_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7905 _0641_ a_22659_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7906 vssd1 a_15795_28879# a_15963_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7907 _0843_ a_9223_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X7908 vccd1 a_9815_14557# a_9983_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7909 vccd1 a_14155_3285# _0313_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X7912 temp1.capload\[0\].cap.Y net49 a_2689_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7913 cal_lut\[87\] a_25439_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7914 a_8795_4943# a_8013_4949# a_8711_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7915 a_25203_10901# net36 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7916 a_10197_25223# _0731_ a_10443_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7917 vccd1 a_25823_23439# a_25991_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7918 a_27774_17567# a_27606_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7919 cal_lut\[139\] a_5843_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7920 a_18390_28853# a_18222_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7922 a_24665_15829# a_24499_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7923 a_8447_7338# _0308_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7924 a_19743_25615# a_18961_25621# a_19659_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7925 a_18255_7663# a_18119_7637# a_17835_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7926 _0051_ a_17415_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7927 a_19256_20969# cal_lut\[52\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X7928 vccd1 _0295_ a_20727_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7929 a_23936_9839# cal_lut\[171\] a_23361_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X7930 vssd1 net46 a_20267_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7931 a_5801_26409# _0409_ _0410_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7932 vccd1 a_18027_19783# _0468_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7933 _0012_ a_20635_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7934 a_18475_5639# _0445_ a_18709_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7935 vssd1 _0361_ a_25051_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7936 vccd1 a_6791_4074# _0133_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7937 vccd1 a_15779_1653# a_15695_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7938 vssd1 a_4277_27221# a_4211_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7939 vssd1 a_25823_23439# a_25991_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7940 a_10317_3311# _0146_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7941 a_17677_25071# _0046_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7942 a_20132_19394# dbg_result[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X7943 a_10034_15823# a_9761_15829# a_9949_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7944 a_17565_13621# _0593_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7946 a_8999_7828# _0303_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7947 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7948 vssd1 cal_lut\[107\] a_17961_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7949 _0038_ a_9411_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7950 _0485_ a_13942_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7951 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7952 a_21997_1685# a_21831_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7953 a_3685_22325# clknet_0_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7954 a_18192_15529# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7955 a_16035_6144# cal_lut\[119\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7957 a_8251_29789# a_7553_29423# a_7994_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7958 vccd1 a_20499_8439# _0583_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X7959 cal_lut\[192\] a_14031_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7960 a_20648_21641# a_20249_21269# a_20522_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7961 vssd1 a_25623_17973# a_25581_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7962 a_4616_17455# _0476_ a_4313_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X7963 a_27498_8863# a_27330_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7964 vccd1 net41 a_14655_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7965 a_22872_21263# _0636_ a_22770_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X7966 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_3056_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X7967 a_17459_29185# _0216_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7968 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7969 _0358_ a_27071_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X7970 cal_lut\[192\] a_14031_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7971 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd _0817_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7972 a_9187_29111# a_9478_29001# a_9429_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7973 vccd1 _0087_ a_21709_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7974 vccd1 a_12927_17723# a_12843_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7975 cal_lut\[67\] a_22955_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7976 a_4897_20719# _0427_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X7977 vssd1 a_21334_4511# a_21292_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7978 _0302_ a_7704_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X7979 a_19664_27497# _0222_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7980 a_6646_21041# _0425_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X7981 a_27219_15253# a_27510_15553# a_27461_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7982 temp1.capload\[7\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7984 vssd1 a_22711_6549# _0343_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X7985 a_8251_9117# a_7387_8751# a_7994_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7986 vccd1 _0811_ a_4528_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X7988 vccd1 _0498_ a_11693_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7990 vccd1 _0431_ a_6375_19095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X7991 a_9021_29575# a_9117_29397# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X7992 a_3299_19061# _0424_ a_3517_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X7993 a_3953_10761# a_3406_10505# a_3606_10660# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7994 a_11416_27247# a_10423_27247# a_11287_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X7995 a_15262_27765# a_15094_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7996 cal_lut\[133\] a_8695_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7997 vssd1 cal_lut\[170\] a_24964_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X7998 _0164_ a_24039_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7999 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4988_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X8000 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8001 vccd1 a_22787_14735# a_22955_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8002 a_7741_13103# _0019_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8003 vssd1 net25 a_11987_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8004 vssd1 _0341_ a_26107_8725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8005 a_15281_12565# a_15115_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8007 a_18637_19631# net18 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X8008 vssd1 _0332_ a_14103_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8009 a_21913_11471# _0449_ a_21997_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8011 vccd1 a_22403_22075# a_22319_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8013 vccd1 a_17197_19777# _0582_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8014 a_18072_26159# a_17673_26159# a_17946_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8015 a_6648_24847# _0792_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X8016 a_1477_10901# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8017 vssd1 temp1.dac.vdac_single.en_pupd a_3247_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8018 vccd1 _0714_ a_8951_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8019 a_14287_8320# cal_lut\[112\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8020 vccd1 cal_lut\[168\] a_25783_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8021 vccd1 a_3606_10660# a_3535_10761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8022 _0414_ a_2419_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8023 a_23263_26935# a_23547_26921# a_23482_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8024 _0866_ a_18192_15529# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X8025 vssd1 a_5843_3829# a_5801_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8026 a_3991_26409# _0414_ _0784_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8027 a_4816_16617# clknet_1_0__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8028 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8029 vccd1 net36 a_22107_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8030 a_6244_25045# _0805_ a_6636_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X8031 a_7553_16367# a_7387_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8032 vccd1 clknet_0__0380_ a_6537_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8033 a_17489_25071# a_17323_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8034 vssd1 a_11605_16055# _0844_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X8036 a_14845_10927# cal_lut\[190\] a_14773_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8037 a_17489_23983# a_17323_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8038 a_9326_20719# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X8041 a_11781_13103# cal_lut\[81\] a_11343_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8042 a_8270_3829# a_8102_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8043 vccd1 a_28031_10205# a_28199_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8044 a_22009_27247# a_21739_27613# a_21919_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X8045 _0052_ a_19531_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8047 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8049 a_15094_29789# a_14655_29423# a_15009_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8050 a_17094_20407# _0582_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X8051 a_8289_14741# a_8123_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8052 _0577_ a_16679_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8053 vccd1 a_18723_3579# a_18639_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8054 temp1.capload\[8\].cap.Y net63 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8055 vccd1 net35 a_19255_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8056 vssd1 _0440_ a_17323_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8057 a_16373_16341# _0613_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X8058 vccd1 a_11579_3829# _0363_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8059 vssd1 a_3575_15797# _0379_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0991 ps=0.955 w=0.65 l=0.15
X8060 vccd1 cal_lut\[107\] a_17536_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8061 a_24846_25437# a_24573_25071# a_24761_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8062 a_8887_15823# a_8105_15829# a_8803_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8063 a_18298_3423# a_18130_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8064 a_25507_10383# a_25327_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8065 vccd1 a_1921_11989# _0200_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8067 vccd1 clknet_1_1__leaf__0380_ a_9319_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.173 ps=1.82 w=0.64 l=0.15
X8068 vssd1 net44 a_16127_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8069 vssd1 a_3759_21495# _0782_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X8070 a_1551_19605# _0761_ a_2614_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8071 vssd1 net26 a_14747_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8072 a_23450_7775# a_23282_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8073 _0220_ a_16904_25321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X8074 a_11715_21379# _0664_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8075 a_11508_20719# _0678_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X8077 a_27521_12559# _0172_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8078 a_22396_28169# a_21997_27797# a_22270_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8079 vssd1 _0421_ a_2931_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8080 a_15469_3855# _0178_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8081 vssd1 a_3995_18793# _0759_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8082 a_25397_7497# a_24407_7125# a_25271_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8083 vssd1 a_20287_28603# a_20245_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8084 a_10236_8751# _0476_ a_10046_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X8085 vssd1 net20 a_19961_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8086 a_20755_22351# a_19973_22357# a_20671_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8087 _0160_ a_25879_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8088 vssd1 _0438_ a_14006_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.107 ps=0.98 w=0.65 l=0.15
X8089 cal_lut\[145\] a_7775_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8090 a_11693_10383# cal_lut\[147\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8091 a_2794_28662# _0419_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X8092 cal_lut\[104\] a_21759_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8093 a_25800_17455# a_25401_17455# a_25674_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8094 vccd1 _0316_ a_5179_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8095 a_7994_8863# a_7826_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8096 vccd1 a_9091_29111# ctr\[12\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8097 vssd1 cal_lut\[13\] a_22388_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X8098 vssd1 net22 a_1917_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8099 _0452_ a_20690_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8100 vssd1 a_24351_14735# a_24519_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8101 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X8102 _0442_ a_14523_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8103 a_4351_31055# _0817_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8104 a_11891_10205# a_11711_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8105 vccd1 _0445_ a_15943_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8106 a_21591_11293# a_20727_10927# a_21334_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8108 dbg_result[0] a_7410_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X8109 vssd1 cal_lut\[7\] a_12533_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8110 a_2722_20175# _0422_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X8111 vccd1 _0454_ a_17231_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8112 vssd1 a_13146_25183# a_13104_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8113 vccd1 _0437_ a_7025_21041# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8114 vccd1 _0433_ a_8297_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8115 a_11966_7119# a_11693_7125# a_11881_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8116 a_22719_27221# net47 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8118 vssd1 _0481_ a_19777_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8120 vccd1 net33 a_22199_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8121 vccd1 net27 a_3799_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8122 vssd1 _0856_ a_23671_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8123 vccd1 a_11195_28701# a_11366_28588# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X8124 a_4892_20175# _0747_ a_4801_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X8125 a_22839_6575# cal_lut\[158\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X8126 a_25203_10901# net36 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8127 vssd1 a_15687_27765# a_15645_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8128 a_21879_16055# _0505_ a_22113_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8129 a_8270_3829# a_8102_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8130 a_10691_29673# net13 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X8131 a_4866_5599# a_4698_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8132 a_21978_21919# a_21810_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8133 vccd1 _0428_ a_4253_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X8134 vccd1 cal_lut\[98\] a_11891_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8135 vssd1 a_25387_5161# a_25394_5065# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8136 a_27035_8181# a_27211_8513# a_27163_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X8137 _0110_ a_19807_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8138 a_23110_3044# a_22903_2985# a_23286_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8140 vssd1 a_20839_22325# a_20797_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8141 _0808_ a_2695_14013# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=1.62 w=1 l=0.15
X8142 vccd1 a_9765_6727# _0309_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X8143 a_21261_11293# a_20727_10927# a_21166_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8145 a_14450_24527# a_14011_24533# a_14365_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8146 vccd1 _0709_ a_11900_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X8147 vccd1 cal_lut\[185\] a_18272_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8148 a_6246_16503# a_6087_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X8150 vccd1 a_19763_4074# _0117_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8151 a_2794_28335# _0419_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X8152 a_11601_3311# a_11435_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8153 a_6737_22351# _0786_ a_6939_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8154 vccd1 _0464_ a_15727_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8155 a_3575_15797# a_4027_16144# a_3985_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8158 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8159 a_7060_31751# net10 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X8160 a_22546_13469# a_22107_13103# a_22461_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8161 vccd1 _0424_ a_2222_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X8162 a_17651_28023# a_17942_27913# a_17893_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8163 vccd1 a_8251_13469# a_8419_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8164 vssd1 a_28199_17723# a_28157_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8165 a_4977_3861# a_4811_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8166 _0172_ a_27351_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8167 a_25161_11293# a_24823_11079# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8168 a_10258_10383# _0513_ a_10178_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8169 net34 a_17415_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X8172 vssd1 a_15909_7809# _0546_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8173 a_25271_24349# a_24407_23983# a_25014_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8174 vssd1 _0425_ _0381_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8175 a_2489_8181# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R20 vssd1 net50 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8176 a_1673_22351# ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8177 a_8335_6941# a_7553_6575# a_8251_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8178 cal_lut\[66\] a_21115_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8179 vssd1 a_15595_21237# a_15553_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8180 a_8286_4943# a_7847_4949# a_8201_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8181 _0673_ a_11191_19659# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X8182 a_4487_13077# _0390_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.178 ps=1.4 w=0.42 l=0.15
X8183 a_15904_25589# net47 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X8184 vccd1 a_4027_16144# a_3575_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X8186 a_23489_22895# _0469_ a_23055_23047# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8187 vccd1 a_19862_4511# a_19789_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8188 a_20322_9269# a_20154_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8189 a_4974_8029# a_4701_7663# a_4889_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8190 a_25271_9117# a_24573_8751# a_25014_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8191 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8192 a_3785_17999# _0421_ a_4143_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8193 vssd1 a_26283_8207# a_26451_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8194 a_15262_27765# a_15094_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8195 _0841_ a_13459_22359# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X8196 a_14353_18793# _0425_ a_14550_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8197 a_20437_3311# _0156_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8198 a_14269_1135# a_14103_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8199 a_14006_19407# _0447_ a_13892_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X8200 a_22205_14013# cal_lut\[174\] a_22133_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8201 a_7975_18909# a_7111_18543# a_7718_18679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8202 vssd1 _0341_ a_24635_8513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8203 a_6940_12937# a_6541_12565# a_6814_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8204 _0795_ _0737_ a_5553_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8205 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8206 _0124_ a_13183_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8207 a_10832_30663# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8208 a_10883_25071# _0718_ _0749_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.106 ps=0.975 w=0.65 l=0.15
X8209 vssd1 _0414_ _0419_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8210 a_18015_5639# _0445_ a_18249_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8211 a_13714_28879# a_13441_28885# a_13629_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8212 a_15695_13647# a_14913_13653# a_15611_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8213 vccd1 a_17095_5639# _0614_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X8214 vccd1 _0352_ a_25695_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8215 a_25594_5220# a_25387_5161# a_25770_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8216 vccd1 a_6703_6549# _0327_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X8217 a_6909_10389# a_6743_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8218 vssd1 a_27371_22075# a_27329_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8219 _0375_ a_5451_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8220 _0107_ a_18519_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8221 a_7994_29535# a_7826_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8222 a_5077_24233# _0796_ a_4931_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X8223 a_5617_15431# a_5713_15253# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X8224 a_17029_18005# a_16863_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8225 vccd1 a_4222_12533# a_4149_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8226 vssd1 a_17565_13621# _0596_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8227 a_15094_27791# a_14821_27797# a_15009_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8228 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8229 vssd1 _0363_ a_11019_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8230 vccd1 a_20141_6005# _0586_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8231 vccd1 a_14703_21972# _0040_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8232 a_10596_17705# _0662_ a_10505_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X8233 a_12610_14557# a_12171_14191# a_12525_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8236 a_23873_16911# a_23535_17143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8237 a_23792_10089# _0510_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X8238 a_20417_13249# _0526_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X8239 vssd1 a_11120_28853# net13 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X8241 a_27701_10205# a_27167_9839# a_27606_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8242 a_5805_16367# a_5639_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8243 a_17627_14735# a_16845_14741# a_17543_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8245 a_5460_15823# clknet_1_0__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8246 a_11172_14191# a_10773_14191# a_11046_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8247 a_5359_8207# a_5179_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8248 vssd1 a_3891_17455# _0755_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X8250 a_7289_25321# _0734_ a_7071_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8251 a_14616_14709# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8253 a_26367_8207# a_25585_8213# a_26283_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8254 _0355_ a_25507_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8255 a_16179_29397# cal_lut\[44\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X8256 a_25559_10927# a_25339_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8257 vccd1 a_11458_27500# dbg_result[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X8258 vssd1 _0626_ a_10562_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8259 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8260 vccd1 _0444_ a_21997_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X8261 a_18475_19783# net18 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8264 temp1.dac_vout_notouch_ net14 a_11868_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X8265 a_14910_7119# a_14637_7125# a_14825_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8266 a_22503_24135# cal_lut\[31\] a_22649_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X8267 a_14550_18793# a_14770_18517# _0472_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8268 a_11723_8751# a_11594_9025# a_11303_8725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8269 a_6651_18793# _0839_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8270 a_13805_9673# a_12815_9301# a_13679_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8271 a_8491_24847# _0713_ a_8397_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X8272 a_15469_20407# _0872_ a_15632_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8273 vssd1 a_24455_19783# cal_lut\[28\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8274 a_7097_6031# _0144_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8275 vssd1 a_7407_7093# a_7365_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8276 a_14457_7663# _0124_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8277 a_22165_10357# _0634_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X8278 a_8483_31599# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X8279 a_2652_28487# _0801_ a_2794_28662# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X8283 a_14710_1247# a_14542_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8284 a_18659_10615# _0514_ a_18893_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8287 vccd1 net44 a_16127_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8288 vssd1 a_14747_20175# net20 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8289 a_14545_5487# a_14379_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8290 vccd1 a_17555_28023# cal_lut\[91\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8291 vccd1 net41 a_7387_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8295 a_2576_26703# a_2327_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X8296 a_13698_23413# a_13530_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8297 vccd1 a_12311_11079# cal_lut\[98\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8298 a_21031_21263# a_20249_21269# a_20947_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8299 a_17244_15113# a_16845_14741# a_17118_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8300 a_15193_15431# _0505_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X8301 a_16340_7913# _0498_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X8302 a_12893_22895# _0081_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8303 a_23286_2767# a_23039_3145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8304 vccd1 a_8263_15444# _0078_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8305 a_20666_13353# _0528_ a_20417_13249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8306 vccd1 _0863_ a_23211_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8307 a_12525_18231# cal_lut\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X8308 a_14747_27497# _0487_ a_14829_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X8309 a_16983_23047# cal_lut\[82\] a_17129_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X8311 a_7439_4373# net1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X8312 vccd1 a_10740_29575# a_10691_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X8314 a_9049_30761# _0817_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8315 vccd1 net7 a_2417_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X8316 vccd1 a_8527_3855# a_8695_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8317 vccd1 a_19683_2197# a_19690_2497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8318 _0834_ a_4003_30006# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X8319 vccd1 temp1.i_precharge_n a_2778_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8320 vccd1 a_18111_25589# net46 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8321 vssd1 cal_lut\[3\] a_9687_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8322 vccd1 a_21334_11039# a_21261_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8323 vccd1 a_9005_24501# _0728_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8324 a_5841_19605# _0737_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X8325 a_15446_2741# a_15278_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8326 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X8327 a_20203_28701# a_19421_28335# a_20119_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8328 a_9358_3855# _0495_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X8329 a_1677_6575# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8331 a_7994_11039# a_7826_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8332 vssd1 a_10239_31055# net14 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8333 vccd1 _0400_ a_6377_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8334 a_3169_25935# _0418_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X8335 a_16481_27247# _0042_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8336 vssd1 net24 a_6743_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8337 vccd1 a_20287_11195# a_20203_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8339 vssd1 a_13691_28500# _0049_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8340 vccd1 cal_lut\[56\] a_23481_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X8342 net8 a_10844_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8343 a_19426_20719# _0559_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X8344 a_13838_19319# _0442_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8345 vccd1 _0341_ a_25603_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8346 vssd1 _0444_ a_20716_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X8347 a_2309_11791# _0389_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8348 vccd1 cal_lut\[93\] a_14283_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8349 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8350 a_6929_21583# _0778_ a_6519_21495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X8351 vssd1 _0376_ a_5639_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8352 a_5227_26935# _0811_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8353 vccd1 a_25187_15041# a_25011_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X8354 vccd1 net36 a_26891_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8355 _0362_ a_25047_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8357 vssd1 a_8803_1679# a_8971_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8358 a_6269_29423# _0209_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8359 vccd1 a_8539_2986# _0180_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8360 _0597_ a_15943_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X8361 a_11857_18517# _0556_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X8362 vssd1 a_16640_4373# net31 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X8363 net18 a_14287_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X8364 cal_lut\[148\] a_13019_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8365 vccd1 _0481_ a_19255_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8366 cal_lut\[1\] a_4831_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8367 a_25755_11989# net36 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8369 a_7157_19319# clknet_1_1__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X8370 a_18271_25437# a_17489_25071# a_18187_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8372 a_25770_4943# a_25523_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8373 _0818_ _0434_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X8374 cal_lut\[184\] a_13111_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8375 a_22177_6575# a_21187_6575# a_22051_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8376 a_21169_11471# cal_lut\[104\] a_21085_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8377 _0189_ a_5639_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8378 a_17105_10357# _0515_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X8379 vccd1 a_25014_24095# a_24941_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8380 vssd1 _0541_ a_15725_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X8381 vccd1 cal_lut\[96\] a_16156_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8382 vccd1 _0495_ a_15943_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X8383 a_8412_5321# a_8013_4949# a_8286_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8384 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8385 a_10961_5487# _0128_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8386 a_4893_14441# _0809_ _0398_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8387 vccd1 a_18326_7637# a_18255_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8388 vssd1 a_16975_11195# a_16933_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8389 _0075_ a_26063_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8390 vccd1 a_4167_16367# _0839_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8391 a_11547_24847# _0711_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8392 a_25271_23261# a_24407_22895# a_25014_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8395 a_27847_7119# a_26983_7125# a_27590_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8396 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8397 vssd1 a_25106_15797# a_25064_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8398 a_7791_27613# a_7093_27247# a_7534_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8399 cal_lut\[157\] a_21115_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8400 a_4663_10205# a_3965_9839# a_4406_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8401 a_15553_21641# a_14563_21269# a_15427_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8402 a_24771_21085# a_24591_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8403 a_9647_14709# cal_lut\[79\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X8404 a_12977_2223# a_11987_2223# a_12851_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8405 _0140_ a_2971_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8406 a_4407_15529# _0387_ a_4091_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X8407 a_25713_12381# a_25375_12167# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X8408 a_4431_26159# ctr\[6\] _0784_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X8409 vccd1 a_7718_18679# a_7652_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X8410 a_2566_15797# a_2398_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8412 vssd1 a_17555_28023# cal_lut\[91\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8413 a_26318_16733# a_25879_16367# a_26233_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8414 _0376_ a_5083_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8416 a_28115_17821# a_27333_17455# a_28031_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8417 vccd1 _0340_ a_19807_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8418 a_14158_26677# a_13990_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8419 a_1639_15444# _0388_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8420 vccd1 a_27774_9951# a_27701_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8421 vccd1 _0363_ a_8951_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8423 a_21081_4399# _0114_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8424 _0444_ a_20943_6369# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X8425 vccd1 net26 a_14103_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8426 vssd1 a_25927_13255# cal_lut\[175\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8427 a_25471_20407# a_25762_20297# a_25713_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8428 vssd1 a_6319_11293# a_6487_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8429 vssd1 _0263_ a_22291_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8430 vccd1 cal_lut\[33\] a_24771_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8431 a_17526_19881# _0580_ a_17446_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8432 a_17861_26159# _0088_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8435 a_10380_19783# _0629_ a_10522_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8436 a_27590_17973# a_27422_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8437 a_15715_5175# _0440_ a_15949_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8438 a_27347_14557# a_27167_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8439 vssd1 _0331_ a_11711_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8441 vssd1 _0561_ a_13091_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8442 a_14655_18115# dbg_result[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8443 a_13035_14557# a_12171_14191# a_12778_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8444 a_13809_4943# a_13275_4949# a_13714_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8445 a_17187_13255# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8446 vccd1 a_6633_26703# a_6739_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X8447 cal_lut\[96\] a_15963_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8448 a_26094_15939# _0246_ a_26012_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8449 _0001_ a_7387_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8450 vccd1 a_15071_13268# _0010_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8451 vssd1 a_18142_28068# a_18071_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X8452 _0454_ a_18519_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X8453 a_10517_23983# _0705_ a_10083_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8454 a_13261_21263# _0039_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8455 a_11157_17705# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.148 ps=1.34 w=0.42 l=0.15
X8456 a_19167_19061# dbg_result[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X8457 _0690_ a_14747_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8458 vssd1 _0154_ a_20237_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8459 _0849_ a_13363_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8460 a_4988_31375# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X8461 vccd1 a_20579_9295# a_20747_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8463 temp1.capload\[6\].cap.Y net61 a_1769_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8464 a_20579_9295# a_19881_9301# a_20322_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8465 a_4678_26311# ctr\[1\] a_4998_26165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8467 a_15101_13647# _0010_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8468 _0410_ ctr\[9\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8470 vssd1 cal_lut\[81\] a_12120_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8471 _0875_ a_23391_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8472 vssd1 a_1959_21807# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8473 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8474 vccd1 net31 a_17691_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8475 a_19583_2741# a_19759_3073# a_19711_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X8476 vccd1 cal_lut\[139\] a_6555_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8477 a_17961_27247# a_17691_27613# a_17871_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X8478 a_16109_10927# a_15943_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8479 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_2576_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X8480 a_18387_9527# a_18678_9417# a_18629_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8481 vccd1 a_16737_13621# _0600_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8482 a_8527_3855# a_7663_3861# a_8270_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8483 vssd1 cal_lut\[13\] a_21825_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8484 vssd1 a_15715_30186# _0044_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8485 a_25397_25071# a_24407_25071# a_25271_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8486 vccd1 _0276_ a_12815_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8487 a_7716_25589# _0734_ a_8108_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X8489 vssd1 _0448_ a_15023_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8490 _0747_ a_3072_19637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X8491 a_6537_19605# clknet_0__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8492 a_25389_19631# a_24842_19905# a_25042_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8493 vssd1 clknet_1_0__leaf_io_in[0] a_4811_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8495 vccd1 _0344_ a_24315_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8497 _0043_ a_17047_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8499 vccd1 a_4277_27221# a_4307_27574# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8500 cal_lut\[14\] a_23139_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8501 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8502 cal_lut\[38\] a_8419_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8504 vssd1 a_15043_24501# a_15001_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8505 _0531_ a_17783_21271# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8506 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8507 a_3111_28662# _0800_ a_2652_28487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8508 vccd1 a_9275_28023# _0816_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X8509 a_12299_3677# a_11435_3311# a_12042_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8510 vccd1 net27 a_7387_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8512 a_12688_18115# cal_lut\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X8515 _0669_ _0663_ a_10055_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8516 net7 a_1407_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X8517 vccd1 a_9371_2741# _0367_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X8519 cal_lut\[105\] a_21759_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8520 a_15453_12015# cal_lut\[192\] a_15381_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8521 vssd1 a_7994_16479# a_7952_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8522 a_8987_14735# a_8289_14741# a_8730_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8523 a_21883_1109# cal_lut\[151\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X8525 a_9482_6031# a_9209_6037# a_9397_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8526 a_21265_7815# _0283_ a_21428_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8527 a_24835_5461# net33 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8528 vssd1 a_1741_30199# a_1554_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8529 a_21362_26133# a_21155_26133# a_21538_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8530 a_9297_12879# cal_lut\[79\] a_8951_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8532 vssd1 a_8270_3829# a_8228_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8534 _0701_ a_9043_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X8535 _0359_ a_27531_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8536 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8537 a_15193_14343# cal_lut\[10\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X8538 a_23815_4087# a_24106_3977# a_24057_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8539 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_2327_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8540 a_11794_8725# a_11594_9025# a_11943_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8541 vccd1 a_11587_8725# a_11594_9025# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8542 vccd1 cal_lut\[163\] a_24262_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X8543 vssd1 a_20417_13249# _0529_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8544 a_27710_15253# a_27510_15553# a_27859_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8545 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8548 a_4443_18793# _0426_ _0427_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8549 a_21675_4765# a_20893_4399# a_21591_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8550 _0306_ a_13592_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X8551 a_2014_14709# a_1846_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8553 a_12035_26324# _0846_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8555 _0437_ a_7111_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X8557 a_24075_19087# a_23377_19093# a_23818_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8558 a_22438_1653# a_22270_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8559 a_21591_10205# a_20893_9839# a_21334_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8561 vccd1 a_13537_15431# _0255_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X8562 a_25401_17455# a_25235_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8563 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8564 a_3370_11177# _0391_ a_3288_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8565 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8567 a_27583_9514# _0356_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8568 vccd1 _0015_ a_25389_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X8569 vssd1 _0773_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8570 a_15531_24135# _0460_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8571 vccd1 a_25375_20407# cal_lut\[34\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8572 _0661_ _0660_ a_12351_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.13 ps=1.26 w=1 l=0.15
X8573 vssd1 a_3081_28309# a_3015_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X8574 a_4211_23983# _0411_ a_3848_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X8575 vssd1 a_6674_16620# a_6632_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X8576 vssd1 net2 a_3155_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X8578 vccd1 _0448_ a_14747_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X8579 a_6184_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X8580 a_11152_30287# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X8581 vssd1 _0465_ a_18731_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8582 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X8583 a_3575_15797# net69 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X8586 vccd1 _0328_ a_7571_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8587 a_7607_6031# a_6909_6037# a_7350_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8588 vccd1 a_15687_29691# a_15603_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8589 vccd1 _0841_ a_8123_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X8590 _0245_ a_25047_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8591 vssd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8592 vccd1 a_9835_26703# _0385_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8593 vccd1 _0451_ a_9595_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X8594 vccd1 a_24635_8513# a_24459_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X8596 a_21825_13103# a_21555_13469# a_21735_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X8597 vssd1 a_9184_20871# _0627_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X8598 _0767_ ctr\[4\] a_5998_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X8599 vssd1 net44 a_22291_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X8600 a_7350_10357# a_7182_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8601 vccd1 a_15255_28500# _0091_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8602 vssd1 a_19915_19087# _0443_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X8603 vccd1 _0630_ a_10454_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X8605 cal_lut\[140\] a_6947_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8606 cal_lut\[141\] a_4831_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8608 vccd1 _0858_ a_14839_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8610 _0100_ a_14287_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8611 a_6647_28585# _0390_ a_6429_28309# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8612 vccd1 cal_lut\[174\] a_21971_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X8613 vccd1 a_25014_23007# a_24941_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8614 a_24591_21085# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8615 a_4437_15055# a_4245_14796# _0205_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X8616 vccd1 a_1736_18517# _0744_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8617 a_8546_15797# a_8378_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8618 a_7005_4551# _0299_ a_7168_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8619 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2419_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8620 vssd1 _0552_ a_17381_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X8621 a_9305_14191# _0079_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8622 _0155_ a_17415_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8623 _0340_ a_19435_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8624 a_26226_6941# a_25787_6575# a_26141_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8625 a_9905_21263# _0591_ a_9821_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8626 _0266_ a_12355_21271# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X8627 vssd1 _0483_ a_9436_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X8628 a_7182_10383# a_6909_10389# a_7097_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8629 vccd1 _0447_ a_12950_16988# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X8630 _0016_ a_14839_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8631 a_4713_21583# ctr\[3\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8632 _0505_ a_17323_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8633 a_4663_9117# a_3965_8751# a_4406_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8634 vccd1 _0281_ a_18335_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8635 a_9749_16617# _0702_ a_9595_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X8636 a_14155_3285# cal_lut\[131\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X8637 vssd1 _0305_ a_11527_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8638 vccd1 _0454_ a_16035_18112# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8639 a_10197_25223# _0718_ a_10347_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X8641 a_11684_22671# _0672_ _0710_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.393 ps=2.51 w=0.65 l=0.15
X8642 a_21919_27613# a_21739_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8643 vssd1 net42 a_26983_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8644 a_8251_16733# a_7387_16367# a_7994_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8645 a_26861_13103# a_26314_13377# a_26514_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
R21 vccd1 temp1.capload\[6\].cap_61.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8647 a_22903_21959# _0460_ a_23077_21835# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8648 a_16771_8751# cal_lut\[125\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8649 a_20706_27791# a_20267_27797# a_20621_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8650 vssd1 a_13771_21263# a_13939_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8651 vccd1 _0453_ a_17783_21271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X8653 a_21591_11293# a_20893_10927# a_21334_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8654 a_17935_28009# net46 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8655 vssd1 _0396_ a_3420_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8656 a_11765_17973# _0587_ a_12052_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X8657 _0354_ a_25783_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8658 _0107_ a_18519_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8659 a_7534_27359# a_7366_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8660 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8662 a_3015_28335# _0801_ a_2652_28487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X8663 a_16076_21379# _0872_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8664 a_10743_19631# dbg_result[5] a_10380_19783# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X8665 vccd1 _0675_ a_10943_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8666 a_6982_17973# a_6823_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8667 a_2708_14191# a_2309_14191# a_2582_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8668 vssd1 a_17105_10357# _0624_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X8671 vssd1 a_25410_10901# a_25339_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X8672 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8673 vccd1 net8 a_10515_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X8674 a_20621_27791# _0053_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8675 a_13257_23445# a_13091_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8676 _0670_ _0667_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8677 vssd1 _0471_ a_21970_18231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8680 a_25502_21781# a_25295_21781# a_25678_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8681 _0571_ a_12539_6144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8682 a_1585_8751# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8683 a_9390_1501# a_9117_1135# a_9305_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8684 a_22719_27221# net47 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8685 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8687 a_4805_19087# _0430_ a_5007_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8688 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8690 a_2108_15529# _0428_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X8691 vssd1 a_7350_10357# a_7308_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8692 a_16109_10927# a_15943_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8694 vssd1 a_2652_28487# _0832_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X8695 vssd1 a_3112_19783# a_3072_19637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8697 a_1541_19087# a_1471_19319# _0423_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X8699 vccd1 _0439_ a_8975_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8700 a_22806_3829# a_22638_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8701 vssd1 _0872_ a_14273_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8702 vccd1 net26 a_13275_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8703 vssd1 a_2722_20175# _0424_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X8704 a_23457_3145# a_22910_2889# a_23110_3044# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X8705 _0015_ a_23763_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8706 vssd1 _0043_ a_17845_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8707 a_15569_27247# cal_lut\[92\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X8710 vccd1 cal_lut\[60\] a_20775_18231# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X8711 vssd1 a_15531_4564# _0178_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8712 a_20157_16917# a_19991_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8713 a_25431_21807# a_25295_21781# a_25011_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8714 _0434_ _0422_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8716 vssd1 a_5142_7775# a_5100_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8717 vccd1 _0715_ a_9858_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X8718 a_16117_18365# _0454_ a_16035_18112# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8719 a_19303_2375# a_19399_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X8720 a_23707_8029# a_22843_7663# a_23450_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8721 a_1584_27023# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X8722 a_23355_10615# cal_lut\[109\] a_23481_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X8723 a_7607_10383# a_6909_10389# a_7350_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8725 a_12141_8751# a_11587_8725# a_11794_8725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8726 _0676_ _0666_ a_10969_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8727 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8728 cal_lut\[30\] a_21023_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8729 vssd1 cal_lut\[16\] a_14565_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X8730 a_19789_5853# a_19255_5487# a_19694_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8731 vssd1 _0237_ a_25187_15041# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8732 _0877_ a_24771_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8733 vssd1 a_25203_10901# a_25210_11201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8735 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8736 vssd1 _0453_ a_18151_21271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8737 a_19659_25615# a_18795_25621# a_19402_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8738 _0637_ a_21923_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X8739 a_4771_20871# net21 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X8740 a_16013_19631# a_15023_19631# a_15887_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8742 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8743 _0410_ _0409_ a_5801_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8744 a_10784_23983# _0681_ a_10699_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8745 a_10317_7119# _0122_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8746 _0265_ a_21872_25731# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X8747 a_3685_22325# clknet_0_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8748 vssd1 _0363_ a_16079_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8749 a_5418_3829# a_5250_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8750 a_12341_2223# _0147_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8751 a_18390_28853# a_18222_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8754 a_18865_12937# a_17875_12565# a_18739_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8755 _0475_ a_18369_18337# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X8756 a_19890_2197# a_19683_2197# a_20066_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8757 a_14269_1135# a_14103_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8758 a_8947_11471# a_8767_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8759 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5087_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X8760 a_25103_5175# a_25394_5065# a_25345_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X8761 a_14967_1501# a_14103_1135# a_14710_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8762 a_9326_21046# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X8763 vssd1 cal_lut\[51\] a_16949_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8764 vccd1 a_11302_16519# _0629_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X8765 a_17961_8751# a_17691_9117# a_17871_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X8766 vssd1 _0836_ a_2773_9991# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8767 vccd1 _0748_ a_7653_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8768 vssd1 _0425_ _0485_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8769 a_8975_18793# _0433_ _0680_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X8770 _0521_ a_8645_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.373 ps=1.75 w=1 l=0.15
X8771 vccd1 _0765_ a_8309_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8772 a_2566_15797# a_2398_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8773 a_12709_27247# _0007_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8774 vccd1 _0452_ a_16803_22689# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8775 a_7550_14557# a_7111_14191# a_7465_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8776 vccd1 a_16147_12533# a_16063_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8777 vccd1 cal_lut\[162\] a_26519_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8778 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_2327_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X8780 vccd1 net46 a_19439_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8781 a_15483_8751# cal_lut\[126\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8782 a_15370_19407# _0442_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X8783 vccd1 a_10835_4161# a_10659_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X8784 a_18807_9673# a_18678_9417# a_18387_9527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8785 a_18659_10615# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X8786 a_14103_27497# _0487_ a_14185_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8787 net81 a_15023_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8788 vssd1 a_22787_14735# a_22955_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8789 vssd1 a_26451_8181# a_26409_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8790 a_23110_3044# a_22910_2889# a_23259_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8791 a_20437_21263# _0065_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8792 vssd1 a_11029_17429# _0663_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X8793 a_2398_15823# a_2125_15829# a_2313_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8794 _0239_ a_25415_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8795 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8796 a_25849_21807# a_25295_21781# a_25502_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8797 a_5805_16367# a_5639_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8798 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8799 _0772_ a_1963_21365# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.1 w=0.65 l=0.15
X8800 a_5376_13103# a_4977_13103# a_5250_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8801 a_26352_6575# a_25953_6575# a_26226_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8802 a_25431_21807# a_25302_22081# a_25011_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X8803 vssd1 a_4310_8439# a_4259_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8804 temp1.capload\[10\].cap.Y net50 a_2505_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8805 _0760_ a_4283_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8806 a_21971_13879# _0505_ a_22205_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8807 a_27802_13924# a_27602_13769# a_27951_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8808 vccd1 _0434_ a_8383_22583# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X8809 vccd1 a_19862_11039# a_19789_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8810 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8811 vssd1 net40 a_14655_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8813 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8814 a_10459_15823# a_9761_15829# a_10202_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8815 a_24035_7119# a_23855_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8816 a_2413_8751# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8817 vssd1 net29 a_15115_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8819 a_6239_27247# a_6019_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8820 a_22837_27069# a_22567_26703# a_22747_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X8821 _0769_ a_4892_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8822 a_10034_15823# a_9595_15829# a_9949_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8823 a_11425_13353# _0501_ a_11509_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8824 a_14160_27907# cal_lut\[92\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X8825 vccd1 a_9021_29575# net71 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8827 a_8951_25321# _0713_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8828 a_5418_3829# a_5250_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X8829 a_11797_25071# _0706_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8831 vssd1 _0344_ a_24315_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8833 _0290_ a_17875_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8834 _0140_ a_2971_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8835 vccd1 cal_lut\[167\] a_18659_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X8836 a_5307_29789# a_4609_29423# a_5050_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8837 vccd1 net28 a_8951_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8839 vssd1 net41 a_7387_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8840 _0111_ a_18519_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8841 vccd1 _0508_ a_23151_10955# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8842 a_14821_29423# a_14655_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8845 a_19100_22351# _0469_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X8846 vssd1 a_1551_19605# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8847 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2879_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X8848 vssd1 a_20775_5639# _0585_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X8849 _0054_ a_21463_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8850 a_6519_21495# _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X8851 a_7239_17999# a_6541_18005# a_6982_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X8852 a_12311_11079# a_12407_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8853 a_9765_6727# cal_lut\[127\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X8854 a_21725_21807# _0030_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8855 vccd1 a_22403_16635# a_22319_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8856 a_25594_5220# a_25394_5065# a_25743_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8857 vssd1 a_7975_18909# a_8146_18796# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8858 vccd1 a_26479_16042# _0072_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8859 a_12310_10615# _0652_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X8860 vccd1 a_15262_23413# a_15189_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8861 vccd1 a_8695_3829# a_8611_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8862 a_14651_6031# a_14471_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8863 vccd1 a_18942_13621# a_18869_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8864 a_15703_2767# a_14839_2773# a_15446_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8865 _0434_ net7 a_2489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8866 _0364_ a_16859_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8867 vssd1 net43 a_21371_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8868 vssd1 a_9933_19061# _0630_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X8869 _0368_ a_9131_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8870 a_20039_2223# a_19819_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8871 vssd1 a_11609_21379# a_11715_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8872 a_17329_5487# cal_lut\[137\] a_17257_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8873 vssd1 _0481_ a_9565_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8875 cal_lut\[46\] a_16423_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8876 _0352_ a_24683_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X8877 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4811_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X8880 vccd1 a_15611_13647# a_15779_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8881 vssd1 _0872_ a_17401_24759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8882 vccd1 a_12467_3579# a_12383_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8883 a_10129_7125# a_9963_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8885 a_10839_15444# _0661_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8886 _0324_ a_5359_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8887 vccd1 a_6055_10602# _0188_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8888 a_16373_13077# _0604_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X8890 _0584_ a_20175_5056# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X8892 vccd1 a_9650_6005# a_9577_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8893 _0835_ a_4187_28918# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X8894 vccd1 a_2023_19319# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8895 a_10379_6740# _0304_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8896 a_21897_12533# _0456_ a_22054_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X8898 vccd1 cal_lut\[17\] a_17168_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8899 a_9671_26481# ctr\[7\] a_9559_26481# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.131 ps=1.05 w=0.64 l=0.15
X8900 a_12042_3423# a_11874_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8901 vccd1 _0371_ a_14379_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8904 vssd1 a_28031_12559# a_28199_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8905 a_11931_15645# a_11233_15279# a_11674_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8906 a_20066_2589# a_19819_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8908 vssd1 _0717_ a_9673_23047# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8909 vccd1 a_17565_13621# _0596_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8910 vccd1 a_23167_26935# cal_lut\[57\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8911 vccd1 a_4066_7396# a_3995_7497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X8912 a_17312_12879# cal_lut\[17\] a_16737_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8913 ctr\[8\] a_5199_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8914 a_1917_19631# net22 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8915 vssd1 a_15446_2741# a_15404_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8916 a_25755_11989# net36 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8917 vssd1 dbg_result[5] _0592_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8918 vssd1 a_18539_26427# a_18497_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8919 _0665_ _0664_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8920 vssd1 cal_lut\[108\] a_20676_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8921 _0495_ a_13714_19407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8922 a_12057_15279# a_11067_15279# a_11931_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8923 a_24045_15279# cal_lut\[69\] a_23973_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8924 a_20676_5059# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8925 vssd1 a_22219_6843# a_22177_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8926 a_23102_27613# a_22855_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X8927 a_9184_20871# _0592_ a_9326_21046# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X8928 dbg_result[3] a_7410_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X8929 vssd1 _0014_ a_24653_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X8931 a_6403_11293# a_5621_10927# a_6319_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8933 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8934 _0414_ a_2419_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8935 vccd1 a_20690_18517# _0452_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X8937 a_10685_28335# _0197_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8938 vssd1 cal_lut\[87\] a_21872_25731# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8939 _0360_ a_25875_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8940 vccd1 a_25203_10901# a_25210_11201# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8941 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8942 a_9131_13647# a_8951_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8943 a_11471_5853# a_10773_5487# a_11214_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8944 vssd1 dbg_result[1] a_14103_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X8945 a_15163_9527# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8946 ctr\[1\] a_2439_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8947 vccd1 net44 a_20083_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8948 vssd1 _0447_ _0448_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8950 a_16845_26703# cal_lut\[43\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8951 a_8105_1685# a_7939_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8953 a_18313_2057# a_17323_1685# a_18187_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8954 a_3969_12559# _0203_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8955 a_27839_9117# a_27057_8751# a_27755_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8956 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8958 a_5709_6409# a_4719_6037# a_5583_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8959 cal_lut\[87\] a_25439_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8961 a_26983_10383# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8962 ctr\[1\] a_2439_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8963 a_14655_18115# _0442_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X8964 vccd1 _0714_ a_8055_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8965 a_17762_25437# a_17323_25071# a_17677_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8966 a_25191_19631# a_24971_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X8968 a_19793_26703# _0052_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8969 vccd1 a_20947_21263# a_21115_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8970 _0345_ a_24771_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X8971 vccd1 net73 _0403_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8972 a_16220_5737# cal_lut\[149\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X8973 a_17302_17999# a_17029_18005# a_17217_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8974 a_15795_17821# a_15097_17455# a_15538_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8975 a_26830_17705# _0246_ a_26748_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8976 _0342_ a_20815_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8977 a_15469_20407# cal_lut\[34\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X8978 a_27732_17455# a_27333_17455# a_27606_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8979 _0197_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8980 a_23457_3145# a_22903_2985# a_23110_3044# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X8981 vssd1 a_20947_21263# a_21115_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8982 vccd1 _0460_ a_10229_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8983 _0378_ a_12351_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X8984 a_15795_28879# a_14931_28885# a_15538_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X8985 _0460_ a_20451_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8987 vccd1 cal_lut\[150\] a_18975_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8989 a_19421_24533# a_19255_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8990 vccd1 net77 a_4893_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8991 a_3062_23983# _0823_ a_2563_23957# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X8992 vssd1 a_26394_6687# a_26352_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8993 vccd1 a_13997_28023# _0271_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X8994 a_4143_17999# _0421_ a_3785_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8995 _0867_ a_20400_15939# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
R22 vssd1 net56 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8996 a_13717_26709# a_13551_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8997 a_2489_8181# temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8998 a_2887_25615# _0414_ _0746_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8999 a_22695_23439# a_21831_23445# a_22438_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9000 a_22983_15431# _0508_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X9001 a_6265_5487# a_6099_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9002 vccd1 a_6607_9514# _0139_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9005 a_6963_5853# a_6099_5487# a_6706_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9006 a_13173_9001# _0573_ a_13091_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9007 a_15465_28879# a_14931_28885# a_15370_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9008 vccd1 a_10627_15797# a_10543_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9010 vccd1 _0481_ a_16771_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9011 a_2401_11471# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X9012 vssd1 net2 a_6927_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X9013 vccd1 _0812_ a_5487_29217# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X9014 a_1673_16911# net6 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9015 _0839_ a_4167_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9016 vssd1 a_9155_14709# a_9113_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9017 a_28031_12559# a_27167_12565# a_27774_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9018 a_18693_22895# _0454_ a_18611_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9019 a_7368_18377# a_6375_18005# a_7239_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X9020 a_22895_16519# cal_lut\[25\] a_23021_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X9021 a_24125_7485# a_23855_7119# a_24035_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X9022 a_1764_21807# ctr\[4\] a_1461_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X9024 a_19496_13353# cal_lut\[18\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X9025 a_26904_21807# a_26505_21807# a_26778_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9026 a_15208_23145# cal_lut\[51\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X9027 vssd1 net12 a_10055_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9028 a_22365_23439# a_21831_23445# a_22270_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9029 vccd1 a_25007_5175# cal_lut\[161\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9031 a_4984_25615# _0744_ a_4811_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X9032 a_14986_5599# a_14818_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9033 vccd1 a_2000_29111# a_1951_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X9034 a_17871_27613# a_17691_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9035 vccd1 net22 a_1963_21365# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X9036 a_10551_13469# a_9687_13103# a_10294_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9037 vccd1 a_17159_27515# a_17075_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9038 a_10233_22895# _0675_ a_10137_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X9040 vssd1 _0281_ a_18335_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9041 vccd1 cal_lut\[72\] a_26094_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X9043 a_8544_17429# net4 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X9044 a_8377_10927# a_7387_10927# a_8251_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9045 vssd1 a_8845_28023# _0408_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X9046 a_10331_20969# _0670_ a_10413_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X9047 a_14986_5599# a_14818_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9048 a_15023_8751# cal_lut\[132\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9049 a_20966_19743# a_20798_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9050 _0755_ a_3891_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9051 a_22871_14735# a_22089_14741# a_22787_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9052 a_25941_5321# a_25387_5161# a_25594_5220# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9055 vssd1 net11 a_8483_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X9056 vccd1 cal_lut\[117\] a_19343_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9057 _0476_ a_23763_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X9058 vccd1 a_25439_7093# a_25355_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9060 a_9509_28157# dec1.i_ones a_9437_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9061 vccd1 cal_lut\[90\] a_17871_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9062 a_10562_19319# _0628_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X9063 vssd1 a_15262_27765# a_15220_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9064 a_13997_3855# _0131_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9065 a_19065_2045# a_18795_1679# a_18975_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X9066 a_10129_1685# a_9963_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9067 vccd1 _0500_ a_11509_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X9068 _0399_ net76 a_7013_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9070 cal_lut\[140\] a_6947_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9071 cal_lut\[141\] a_4831_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9072 a_6633_26703# a_6397_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X9073 a_17669_9673# a_16679_9301# a_17543_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9074 vssd1 a_4789_11703# net75 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X9075 a_8527_3855# a_7829_3861# a_8270_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9076 a_17919_3073# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X9077 a_19890_2197# a_19690_2497# a_20039_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9078 a_10360_10383# _0494_ a_10258_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X9079 a_2355_12559# a_1573_12565# a_2271_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9080 vssd1 cal_lut\[174\] a_25965_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9081 vssd1 _0467_ a_17661_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9082 a_12870_13215# a_12702_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9083 vccd1 a_9595_26703# a_9947_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.229 ps=1.36 w=0.64 l=0.15
X9084 _0779_ _0432_ a_5915_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9085 vssd1 _0279_ a_14287_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9086 a_12161_25321# _0708_ _0729_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9087 vssd1 a_14675_3829# a_14633_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R23 temp1.capload\[12\].cap_52.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9088 vssd1 a_6982_12127# a_6940_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9089 a_9000_19783# _0703_ a_9142_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9090 a_8951_13647# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9091 a_3327_25935# ctr\[3\] _0746_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X9092 a_25401_17455# a_25235_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9093 vccd1 net43 a_21371_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9094 a_24835_19605# net43 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9095 cal_lut\[151\] a_20931_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9096 vssd1 net31 a_16863_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9097 vccd1 cal_lut\[24\] a_20296_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X9098 vccd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9099 vssd1 _0247_ a_26063_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9101 vccd1 a_23875_7931# a_23791_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9102 _0691_ a_16679_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X9103 vccd1 a_3081_28309# a_3111_28662# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9104 a_14637_8029# a_14103_7663# a_14542_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9105 a_22926_27221# a_22719_27221# a_23102_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9106 net39 a_3155_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X9107 a_4495_21495# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X9108 a_20893_19997# a_20359_19631# a_20798_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9109 vssd1 _0354_ a_26155_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9110 _0316_ a_10108_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X9111 vssd1 a_3325_8903# _0323_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X9114 a_26663_13103# a_26443_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9115 a_8951_25321# _0721_ _0748_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.175 ps=1.35 w=1 l=0.15
X9116 _0032_ a_24591_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9117 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2043_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X9118 vccd1 a_3851_15253# _0198_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X9119 a_18107_7338# _0293_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9120 _0652_ a_11343_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X9121 a_2576_29673# a_2327_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X9122 vccd1 _0838_ a_13459_22359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X9124 vccd1 _0557_ _0819_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9125 vssd1 a_28031_11471# a_28199_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9126 _0804_ _0410_ a_2413_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9127 a_10402_7119# a_9963_7125# a_10317_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9128 vccd1 net23 a_8583_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9129 vccd1 clknet_0__0380_ a_8390_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9130 a_24793_19997# a_24455_19783# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X9134 _0868_ a_23759_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X9135 vccd1 cal_lut\[87\] a_21954_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X9136 vssd1 a_7527_15444# _0036_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9137 a_12797_13469# a_12263_13103# a_12702_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9139 a_20119_28701# a_19255_28335# a_19862_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9140 a_19433_4221# a_19163_3855# a_19343_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X9141 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9142 vccd1 a_7631_17171# _0425_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9143 net14 a_10239_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X9144 vssd1 _0421_ a_2742_18082# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X9145 dbg_result[1] a_6674_16620# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X9146 a_8999_7828# _0303_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9147 a_11243_30511# net13 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X9148 vssd1 a_23811_4564# _0115_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9149 vccd1 a_22503_24135# _0685_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X9151 a_22461_13103# _0013_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9153 ctr\[11\] a_8419_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9154 vccd1 cal_lut\[32\] a_24679_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9155 vccd1 _0836_ a_3370_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X9156 a_12920_27247# a_12521_27247# a_12794_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9157 _0438_ a_13459_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9158 a_7751_13647# a_7571_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9159 vccd1 _0216_ a_15299_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X9160 a_18878_9572# a_18671_9513# a_19054_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X9162 vssd1 a_11639_14459# a_11597_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9163 a_20661_8573# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X9164 a_7527_15444# _0880_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9166 a_11789_3311# _0129_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9167 vccd1 _0630_ _0631_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X9168 vssd1 a_18107_8439# _0607_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9169 a_4491_13879# ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9170 a_11674_15391# a_11506_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9171 a_4732_28169# a_4333_27797# a_4606_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9172 a_2778_24527# temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9173 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X9174 _0383_ a_6979_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9176 vccd1 cal_lut\[19\] a_7751_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9178 a_19061_21629# _0453_ a_18979_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9179 vccd1 _0446_ a_14417_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X9180 a_24455_19783# a_24551_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9181 a_12686_1653# a_12518_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9183 vccd1 a_25755_11989# a_25762_12289# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9184 _0797_ _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X9185 a_5326_6005# a_5158_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9186 a_18187_25437# a_17323_25071# a_17930_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9187 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9188 _0418_ a_2327_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9189 a_12626_10927# a_12311_11079# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9190 a_7716_22325# _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X9191 io_out[2] a_2511_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9193 a_21555_18909# _0442_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9194 a_18685_16917# a_18519_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9195 cal_lut\[134\] a_7315_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9196 a_14778_14441# _0851_ a_14696_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9197 vssd1 a_10659_7637# net26 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X9198 vccd1 a_15538_28853# a_15465_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9199 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9200 a_20943_12043# _0505_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X9202 vccd1 net23 a_9043_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9203 a_14151_4564# _0313_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9204 vssd1 _0711_ a_11547_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9205 vssd1 net24 a_4535_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9206 net28 a_6007_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9208 vccd1 a_16373_13077# _0609_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X9209 vssd1 cal_lut\[181\] a_9221_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9210 vssd1 a_9650_6005# a_9608_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9211 a_13714_19407# a_13459_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.312 ps=2.12 w=1 l=0.15
X9212 _0434_ _0422_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9213 cal_lut\[29\] a_19551_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9215 vccd1 cal_lut\[59\] a_20022_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X9216 vccd1 a_22438_23413# a_22365_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9217 vssd1 a_18475_5639# _0615_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9218 cal_lut\[126\] a_15503_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9220 vssd1 _0422_ _0741_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9221 vccd1 cal_lut\[142\] a_4163_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9222 vccd1 _0239_ a_25787_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9223 a_6979_19061# _0439_ a_7188_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X9224 a_5728_24847# _0794_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X9225 _0708_ _0681_ a_11142_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X9226 a_13809_3861# a_13643_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9227 vssd1 cal_lut\[82\] a_17041_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9228 vccd1 _0423_ a_2447_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9229 a_15325_9661# net20 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X9230 vssd1 _0808_ a_3877_11703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9231 a_11756_22671# _0674_ a_11684_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0683 ps=0.86 w=0.65 l=0.15
X9232 a_22523_5175# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X9234 a_15494_19319# dbg_result[1] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X9235 vssd1 _0025_ a_24469_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9236 a_17560_4917# _0440_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X9237 vccd1 net38 a_19255_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9238 _0814_ a_5915_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9239 a_21166_10205# a_20893_9839# a_21081_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9240 a_4897_27247# _0812_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9241 vccd1 net67 a_3882_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9243 a_28031_11471# a_27167_11477# a_27774_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
R24 vccd1 temp1.capload\[7\].cap_62.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9244 vccd1 cal_lut\[173\] a_17187_13255# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X9245 a_7025_21041# _0735_ a_6516_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X9246 a_15093_1135# a_14103_1135# a_14967_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9247 a_5341_17429# clknet_0_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9248 cal_lut\[105\] a_21759_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9249 net4 a_1407_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X9250 a_25757_10927# a_25210_11201# a_25410_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9251 a_8544_17429# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X9253 a_6823_14735# a_6541_14741# a_6729_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X9254 _0853_ a_17732_14441# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X9256 vssd1 a_18907_12533# a_18865_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9259 vssd1 _0745_ a_2023_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X9260 vccd1 a_20775_14967# _0527_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9261 vssd1 a_13942_20149# _0485_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9262 a_21879_6250# _0342_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9263 vssd1 _0467_ a_12693_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9264 a_19956_22057# cal_lut\[64\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X9265 vccd1 net56 temp1.capload\[1\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9266 vssd1 a_4912_8439# net24 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X9267 a_18318_27791# a_18071_28169# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9268 vssd1 ctr\[8\] _0410_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9269 vccd1 a_2209_25589# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X9270 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9271 vccd1 a_4771_4917# _0320_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X9273 vccd1 a_15871_2741# a_15787_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9274 vccd1 _0505_ a_19071_11584# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9275 a_20237_2223# a_19683_2197# a_19890_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9276 a_3985_16189# net69 a_3885_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X9277 a_20194_13647# _0532_ a_20114_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9278 vccd1 _0362_ a_25419_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9279 vccd1 a_20966_19743# a_20893_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9280 a_1683_17455# net5 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9281 vccd1 _0609_ a_11895_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9282 a_22615_19631# a_22395_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X9283 a_11545_9117# a_11207_8903# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X9284 vccd1 a_17498_29397# a_17427_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9286 a_7571_13647# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9287 a_19694_28701# a_19255_28335# a_19609_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9288 vssd1 temp1.dac_vout_notouch_ a_3607_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X9289 vccd1 a_17560_4917# _0441_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9290 a_22481_9839# cal_lut\[177\] a_22409_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9291 a_4238_10205# a_3799_9839# a_4153_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9292 vccd1 _0841_ a_23027_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X9293 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_2576_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X9294 vccd1 _0818_ a_5545_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X9295 _0672_ a_10372_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X9296 vssd1 a_12391_7119# a_12559_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9297 _0176_ a_25419_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9298 vccd1 a_22971_13469# a_23139_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9300 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9301 a_20641_16367# cal_lut\[30\] a_20569_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9302 vccd1 net25 a_11435_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9303 a_13353_12559# _0191_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9304 vssd1 a_20287_24501# a_20245_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9305 a_14896_15529# cal_lut\[35\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X9306 a_22553_25071# _0085_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9307 a_16105_4233# a_15115_3861# a_15979_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9308 a_20237_2223# a_19690_2497# a_19890_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9309 a_10851_11079# _0495_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X9310 vccd1 a_15687_27765# a_15603_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9311 vssd1 _0755_ a_5444_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9312 a_18107_8439# _0514_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9313 a_14747_27497# _0487_ a_14829_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9314 _0219_ a_15479_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9315 vccd1 net45 a_15391_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9316 a_15370_17821# a_15097_17455# a_15285_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9317 a_5250_9295# a_4977_9301# a_5165_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9318 vssd1 cal_lut\[176\] a_25137_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9319 a_13512_13621# _0575_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X9320 a_19054_9295# a_18807_9673# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X9321 a_6182_22895# clknet_0_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9322 a_16189_18365# cal_lut\[95\] a_16117_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9323 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9324 vssd1 a_20874_27765# a_20832_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9325 a_4174_25654# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X9326 vssd1 a_3155_16911# _0421_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X9327 a_17894_13647# _0594_ a_17814_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9328 a_26137_18543# a_25971_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9329 a_10528_7497# a_10129_7125# a_10402_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9330 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X9331 a_27847_17999# a_27149_18005# a_27590_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9332 _0858_ a_14604_13353# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X9333 a_3851_15253# net68 a_4189_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.12 ps=1.02 w=0.65 l=0.15
X9334 a_20893_4399# a_20727_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9335 a_25389_13103# a_24835_13077# a_25042_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9336 _0427_ _0426_ a_4443_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9337 a_10141_9615# cal_lut\[121\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X9338 a_18041_12565# a_17875_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9339 a_12978_23261# a_12539_22895# a_12893_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9340 a_19467_16911# a_18685_16917# a_19383_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9341 vccd1 net6 a_1683_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9342 vccd1 a_1743_18259# _0422_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X9343 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6184_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X9344 _0092_ a_13275_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9345 a_4714_23483# _0797_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X9346 a_3882_22895# clknet_0_temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9347 _0071_ a_27351_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9348 vssd1 net25 a_9963_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9349 vccd1 a_1673_22351# a_1773_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9350 a_14163_8903# _0440_ a_14337_8779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X9351 vccd1 net42 a_25235_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9352 vssd1 net72 _0397_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9353 vccd1 a_6522_29535# a_6449_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9354 a_23483_18909# a_23303_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9355 a_16373_13077# _0608_ a_16753_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X9356 a_15193_2767# _0179_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9357 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd _0773_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9359 vccd1 a_6955_23671# _0753_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X9360 vssd1 a_22891_20871# _0636_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9361 vssd1 a_7718_18679# a_7656_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X9362 a_5141_21781# _0432_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X9363 vssd1 a_10839_15444# net12 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9364 a_14345_9269# _0562_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9366 _0237_ a_12723_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9367 a_12475_7119# a_11693_7125# a_12391_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9369 vccd1 a_5475_29691# a_5391_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9370 a_17037_20719# _0531_ a_16955_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9371 a_20245_5487# a_19255_5487# a_20119_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9372 a_15170_10357# a_15002_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9373 _0172_ a_27351_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9374 a_4521_27791# _0207_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9375 vccd1 a_11765_17973# _0589_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X9376 _0182_ a_10055_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9377 a_17930_25183# a_17762_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9378 a_16679_24527# _0484_ a_16761_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9379 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9381 a_16566_27613# a_16127_27247# a_16481_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9382 vssd1 net30 a_12171_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9384 vccd1 a_22843_9295# _0451_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9385 _0649_ a_10699_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9386 a_21954_24643# _0260_ a_21872_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9387 vssd1 _0724_ a_7523_24833# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9388 a_19793_28879# _0048_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9389 vssd1 clknet_0_temp1.i_precharge_n a_1753_26133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9390 vccd1 a_9375_29397# a_9117_29397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X9391 _0428_ _0411_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9392 a_9831_24501# _0720_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X9393 a_6503_16733# a_5639_16367# a_6246_16503# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9395 a_15722_12533# a_15554_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9396 a_12249_17455# _0005_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9398 vccd1 _0875_ a_23763_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9400 vccd1 cal_lut\[159\] a_23943_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9401 vssd1 a_8419_13371# a_8377_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9402 a_13997_28023# cal_lut\[92\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X9403 vssd1 temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X9404 a_16481_21807# _0041_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9405 _0098_ a_12263_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9406 vssd1 a_6519_21495# _0780_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X9408 a_18107_8439# _0514_ a_18341_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9409 a_18751_23671# _0459_ a_18985_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9410 vccd1 a_12778_3829# a_12705_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9411 _0137_ a_4443_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9412 _0744_ a_1736_18517# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X9413 vccd1 _0290_ a_18335_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X9414 _0124_ a_13183_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9415 a_22365_25071# a_22199_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9416 a_1867_23759# _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9417 a_6982_14709# a_6823_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X9418 vssd1 net25 a_14839_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9420 vccd1 _0483_ a_9043_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X9421 a_1921_11989# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X9422 a_15554_12559# a_15281_12565# a_15469_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9423 a_13219_27613# a_12521_27247# a_12962_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9424 a_21739_27613# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9425 vssd1 cal_lut\[31\] a_23481_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9426 a_20775_14967# _0459_ a_21009_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9427 a_21626_6941# a_21353_6575# a_21541_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9429 a_27333_17455# a_27167_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9430 a_15943_12015# cal_lut\[191\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9432 a_23053_20719# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X9433 a_10968_27247# a_10589_27247# a_10871_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X9434 vccd1 net22 a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9435 vssd1 clknet_1_0__leaf_io_in[0] a_1959_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9436 a_5483_8029# a_4701_7663# a_5399_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9437 vccd1 _0352_ a_27351_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X9438 a_13997_28023# _0260_ a_14160_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9439 vssd1 a_22926_27221# a_22855_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9440 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9441 a_15974_15823# _0542_ a_15725_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X9442 a_26141_6575# _0161_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9443 _0501_ a_19977_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X9444 a_21166_10205# a_20727_9839# a_21081_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9445 a_9563_28487# _0815_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X9446 a_23815_12791# a_24106_12681# a_24057_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9448 vccd1 _0557_ a_10715_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9449 a_11421_15279# _0004_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9450 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9451 _0863_ a_13144_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X9452 a_5517_10761# a_4970_10505# a_5170_10660# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9453 vssd1 a_5105_25045# a_5039_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X9454 a_23077_21835# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X9455 a_4153_8751# _0140_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9456 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9457 a_24938_15823# a_24665_15829# a_24853_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9458 _0329_ a_10051_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9459 _0369_ a_9591_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9460 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9461 a_7607_6031# a_6743_6037# a_7350_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9463 a_6909_12381# a_6375_12015# a_6814_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9464 vssd1 net8 a_10515_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9465 vccd1 ctr\[5\] a_5555_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9466 vccd1 a_17935_28009# a_17942_27913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9467 vccd1 _0438_ _0439_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9468 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9470 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9471 _0348_ a_24035_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9472 vccd1 net30 a_12999_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9473 vssd1 a_24827_24501# _0238_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X9474 a_6939_22351# _0787_ a_6737_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9475 vssd1 a_16734_21919# a_16692_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9476 vccd1 _0411_ a_4091_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X9478 a_10943_23671# _0679_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X9479 vssd1 cal_lut\[29\] a_19756_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9480 a_7182_6031# a_6743_6037# a_7097_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9481 vssd1 a_2566_15797# a_2524_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9482 a_21883_1109# a_22059_1109# a_22011_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X9483 vssd1 a_14158_26677# a_14116_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9485 _0725_ a_8971_22895# a_9209_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X9486 _0283_ a_13459_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X9487 _0288_ a_20676_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X9489 vccd1 _0483_ a_15943_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9490 a_3056_29199# temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X9491 vssd1 cal_lut\[25\] a_23849_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9493 vssd1 _0839_ _0196_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9494 vssd1 a_2933_14709# _0202_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9495 vssd1 a_25014_8863# a_24972_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9496 a_11302_16519# _0609_ a_11439_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9498 a_20775_5639# _0441_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9499 cal_lut\[96\] a_15963_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9500 a_22619_15253# net38 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X9501 a_18545_5309# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X9502 vccd1 a_20471_26677# a_20387_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9503 a_21879_19783# a_21975_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9504 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd a_1584_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X9505 a_19303_23047# _0454_ a_19537_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9506 a_4364_9839# a_3965_9839# a_4238_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9508 a_4032_25847# ctr\[1\] a_4174_25654# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X9509 vssd1 a_22625_17973# _0643_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X9510 a_9117_8207# a_8583_8213# a_9022_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9511 _0842_ a_8303_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9512 a_6522_29535# a_6354_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9513 a_20775_26311# a_20871_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X9514 cal_lut\[30\] a_21023_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9515 a_22438_1653# a_22270_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9516 a_15427_10383# a_14729_10389# a_15170_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9517 vccd1 a_24243_19061# a_24159_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9518 vccd1 a_21362_26133# a_21291_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9519 vccd1 a_19303_23047# _0619_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X9521 a_10839_19958# _0629_ a_10380_19783# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X9522 a_8059_18909# a_7277_18543# a_7975_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X9523 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9525 a_4238_9117# a_3799_8751# a_4153_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9526 vssd1 _0211_ a_10025_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X9527 a_25011_21781# a_25302_22081# a_25253_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9528 a_6354_9117# a_5915_8751# a_6269_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9529 _0724_ a_9372_24135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X9530 vccd1 net10 a_7847_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X9531 a_28115_10205# a_27333_9839# a_28031_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9532 a_19961_22895# cal_lut\[90\] a_19889_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9533 a_15979_12559# a_15281_12565# a_15722_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9534 vccd1 a_1945_15431# _0388_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X9535 vssd1 a_25927_10602# _0169_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9536 a_12679_28010# _0847_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9537 vccd1 _0755_ a_5915_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X9538 vccd1 _0483_ a_10607_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9539 a_15554_12559# a_15115_12565# a_15469_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9540 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9541 vssd1 _0697_ a_9043_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9542 vssd1 a_7410_17973# a_7368_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9543 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9544 vccd1 ctr\[12\] a_8329_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9545 _0869_ a_23483_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X9546 vccd1 a_14273_15431# _0880_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X9547 a_16155_22923# _0464_ a_16069_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X9548 a_26735_6941# a_25953_6575# a_26651_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9549 vssd1 _0259_ a_17323_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9550 _0544_ a_15943_7232# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X9552 a_10699_24233# _0707_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9553 net40 a_12723_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X9554 vssd1 ctr\[1\] a_2685_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9555 _0230_ a_21919_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X9556 a_23205_17455# _0473_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X9558 vssd1 net42 a_23211_19093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9560 vccd1 a_18645_12043# _0502_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X9561 a_3575_7351# a_3866_7241# a_3817_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9562 a_8055_25321# _0721_ a_7755_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X9563 _0001_ a_7387_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9564 a_23055_23047# cal_lut\[32\] a_23201_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X9565 a_1860_22711# a_1673_22351# a_1773_22467# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X9566 a_12705_3855# a_12171_3861# a_12610_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9567 a_6637_3311# _0133_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9568 _0280_ a_15524_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X9569 vccd1 _0420_ a_1625_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X9570 a_25030_17999# a_24591_18005# a_24945_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9571 a_22695_1679# a_21997_1685# a_22438_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9572 a_8937_8207# _0121_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9573 _0249_ a_26012_15939# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X9574 vssd1 a_25439_24251# a_25397_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9575 a_17197_19777# _0581_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9576 _0680_ _0433_ a_8975_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9577 vccd1 net34 a_23211_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X9578 vccd1 _0706_ a_12265_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9579 _0252_ a_25552_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X9580 a_16737_13621# _0599_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9581 vccd1 _0377_ a_6099_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9582 a_16803_22689# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X9583 a_14365_24527# _0093_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9585 a_3852_14165# ctr\[3\] a_3981_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9586 cal_lut\[147\] a_10995_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9587 vssd1 _0462_ a_22813_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9588 a_12521_27247# a_12355_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9590 _0664_ a_10596_17705# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9591 vccd1 a_6246_16503# a_6180_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X9592 vssd1 a_26307_13077# a_26314_13377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9593 vccd1 net81 a_14287_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9594 a_24485_17607# _0246_ a_24648_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9595 cal_lut\[170\] a_26635_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9596 vssd1 a_9429_19605# a_9363_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X9597 _0190_ a_6099_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9598 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9600 a_13028_7913# _0570_ a_12926_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X9601 vssd1 a_5779_8426# _0141_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9603 a_4771_20871# _0438_ a_4897_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X9604 vccd1 a_17314_4132# a_17243_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X9605 a_15009_23439# _0094_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9606 vccd1 _0450_ a_22659_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9607 vssd1 _0569_ a_13091_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X9608 vssd1 _0340_ a_19807_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9610 _0737_ a_3799_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9611 a_21879_6250# _0342_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9612 _0293_ a_16996_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X9613 vssd1 _0503_ a_8951_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9614 a_19694_28701# a_19421_28335# a_19609_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9615 vssd1 a_8268_24501# _0722_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X9616 a_15821_20719# cal_lut\[40\] a_15749_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9617 a_1743_18259# net5 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X9618 a_20119_15645# a_19421_15279# a_19862_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9619 a_11759_4564# _0311_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9620 a_24761_25071# _0086_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9621 cal_lut\[101\] a_15595_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9622 vssd1 cal_lut\[72\] a_26012_15939# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9624 a_2773_9991# _0836_ a_2936_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9625 _0075_ a_26063_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9626 vccd1 a_9815_1501# a_9983_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9627 a_16390_5487# cal_lut\[149\] a_16309_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X9628 vccd1 a_7071_25045# _0735_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9629 a_17682_16100# a_17482_15945# a_17831_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X9630 a_27333_15829# a_27167_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9631 _0476_ a_23763_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9632 _0391_ _0389_ a_2401_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9633 a_5060_31055# a_4811_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X9634 a_8951_28335# _0407_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X9635 a_19862_4511# a_19694_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9636 a_11509_13353# cal_lut\[21\] a_11425_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9637 a_8665_28585# _0815_ _0407_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9638 a_4774_27765# a_4606_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9639 vssd1 cal_lut\[159\] a_24033_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9640 a_21292_9839# a_20893_9839# a_21166_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9641 a_15535_24501# a_15711_24833# a_15663_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X9642 cal_lut\[180\] a_15871_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9643 a_19881_9301# a_19715_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9645 _0794_ _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X9646 a_18765_22895# cal_lut\[83\] a_18693_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9647 vccd1 a_16055_19899# a_15971_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9648 a_19862_5599# a_19694_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9649 _0718_ _0716_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9650 _0845_ a_12856_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X9651 vssd1 _0810_ a_5179_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X9652 a_9397_6031# _0127_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9653 a_16636_5737# _0615_ a_16534_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X9654 cal_lut\[170\] a_26635_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9655 vssd1 _0730_ a_11797_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X9656 vccd1 a_2439_14709# a_2355_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9657 a_19333_13255# _0851_ a_19496_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9658 a_5630_21583# _0755_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X9659 vccd1 a_27590_17973# a_27517_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9661 a_1573_14741# a_1407_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9662 vssd1 _0690_ a_16679_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9663 vssd1 a_25011_14709# _0244_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X9664 a_2309_14191# a_2143_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9666 vssd1 dec1.i_ones _0720_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9667 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X9668 vccd1 ctr\[10\] a_7133_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9669 a_18647_28879# a_17949_28885# a_18390_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9670 a_17095_16055# a_17191_16055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9671 vccd1 a_8723_17130# _0002_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9673 _0510_ a_22875_9867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X9674 a_22649_23983# _0468_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X9675 vssd1 a_10551_11471# a_10719_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9676 a_9853_11477# a_9687_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9677 a_10938_28471# a_10779_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X9678 vssd1 a_9372_24135# _0724_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X9679 a_5725_22351# ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9680 a_9184_20871# _0626_ a_9326_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9682 a_7308_6409# a_6909_6037# a_7182_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9683 temp1.capload\[12\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9684 a_21334_11039# a_21166_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9685 a_6699_13268# _0860_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9686 vssd1 a_25962_11989# a_25891_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X9687 _0801_ _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9688 vccd1 net26 a_14471_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9689 vssd1 _0586_ a_17094_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X9690 _0472_ a_14770_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9691 a_9542_4649# cal_lut\[182\] a_9385_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9692 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9693 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9695 a_2398_15823# a_1959_15829# a_2313_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9697 a_11723_8751# a_11587_8725# a_11303_8725# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9698 a_23426_4649# _0283_ a_23344_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9699 a_9034_6825# _0498_ a_9034_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X9700 vssd1 _0328_ a_7571_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9701 vccd1 a_7775_10357# a_7691_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9702 a_25047_11471# a_24867_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9703 vssd1 _0418_ a_5995_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0894 ps=0.925 w=0.65 l=0.15
X9704 net6 a_1407_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9705 vssd1 a_4406_9951# a_4364_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9706 a_2518_30006# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X9707 a_16566_27613# a_16293_27247# a_16481_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9708 a_2489_17455# net7 _0434_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9709 vccd1 _0706_ a_12161_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9710 vssd1 cal_lut\[84\] a_20997_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9711 _0086_ a_23763_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9712 _0260_ a_13367_10391# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X9714 vssd1 _0481_ a_10853_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9715 a_25125_17999# a_24591_18005# a_25030_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9716 vccd1 a_1407_10383# net4 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9718 cal_lut\[43\] a_17159_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9719 a_17129_22895# _0500_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X9720 a_21725_16367# _0024_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9721 a_8377_29423# a_7387_29423# a_8251_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9722 a_19225_9673# a_18678_9417# a_18878_9572# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X9723 vccd1 _0412_ a_2139_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X9724 vssd1 _0600_ a_16373_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9725 vssd1 a_5843_13371# a_5801_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9726 vccd1 a_11471_5853# a_11639_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9727 a_4364_8751# a_3965_8751# a_4238_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9728 a_6480_8751# a_6081_8751# a_6354_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9729 io_out[0] a_2023_19319# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.5 ps=3 w=1 l=0.15
X9730 vssd1 _0442_ a_19715_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X9731 cal_lut\[184\] a_13111_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9732 vccd1 a_25271_9117# a_25439_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9733 a_15378_22895# _0646_ a_15624_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X9735 vccd1 a_3479_7351# cal_lut\[142\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9736 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9737 a_17927_4917# _0440_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X9738 vccd1 _0451_ a_10699_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9739 a_1913_28023# _0744_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X9740 vssd1 cal_lut\[162\] a_26609_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9741 vssd1 a_8565_28879# a_8671_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X9742 _0520_ _0433_ a_9135_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9743 a_12943_1679# a_12079_1685# a_12686_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9744 a_5643_22671# _0747_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X9745 a_9043_16733# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9746 vssd1 a_25755_11989# a_25762_12289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9747 a_15519_27791# a_14821_27797# a_15262_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9748 a_15663_24893# cal_lut\[94\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X9749 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9750 a_11142_24233# a_10784_23983# _0708_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9751 a_13146_23007# a_12978_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9752 vssd1 a_13714_19407# _0495_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9753 _0168_ a_26155_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9754 vssd1 a_21897_12533# _0683_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X9755 a_26413_16733# a_25879_16367# a_26318_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9756 a_10953_3311# a_9963_3311# a_10827_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9757 vccd1 _0801_ temp1.dac.vdac_single.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9759 a_15262_23413# a_15094_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9760 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9761 vssd1 _0875_ a_23763_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9764 vccd1 a_2288_17973# _0420_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9765 a_8377_6575# a_7387_6575# a_8251_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9766 a_6319_11293# a_5455_10927# a_6062_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9767 a_9091_29111# a_9187_29111# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9768 a_12455_18793# _0556_ _0557_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9769 _0452_ a_20690_18517# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9770 vccd1 a_1651_14165# _0411_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X9771 vssd1 cal_lut\[63\] a_25505_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9772 a_13823_1679# a_13643_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9773 a_11707_1679# a_11527_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9774 a_6909_12559# a_6375_12565# a_6814_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9775 a_20246_22351# a_19807_22357# a_20161_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9776 a_21683_14557# a_20819_14191# a_21426_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9777 a_20329_5309# cal_lut\[154\] a_20257_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9778 _0137_ a_4443_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9779 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9781 a_1917_19881# _0762_ a_1551_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9782 vccd1 a_21265_7815# _0292_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X9785 vssd1 a_22259_19605# a_22266_19905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9786 _0108_ a_21371_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9787 vccd1 a_2271_12559# a_2439_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9788 vssd1 _0390_ a_6914_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X9789 vssd1 a_7410_14709# dbg_result[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X9790 cal_lut\[134\] a_7315_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9791 a_22270_8207# a_21997_8213# a_22185_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9793 a_12460_17455# a_12061_17455# a_12334_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9794 vccd1 a_11207_8903# cal_lut\[99\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9796 vccd1 _0531_ a_16955_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9797 vssd1 a_12686_1653# a_12644_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9798 vssd1 net34 a_23211_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9799 a_25287_12533# cal_lut\[175\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X9800 vssd1 _0806_ a_2959_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9801 vssd1 a_2939_23047# _0417_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X9802 vccd1 a_25271_25437# a_25439_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9803 a_27583_9514# _0356_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9804 a_2652_28487# _0800_ a_2794_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9805 a_3990_23983# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X9806 a_6541_18005# a_6375_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9807 a_24757_18005# a_24591_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9808 _0810_ a_4843_15307# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X9809 a_15557_27497# cal_lut\[44\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9810 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd _0817_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9811 a_19133_21629# cal_lut\[64\] a_19061_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9812 vccd1 _0168_ a_26677_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9813 a_5675_3855# a_4977_3861# a_5418_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9814 a_10551_11471# a_9687_11477# a_10294_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9815 net19 a_21095_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9816 vssd1 a_15255_28500# _0091_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9817 a_8055_25321# _0714_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9818 a_19838_16617# _0872_ a_19756_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9819 a_21353_14557# a_20819_14191# a_21258_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9820 vccd1 a_17927_4917# _0445_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9821 a_3425_18319# _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9822 vssd1 net38 a_19255_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9823 vssd1 a_4491_13879# _0809_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X9824 a_15715_30186# _0218_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9826 a_3869_11989# clknet_0_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9827 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9828 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9830 vccd1 a_24731_6740# _0163_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9831 a_9767_26159# _0592_ a_9559_26481# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.173 ps=1.25 w=0.42 l=0.15
X9832 a_19399_2197# a_19690_2497# a_19641_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X9833 vssd1 a_17783_21271# _0531_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9835 vccd1 _0420_ a_3615_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9836 a_23489_17455# _0475_ a_23079_17607# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X9837 a_14250_3829# a_14082_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9838 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_5060_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X9839 a_17291_29397# net45 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9840 a_18669_22325# _0618_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9841 vssd1 net44 a_20359_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9844 _0154_ a_19439_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9845 _0749_ _0718_ a_10965_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.105 ps=1.21 w=1 l=0.15
X9846 vccd1 _0097_ a_13245_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9847 vssd1 a_10294_13215# a_10252_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9848 vssd1 net10 a_8299_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X9849 cal_lut\[121\] a_8419_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9850 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9851 vccd1 a_21794_6687# a_21721_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9852 a_8335_11293# a_7553_10927# a_8251_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9853 a_13947_12559# a_13165_12565# a_13863_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9854 vssd1 _0858_ a_14839_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9855 a_9187_29111# a_9471_29097# a_9406_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X9856 a_4077_18793# _0426_ a_3995_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9857 vccd1 net33 a_21831_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9859 a_23273_27247# a_22719_27221# a_22926_27221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X9860 vssd1 a_21334_9951# a_21292_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9862 vssd1 net29 a_12263_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9864 vccd1 _0843_ a_9595_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9865 vssd1 a_19862_15391# a_19820_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9866 a_20905_6575# a_20635_6941# a_20815_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X9868 a_19421_4399# a_19255_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9869 vssd1 a_3852_14165# _0394_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X9871 a_15909_7809# _0545_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9872 vccd1 a_7775_6005# a_7691_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9873 _0016_ a_14839_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9874 vssd1 a_7369_28879# a_7475_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X9875 vccd1 _0486_ a_15208_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X9876 vssd1 a_20966_19743# a_20924_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9877 vssd1 a_28015_17973# a_27973_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9878 vssd1 _0839_ _0192_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9879 a_5284_15113# a_4885_14741# a_5158_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9880 a_11046_5853# a_10607_5487# a_10961_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9882 _0259_ a_16951_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X9883 a_25505_22717# a_25235_22351# a_25415_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X9884 vssd1 a_16727_21482# _0041_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9885 cal_lut\[12\] a_19367_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9888 vccd1 net35 a_17875_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9889 a_4253_19087# _0429_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X9890 a_21975_2741# cal_lut\[153\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X9891 vssd1 _0216_ a_14331_29397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9892 vccd1 a_18815_28853# a_18731_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9893 vssd1 _0251_ a_24315_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9894 vccd1 cal_lut\[84\] a_20907_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9895 a_2953_20719# ctr\[2\] _0419_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X9896 a_19126_16885# a_18958_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9897 vccd1 _0152_ a_23457_3145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X9898 a_22787_14735# a_21923_14741# a_22530_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X9899 cal_lut\[12\] a_19367_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9900 a_2839_27221# _0830_ a_3066_27569# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X9901 a_17033_9295# _0106_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9903 a_10045_9295# _0493_ a_10129_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9904 a_16727_21482# _0214_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9905 vssd1 a_12870_13215# a_12828_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9906 temp1.dac_vout_notouch_ net13 a_11796_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X9907 vccd1 a_25198_17973# a_25125_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9909 a_12539_6144# cal_lut\[130\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9910 vccd1 _0850_ a_24683_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X9911 vccd1 a_15078_7093# a_15005_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9912 a_12995_26525# a_12815_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9913 vccd1 ctr\[7\] a_6397_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9914 a_9129_13103# cal_lut\[20\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X9915 _0467_ a_15370_19407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9916 a_23039_3145# a_22910_2889# a_22619_2999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X9917 a_2000_26935# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X9919 a_14250_3829# a_14082_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9920 a_15002_10383# a_14563_10389# a_14917_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9921 _0740_ _0739_ a_4627_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9922 vssd1 a_12559_7093# a_12517_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9923 vccd1 a_9647_14709# _0256_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X9924 a_22457_14735# a_21923_14741# a_22362_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9925 a_20506_1653# a_20338_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X9928 vccd1 net36 a_25603_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9929 vccd1 a_1735_27765# _0825_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X9930 a_15469_26935# _0260_ a_15632_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9931 a_23055_23047# cal_lut\[62\] a_23201_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9932 _0413_ a_1773_22467# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X9933 vccd1 a_24835_19605# a_24842_19905# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9934 vssd1 net42 a_25235_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9935 a_5173_29199# _0814_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9936 cal_lut\[80\] a_9983_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9938 _0824_ a_2563_23957# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9939 vssd1 _0809_ a_4929_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9940 vssd1 a_4406_8863# a_4364_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X9941 a_14733_15431# _0872_ a_14896_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9942 vssd1 net28 a_7111_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X9943 vccd1 clknet_0__0380_ a_8390_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9944 vccd1 a_26486_16479# a_26413_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9945 vccd1 _0859_ a_17599_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9946 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9568_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X9947 a_7347_24501# _0728_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X9948 a_18913_23805# _0481_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X9949 vccd1 _0759_ a_5507_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X9950 a_22175_5263# cal_lut\[151\] a_22079_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.107 ps=0.98 w=0.65 l=0.15
X9951 vssd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_2409_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9952 _0836_ a_3155_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X9953 vssd1 a_20287_5755# a_20245_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9954 vccd1 a_3155_7663# net39 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9955 a_10911_7119# a_10129_7125# a_10827_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9956 vssd1 _0671_ a_12437_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9959 vccd1 clknet_1_0__leaf__0380_ a_5460_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9960 vssd1 _0295_ a_20727_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9962 vssd1 _0438_ _0455_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X9963 vssd1 a_6791_4074# _0133_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X9964 _0127_ a_8767_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9965 vccd1 net31 a_19899_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9966 a_24941_24349# a_24407_23983# a_24846_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X9968 a_27422_7119# a_27149_7125# a_27337_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9969 cal_lut\[46\] a_16423_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9970 vccd1 _0467_ a_9595_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X9971 a_9907_6031# a_9209_6037# a_9650_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9972 vccd1 _0711_ _0730_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9973 _0017_ a_17599_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X9974 a_19345_20719# _0486_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X9975 vssd1 _0382_ _0193_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9976 a_22711_6549# a_22887_6549# a_22839_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X9978 a_9687_17455# _0519_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X9979 vssd1 a_24485_17607# _0251_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X9980 a_21426_14303# a_21258_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9981 a_6603_11777# _0836_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X9982 a_20345_16911# _0029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X9983 a_4789_11703# a_4885_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X9984 vssd1 a_21591_25437# a_21759_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9985 a_2569_22671# _0414_ a_2485_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X9986 a_19426_20719# _0560_ a_19672_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X9987 vccd1 _0336_ a_22659_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X9988 vccd1 _0495_ a_12539_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X9989 _0421_ a_3155_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X9990 vccd1 a_21426_14303# a_21353_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X9991 a_10317_3311# _0146_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X9993 net3 a_1407_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9994 a_19862_28447# a_19694_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X9995 a_27606_10205# a_27167_9839# a_27521_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9996 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9956_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X9997 vccd1 a_20543_18543# a_20690_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X9998 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9999 vccd1 a_18390_28853# a_18317_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10000 a_5069_8029# a_4535_7663# a_4974_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10001 a_14594_9295# _0564_ a_14345_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10002 vssd1 _0257_ a_10699_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10003 a_19865_13621# _0533_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10005 vccd1 a_20775_27412# _0053_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10006 vccd1 dbg_result[3] a_21721_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X10007 a_27333_17455# a_27167_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10008 a_19789_15645# a_19255_15279# a_19694_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10009 _0312_ a_12535_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X10010 a_21721_6941# a_21187_6575# a_21626_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10011 a_13441_28885# a_13275_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10012 a_7256_21237# _0755_ a_7648_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X10013 vssd1 a_26479_16042# _0072_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10015 a_19283_13647# a_18501_13653# a_19199_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10016 a_5545_23439# _0819_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X10017 a_14417_19881# _0438_ a_14321_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X10018 a_6916_17999# a_6375_18005# a_6823_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X10019 vccd1 a_24455_19783# cal_lut\[28\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10020 a_28057_15279# a_27503_15253# a_27710_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10021 vssd1 a_5687_4564# _0134_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10022 _0616_ a_16127_5056# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10025 cal_lut\[29\] a_19551_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10027 vssd1 a_22051_6941# a_22219_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10028 vssd1 a_22695_27791# a_22863_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10029 vccd1 a_2327_22895# _0418_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10030 a_20871_26133# a_21155_26133# a_21090_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10031 a_8951_12559# _0501_ a_9033_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10032 a_2747_18517# _0423_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X10033 _0080_ a_10699_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10034 vccd1 a_12223_2741# _0330_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10035 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10037 a_24041_10927# _0509_ a_23631_11079# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X10038 vccd1 a_15439_17130# _0095_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10041 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7840_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X10042 a_9595_16367# _0519_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X10043 a_10570_3423# a_10402_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10044 a_4882_29789# a_4609_29423# a_4797_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10045 a_2790_24305# a_2741_24135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X10046 a_15715_5175# _0452_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X10047 vssd1 a_24407_15279# _0246_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X10048 vccd1 a_7255_20871# _0768_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X10050 vccd1 a_2287_22325# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10051 vccd1 _0422_ _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10052 a_9021_29575# a_9117_29397# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X10053 _0481_ a_12263_20495# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10054 vssd1 _0246_ a_24485_17607# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10055 a_17565_13621# _0595_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10056 _0416_ a_2010_24759# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10057 vccd1 a_5499_5249# a_5323_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X10058 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10059 a_26505_21807# a_26339_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10060 a_13809_15829# a_13643_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10061 a_11142_23983# _0707_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10062 a_19496_24233# cal_lut\[83\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X10063 a_11555_14557# a_10773_14191# a_11471_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10064 _0392_ a_3288_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X10065 a_18111_25589# net47 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X10066 vssd1 io_in[1] a_1407_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X10067 a_26919_18909# a_26137_18543# a_26835_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10068 a_19915_19453# dbg_result[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X10070 a_11172_5487# a_10773_5487# a_11046_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10071 a_3117_12533# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X10073 a_10699_24233# _0681_ a_10784_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10075 cal_lut\[36\] a_14675_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10076 _0022_ a_15575_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X10077 a_23973_15279# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10078 a_15925_25437# a_15391_25071# a_15830_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10079 a_12705_22895# a_12539_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10081 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4068_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X10082 a_10331_20969# _0670_ a_10413_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10084 vccd1 a_13571_25339# a_13487_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10085 a_16238_7913# _0544_ a_16158_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10087 a_7381_20969# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X10088 vccd1 a_17895_17973# a_17811_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10089 _0296_ a_22240_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X10091 a_2023_19319# _0745_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X10092 vccd1 a_14507_3855# a_14675_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10093 a_13629_4943# _0118_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10094 a_9750_23983# _0720_ a_9372_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X10095 a_21591_2589# a_20727_2223# a_21334_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10096 a_3851_25045# _0802_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X10097 a_9681_2045# a_9411_1679# a_9591_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10098 a_27802_13924# a_27595_13865# a_27978_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X10099 a_9068_10703# cal_lut\[187\] a_8948_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X10100 a_11704_29423# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X10101 vccd1 _0878_ a_14747_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10102 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10103 vccd1 a_23547_26921# a_23554_26825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10104 vccd1 _0486_ a_19256_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X10105 vccd1 a_4584_24759# _0799_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X10106 vccd1 _0784_ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10107 a_28031_11471# a_27333_11477# a_27774_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10108 a_7564_31599# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X10110 a_21717_4399# a_20727_4399# a_21591_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10111 _0382_ clknet_1_0__leaf__0380_ a_6391_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10114 vccd1 _0290_ a_12355_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X10116 vssd1 net65 a_10875_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X10117 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd a_2879_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10118 a_1952_27247# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X10119 a_6182_22895# clknet_0_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X10120 a_10379_6740# _0304_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R25 temp1.capload\[10\].cap_50.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
R26 temp1.capload\[1\].cap_56.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10121 vssd1 net6 a_1837_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10122 vccd1 cal_lut\[134\] a_9542_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10123 vssd1 a_22403_22075# a_22361_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10124 vssd1 a_3155_16911# _0421_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10126 cal_lut\[51\] a_15687_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10127 a_4277_27221# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X10128 _0473_ a_22875_17249# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X10129 vssd1 net45 a_17323_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10130 vssd1 a_2014_14709# a_1972_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10132 a_22185_27791# _0054_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10133 a_14829_27497# cal_lut\[7\] a_14747_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10134 _0000_ a_1867_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10135 a_4153_9839# _0000_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10136 a_2137_20719# _0744_ a_1919_20693# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X10137 a_23818_19061# a_23650_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10139 vccd1 a_5583_6031# a_5751_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10142 _0214_ a_16076_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X10143 vssd1 a_21878_17143# _0692_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X10144 a_16585_16617# _0613_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X10145 a_12521_27247# a_12355_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10146 vccd1 _0807_ a_2564_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X10147 vssd1 a_19333_25223# _0221_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X10148 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10149 cal_lut\[122\] a_9615_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10150 vccd1 _0705_ a_10607_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10152 a_20112_12265# _0444_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10153 a_7917_27247# a_6927_27247# a_7791_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10156 a_22813_19631# a_22266_19905# a_22466_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10157 a_24941_23261# a_24407_22895# a_24846_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10158 a_4708_16143# _0411_ _0387_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X10159 vssd1 a_19763_4074# _0117_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10160 _0225_ a_14375_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10161 vssd1 cal_lut\[115\] a_22240_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10162 a_23650_19087# a_23377_19093# a_23565_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10163 vssd1 cal_lut\[4\] a_10832_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10164 vssd1 a_23763_4943# _0476_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10165 vccd1 a_2235_9303# _0838_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10166 a_19862_11039# a_19694_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10167 vccd1 _0353_ a_27259_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10168 cal_lut\[147\] a_10995_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10169 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10170 _0144_ a_6375_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X10171 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10172 cal_lut\[185\] a_15779_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10173 vssd1 net23 a_7847_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10174 a_27732_9839# a_27333_9839# a_27606_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10175 a_10083_24135# _0712_ a_10229_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10176 vssd1 _0584_ a_20141_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10177 a_4805_19087# _0427_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X10178 a_6541_14741# a_6375_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10179 a_19763_28010# _0223_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X10180 a_4705_27552# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10181 a_9647_14709# a_9823_15041# a_9775_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X10182 a_4277_27221# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X10183 a_3656_25847# temp1.dac_vout_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X10186 _0451_ a_22843_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X10188 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10189 vccd1 cal_lut\[7\] a_12443_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10190 a_6391_16911# _0447_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10192 cal_lut\[45\] a_15963_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10193 vccd1 a_23361_9985# _0659_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X10194 a_1932_22711# _0410_ a_1860_22711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X10195 vssd1 _0674_ a_11348_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X10196 a_5796_31849# a_5547_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10197 vccd1 a_2564_25045# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10198 a_27163_8573# cal_lut\[166\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X10199 _0436_ a_1683_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10200 vccd1 net75 _0395_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10201 vssd1 a_8543_30485# net11 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X10202 a_17673_26159# a_17507_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10204 vccd1 dbg_result[3] a_13942_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10205 vssd1 clknet_1_0__leaf__0380_ _0384_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10207 vssd1 net27 a_3799_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10209 _0356_ a_27163_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X10210 vssd1 _0216_ a_16355_29397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10211 vccd1 dbg_result[1] a_21721_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X10212 a_14185_27247# cal_lut\[8\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X10213 _0765_ _0752_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10214 vssd1 a_5644_12533# a_5404_12797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.07 as=0.172 ps=1.83 w=0.65 l=0.25
X10215 cal_lut\[61\] a_22863_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10216 vccd1 a_18151_21271# _0464_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10217 a_10488_31849# a_10239_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10218 _0108_ a_21371_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10219 _0267_ a_17135_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10220 a_13530_23439# a_13091_23445# a_13445_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10222 _0513_ a_9779_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X10223 a_22383_18793# _0647_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X10224 a_22779_1679# a_21997_1685# a_22695_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10225 a_12433_1679# _0183_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10226 cal_lut\[61\] a_22863_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10227 vssd1 a_8146_18796# a_8104_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X10228 a_12061_17455# a_11895_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10229 a_17870_28157# a_17555_28023# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10230 vccd1 net31 a_17323_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10231 a_9933_19061# _0589_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X10232 a_26123_14165# net37 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10233 a_5377_18319# net72 _0195_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10235 a_7952_13103# a_7553_13103# a_7826_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10236 a_17107_4073# net31 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10237 a_7102_21807# _0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10238 _0651_ a_10699_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10239 vccd1 a_6799_28853# a_6541_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X10241 vccd1 cal_lut\[66\] a_20775_14967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10242 vssd1 _0495_ a_15821_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10243 a_5825_17999# _0384_ a_5460_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10244 vccd1 a_11931_15645# a_12099_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10245 vccd1 temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10246 a_2044_29423# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X10247 a_9671_21495# _0627_ a_9905_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X10248 cal_lut\[179\] a_16147_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10249 vccd1 a_15998_25183# a_15925_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10251 a_13254_9295# a_12981_9301# a_13169_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10252 a_10832_30663# net8 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X10253 a_2959_25071# _0807_ a_2564_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X10254 a_21331_18543# _0442_ a_21217_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.137 ps=1.07 w=0.65 l=0.15
X10255 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10256 vccd1 net42 a_27167_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10257 vccd1 cal_lut\[67\] a_23299_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10258 a_20032_10499# _0260_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10259 vccd1 net78 a_8665_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X10260 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10261 a_7607_2589# a_6909_2223# a_7350_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10263 a_26505_21807# a_26339_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10265 vccd1 _0455_ a_16311_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10266 a_4066_7396# a_3859_7337# a_4242_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X10267 vssd1 _0452_ a_18765_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10268 vssd1 a_11214_5599# a_11172_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10269 vssd1 a_17930_24095# a_17888_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10270 vssd1 a_6607_9514# _0139_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10271 vssd1 _0748_ _0776_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10272 a_26111_20541# a_25891_20553# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10273 vccd1 a_8544_17429# _0433_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10274 a_26081_14557# a_25743_14343# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10275 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10276 vssd1 a_25198_17973# a_25156_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10277 a_13119_3855# a_12337_3861# a_13035_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10278 a_11019_2197# _0363_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X10279 a_21003_8320# cal_lut\[111\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10280 vssd1 clknet_1_1__leaf_io_in[0] a_5915_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10281 a_11965_8527# cal_lut\[99\] a_11527_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10282 vccd1 _0090_ a_18489_28169# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10283 a_26410_18909# a_25971_18543# a_26325_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10284 a_21081_9839# _0104_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10285 a_3991_26409# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X10286 cal_lut\[139\] a_5843_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10287 _0232_ a_23391_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X10288 a_9305_14191# _0079_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10289 a_9775_15101# cal_lut\[79\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X10290 a_3128_28879# a_2879_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10291 _0237_ a_12723_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10292 a_12610_14557# a_12337_14191# a_12525_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10293 a_22790_11471# cal_lut\[14\] a_22633_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10294 a_26233_16367# _0072_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10295 vccd1 a_17543_14735# a_17711_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10296 vccd1 a_16731_1653# _0333_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X10298 a_19756_16617# _0872_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10299 a_11693_10383# cal_lut\[39\] a_11609_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10300 vssd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X10301 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6467_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10302 a_15462_19997# a_15189_19631# a_15377_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10304 _0127_ a_8767_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10305 a_14151_11079# _0474_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X10306 a_9209_22895# _0712_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10307 a_1846_14735# a_1573_14741# a_1761_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10308 a_12985_10615# _0260_ a_13148_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10309 a_22714_13215# a_22546_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10310 vccd1 a_14967_1501# a_15135_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10311 a_22011_1135# cal_lut\[151\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X10312 _0196_ _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10313 vssd1 cal_lut\[2\] a_8393_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10314 vssd1 a_11366_28588# dbg_result[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X10315 a_16373_16341# _0621_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X10316 a_21975_2741# a_22151_3073# a_22103_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X10317 a_1761_12559# _0200_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10318 a_3974_13103# _0808_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X10320 vssd1 _0316_ a_7891_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10321 cal_lut\[121\] a_8419_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10322 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10323 a_24551_5461# a_24842_5761# a_24793_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X10324 vssd1 a_8419_6843# a_8377_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10325 vccd1 _0450_ a_22843_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X10326 a_24971_5487# a_24842_5761# a_24551_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10327 a_25125_23445# a_24959_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10329 a_14177_24533# a_14011_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10330 vssd1 a_3848_24135# _0823_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X10331 vccd1 a_13968_17218# a_13751_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.0672 ps=0.74 w=0.42 l=0.15
X10333 vccd1 a_20775_26311# cal_lut\[88\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10334 net48 a_6927_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X10336 a_20417_13249# _0528_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10337 a_7381_20969# _0766_ a_7583_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10338 _0379_ a_3575_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X10339 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10340 vccd1 _0234_ a_20359_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10341 vccd1 a_21759_10107# a_21675_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10342 a_14523_16885# dbg_result[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X10343 a_13135_15253# _0266_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X10344 a_4653_14013# _0808_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10345 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd _0817_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10346 a_6546_26159# _0399_ a_6460_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X10347 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10348 _0294_ a_18515_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10349 vccd1 a_27590_7093# a_27517_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10350 dbg_result[3] a_7410_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X10351 a_24938_15823# a_24499_15829# a_24853_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10352 vccd1 cal_lut\[171\] a_27163_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10353 a_14441_22895# cal_lut\[9\] a_14369_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10355 vccd1 a_17187_13255# _0601_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10356 vssd1 cal_lut\[122\] a_10325_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10357 vssd1 _0386_ _0197_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10359 a_23855_7119# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10360 a_4153_8751# _0140_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10361 a_2313_15823# _0198_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10362 a_22638_25437# a_22199_25071# a_22553_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10364 a_6459_32463# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X10365 _0764_ _0521_ a_8117_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10366 vccd1 a_25143_6031# _0341_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10367 vssd1 a_18326_7637# a_18255_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X10368 a_12613_10499# _0655_ a_12541_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10369 a_7895_11690# _0881_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10370 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_5796_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X10371 a_3421_24233# _0412_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X10372 _0873_ a_19756_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X10373 a_12778_14303# a_12610_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10374 vssd1 a_27774_9951# a_27732_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10375 a_22838_3133# a_22523_2999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10376 a_6814_7119# a_6541_7125# a_6729_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10378 vccd1 _0814_ a_7111_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X10379 vccd1 a_19303_17607# _0610_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10380 vssd1 cal_lut\[121\] a_8164_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10381 a_19011_19407# _0442_ a_18907_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X10382 vccd1 a_23707_8029# a_23875_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10384 a_15170_21237# a_15002_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10385 vssd1 a_8539_2986# _0180_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10386 a_17743_2741# cal_lut\[155\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X10387 a_7291_25615# _0724_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10388 a_13047_10927# a_12827_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10389 _0670_ _0669_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10390 vssd1 _0387_ a_3851_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.133 ps=1.06 w=0.65 l=0.15
X10391 a_10347_25071# _0720_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10392 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10393 cal_lut\[68\] a_24519_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10394 vssd1 a_15779_1653# a_15737_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10395 vssd1 _0733_ a_7553_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X10396 a_12352_5487# _0451_ a_12162_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X10397 vccd1 net44 a_16863_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10398 a_6467_15823# _0839_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10399 a_23063_3855# a_22199_3861# a_22806_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10401 cal_lut\[113\] a_18171_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10402 vssd1 _0416_ a_1683_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10404 a_4801_20175# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X10406 a_9815_1501# a_9117_1135# a_9558_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10407 _0450_ a_17651_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10408 vssd1 _0456_ a_17312_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X10409 a_21307_19997# a_20525_19631# a_21223_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10410 vssd1 a_7239_17999# a_7410_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X10411 a_21717_10927# a_20727_10927# a_21591_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10412 a_8393_17277# a_8123_16911# a_8303_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10413 vccd1 a_9275_15444# _0079_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10414 a_24972_23983# a_24573_23983# a_24846_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10415 vccd1 a_15963_17723# a_15879_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10416 vccd1 cal_lut\[171\] a_23792_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10419 _0243_ a_23299_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10420 a_9678_5737# _0498_ a_9678_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X10422 _0536_ a_20359_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10423 a_14699_6549# _0290_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X10424 a_4242_7119# a_3995_7497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10425 vssd1 net27 a_3799_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10426 vssd1 clknet_1_0__leaf__0380_ _0381_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10427 vccd1 a_6674_16620# dbg_result[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10428 a_17543_14735# a_16679_14741# a_17286_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10429 a_26677_14191# a_26123_14165# a_26330_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10430 vccd1 cal_lut\[9\] a_13363_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10431 a_26983_9295# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10432 vssd1 a_2931_22325# _0783_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10433 vccd1 a_21721_18909# _0465_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X10434 a_12691_10901# net29 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10435 a_24306_12836# a_24106_12681# a_24455_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10436 a_10488_30761# a_10239_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10437 a_6705_23759# _0720_ _0827_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10439 a_5759_3855# a_4977_3861# a_5675_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10440 a_9403_32143# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X10441 a_2222_20969# _0746_ a_1919_20693# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X10442 a_4885_6037# a_4719_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10443 a_7079_24233# _0437_ a_6987_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X10444 a_18975_1679# a_18795_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10445 a_8951_6825# cal_lut\[127\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X10447 vssd1 a_8527_3855# a_8695_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10448 vssd1 _0462_ a_22175_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X10449 _0429_ a_3615_17999# a_4143_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10450 vccd1 a_21975_2741# _0337_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X10451 a_12978_23261# a_12705_22895# a_12893_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10453 a_10761_9839# cal_lut\[189\] a_10689_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10455 a_9117_1135# a_8951_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10456 a_13926_17277# a_13551_16911# a_13835_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.064 ps=0.725 w=0.42 l=0.15
X10457 vssd1 a_20414_22325# a_20372_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10458 vccd1 _0420_ a_4077_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10459 a_18873_16911# _0028_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10460 vccd1 net42 a_27167_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10461 net28 a_6007_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10463 vccd1 _0864_ a_11987_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10464 a_4259_13103# _0397_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X10466 vccd1 a_26210_9951# a_26137_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10467 cal_lut\[151\] a_20931_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10468 vccd1 a_15531_24135# _0645_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10471 a_3850_23759# _0790_ a_4040_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10472 vssd1 a_13052_15797# _0519_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X10473 vccd1 clknet_1_1__leaf_io_in[0] a_4443_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10474 a_7277_18543# a_7111_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10475 a_16574_17455# _0612_ a_16820_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X10476 a_14265_29257# a_13275_28885# a_14139_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10477 a_9831_24501# _0718_ a_10049_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X10478 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10479 vccd1 a_6674_16620# dbg_result[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X10480 a_20763_1679# a_19899_1685# a_20506_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10482 vssd1 clknet_1_0__leaf_io_in[0] a_1407_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10484 vccd1 a_28031_15823# a_28199_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10485 a_17105_10357# _0623_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X10486 _0092_ a_13275_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10488 vssd1 _0694_ a_10746_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10489 a_2366_25615# _0801_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X10490 a_10497_7119# a_9963_7125# a_10402_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10491 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10492 vccd1 a_5883_27221# a_5890_27521# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10494 a_22270_1679# a_21831_1685# a_22185_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10495 net36 a_24499_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X10496 a_12955_25834# _0848_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10497 vccd1 _0237_ a_16771_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X10498 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10499 a_21265_7815# cal_lut\[111\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X10501 vccd1 _0154_ a_20237_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10502 vccd1 net29 a_9687_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10503 net46 a_18111_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10504 vssd1 a_16373_16341# _0625_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X10505 net31 a_16640_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10506 vssd1 cal_lut\[5\] a_12856_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10507 a_7289_25321# _0724_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10508 vssd1 net40 a_12539_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10509 vssd1 _0425_ _0472_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10510 a_9551_2388# _0368_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X10511 a_3128_27791# a_2879_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10512 a_10505_17705# net12 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X10513 _0346_ a_25783_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10515 vssd1 cal_lut\[90\] a_17961_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10516 vssd1 _0478_ a_22988_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X10518 a_13771_21263# a_12907_21269# a_13514_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10519 vccd1 a_11207_14954# _0004_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10520 vssd1 a_20506_1653# a_20464_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10521 a_4169_21583# _0780_ a_3759_21495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X10522 vccd1 a_2511_21263# io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10523 a_4143_17999# a_3615_17999# _0429_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10524 vssd1 _0057_ a_24377_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10525 cal_lut\[125\] a_15135_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10526 a_15427_21263# a_14729_21269# a_15170_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10527 a_24435_14735# a_23653_14741# a_24351_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10528 vssd1 a_7775_6005# a_7733_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10529 vccd1 _0459_ a_19623_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10530 vssd1 a_6982_14709# a_6920_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X10531 a_9126_11177# cal_lut\[38\] a_9043_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10532 _0748_ _0721_ a_8951_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.26 ps=2.52 w=1 l=0.15
X10533 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10534 vccd1 _0033_ a_26309_20553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10535 vccd1 _0425_ a_5639_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10536 vccd1 a_16991_27613# a_17159_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10537 vssd1 _0685_ a_22291_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10538 a_9558_1247# a_9390_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10539 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10540 a_13441_21263# a_12907_21269# a_13346_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10541 a_10356_8751# cal_lut\[140\] a_10236_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X10543 a_14237_19881# a_14167_19783# _0448_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
X10547 a_18985_23805# cal_lut\[47\] a_18913_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10548 vccd1 a_9673_23047# _0726_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X10549 a_12161_7663# _0441_ a_12079_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10550 _0741_ a_2742_18082# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
R27 vccd1 temp1.capload\[11\].cap_51.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10552 vssd1 ctr\[2\] a_2153_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X10553 a_16679_26703# _0484_ a_16857_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10555 a_20322_7775# a_20154_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10556 vssd1 a_23139_13371# a_23097_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10557 a_26486_16479# a_26318_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10558 a_26283_8207# a_25585_8213# a_26026_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10559 a_27333_9839# a_27167_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10560 a_5278_12533# a_5404_12797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.217 pd=2.17 as=0.273 ps=1.61 w=0.82 l=0.25
X10561 vssd1 _0744_ a_2234_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X10562 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10563 a_22638_3855# a_22199_3861# a_22553_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10564 a_9941_14191# a_8951_14191# a_9815_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10565 a_23903_18695# _0460_ a_24137_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10566 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10567 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10569 vccd1 a_24835_5461# a_24842_5761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10570 a_25138_10927# a_24823_11079# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10571 _0071_ a_27351_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10572 a_21997_11471# cal_lut\[103\] a_21913_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10575 vssd1 a_14103_17455# _0447_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X10576 temp1.dac_vout_notouch_ net13 a_10232_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X10577 a_23063_25437# a_22199_25071# a_22806_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10578 _0420_ a_2288_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10579 vccd1 a_27035_8181# _0351_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X10580 vccd1 _0226_ a_17415_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10581 _0840_ a_6647_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X10582 a_12223_2741# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X10583 vccd1 cal_lut\[121\] a_8246_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X10584 _0557_ _0556_ a_12455_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.36 ps=2.72 w=1 l=0.15
X10585 vccd1 cal_lut\[118\] a_20775_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10586 a_7005_4551# cal_lut\[133\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X10587 vccd1 net25 a_15115_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10588 a_19819_2223# a_19690_2497# a_19399_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X10589 cal_lut\[126\] a_15503_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10590 vccd1 net10 a_10239_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X10591 vccd1 a_4678_26311# _0800_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X10592 a_8397_20983# dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10593 a_28031_17821# a_27167_17455# a_27774_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10594 vccd1 clknet_1_1__leaf_io_in[0] a_10331_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10595 a_20874_27765# a_20706_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10596 a_20572_6031# _0444_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10598 vssd1 clknet_0_temp1.i_precharge_n a_3882_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10599 _0182_ a_10055_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10600 _0838_ a_2235_9303# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10601 vccd1 a_20119_5853# a_20287_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10603 a_23690_10089# _0657_ a_23610_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10604 cal_lut\[22\] a_13295_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10605 a_23377_19093# a_23211_19093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10606 a_9568_31055# a_9319_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10607 net13 a_11120_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10608 a_3869_11989# clknet_0_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10609 vccd1 _0492_ a_16404_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X10610 vccd1 _0482_ a_16845_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X10611 a_20939_16911# a_20157_16917# a_20855_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10613 a_2329_18793# _0421_ a_2234_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0683 ps=0.745 w=0.42 l=0.15
X10614 vccd1 a_15170_10357# a_15097_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10615 vssd1 cal_lut\[89\] a_18560_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10616 vccd1 a_25014_8863# a_24941_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10617 vssd1 _0414_ _0773_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10618 vssd1 clknet_1_0__leaf_io_in[0] a_6375_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10619 a_15745_25071# _0045_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10620 a_6982_12127# a_6814_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10621 _0723_ a_8397_20983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X10622 vccd1 a_9452_32375# a_9403_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X10623 vssd1 dbg_result[1] a_14655_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10624 a_15909_7809# _0515_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X10625 _0451_ a_22843_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10626 a_11895_16617# _0609_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10627 vccd1 a_3859_7337# a_3866_7241# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10628 a_1951_28879# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X10629 vccd1 _0216_ a_14195_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X10631 vssd1 a_13203_14459# a_13161_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10632 vccd1 clknet_0_temp1.i_precharge_n a_1753_26133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10634 a_16297_10927# _0101_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10635 a_11981_11837# a_11711_11471# a_11891_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10636 a_10504_10703# cal_lut\[98\] a_9929_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X10638 _0609_ a_16373_13077# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.91 w=0.65 l=0.15
X10639 a_26778_22173# a_26505_21807# a_26693_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10640 vssd1 temp_delay_last a_4351_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X10641 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10642 a_4238_9117# a_3965_8751# a_4153_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10643 a_4075_14191# ctr\[1\] a_3981_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X10644 a_17835_7637# a_18119_7637# a_18054_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10645 a_6354_9117# a_6081_8751# a_6269_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10646 vccd1 a_7716_25589# _0750_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X10647 a_6729_17999# _0195_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X10648 vccd1 _0460_ a_10851_11079# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X10649 vssd1 _0619_ a_18669_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X10650 _0688_ a_21889_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.112 ps=0.995 w=0.65 l=0.15
X10651 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_2419_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X10652 a_25389_5487# a_24835_5461# a_25042_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10653 a_16853_8751# _0445_ a_16771_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10654 a_12691_10901# net29 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10656 vccd1 a_13422_9269# a_13349_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10657 a_25589_17455# _0069_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10658 a_10551_11471# a_9853_11477# a_10294_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10659 a_12455_18793# net16 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X10660 a_20963_15797# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X10661 vssd1 a_11458_27500# dbg_result[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X10662 vccd1 _0232_ a_23579_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10663 a_19333_24135# _0260_ a_19496_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10666 a_17651_28023# a_17935_28009# a_17870_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X10667 vssd1 a_23707_8029# a_23875_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10669 vssd1 a_21759_4667# a_21717_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10670 vssd1 a_20471_26677# a_20429_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10672 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10674 vssd1 a_5013_24825# a_4947_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10676 a_2010_24759# _0410_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10677 a_24915_21959# a_25011_21781# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10678 vssd1 a_2991_15797# a_2949_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10680 _0057_ a_23579_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X10681 a_10055_17455# _0662_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X10682 temp1.capload\[4\].cap.Y clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10683 _0167_ a_27259_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10684 vccd1 a_19199_13647# a_19367_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10685 vccd1 a_7410_14709# a_7323_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X10686 cal_lut\[113\] a_18171_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10687 a_2000_29111# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X10688 a_22396_2057# a_21997_1685# a_22270_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10690 vccd1 a_22291_20175# net43 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10691 vssd1 a_16550_11039# a_16508_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10692 a_3877_11703# _0808_ a_4040_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10693 a_4701_27791# a_4167_27797# a_4606_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10694 a_2701_21583# _0744_ a_2511_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.127 ps=1.04 w=0.65 l=0.15
X10695 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10696 a_3885_16189# _0411_ a_3796_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0619 ps=0.715 w=0.42 l=0.15
X10697 a_7741_8751# _0120_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10698 vssd1 a_19199_13647# a_19367_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10699 _0815_ a_7847_28992# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X10700 vssd1 net46 a_17783_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10701 a_17041_23805# a_16771_23439# a_16951_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10702 vssd1 a_12927_17723# a_12885_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10703 a_5418_9269# a_5250_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10705 _0850_ a_10699_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X10706 a_5250_3855# a_4811_3861# a_5165_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10707 vccd1 _0483_ a_15299_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10709 vssd1 _0265_ a_21279_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10710 net21 a_4995_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X10711 a_8348_32375# net10 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X10714 vssd1 a_20747_9269# a_20705_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10716 a_14195_10205# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10720 vssd1 _0290_ a_10835_4161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10721 a_18003_6941# a_17305_6575# a_17746_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10722 a_8108_22351# _0785_ a_7853_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X10723 _0234_ a_19940_19881# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X10724 net44 a_17875_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X10725 vssd1 net35 a_20819_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10726 a_20937_5487# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10728 vccd1 a_13514_21237# a_13441_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10729 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10730 vssd1 _0452_ a_16005_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10731 vssd1 a_9671_21495# _0677_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X10732 _0087_ a_21279_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10733 a_1679_22057# _0417_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10735 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10736 vccd1 _0464_ a_18611_20288# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10737 a_14250_15797# a_14082_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10738 a_7975_14557# a_7111_14191# a_7718_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10739 a_18918_22351# _0620_ a_18669_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10741 a_23299_24349# a_23119_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10742 a_24122_17188# a_23922_17033# a_24271_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X10743 vccd1 _0668_ a_11191_19659# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10744 vccd1 _0266_ a_14195_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X10745 a_8201_4943# _0145_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10746 a_18482_12533# a_18314_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10747 vccd1 a_8999_7828# _0121_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10748 cal_lut\[109\] a_22863_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10749 vccd1 net41 a_15023_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10750 a_4929_15307# ctr\[6\] a_4843_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X10751 a_24573_8751# a_24407_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10752 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10753 a_15561_18231# cal_lut\[95\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X10754 vccd1 a_23763_4943# _0476_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10755 vccd1 _0043_ a_17845_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10757 a_18731_12043# _0440_ a_18645_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X10758 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10759 vccd1 net42 a_25879_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10760 a_18642_27497# _0260_ a_18560_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10761 a_20758_9001# _0283_ a_20676_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10762 a_12161_12559# _0515_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10763 a_1735_27765# _0824_ a_1962_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X10764 a_5900_24527# _0795_ a_5645_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X10765 vssd1 a_5141_21781# _0756_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10766 _0385_ a_9835_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.178 ps=1.41 w=1 l=0.15
X10767 a_7645_14557# a_7111_14191# a_7550_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10768 a_11868_29967# a_11619_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X10769 _0386_ a_9559_26481# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10770 a_22764_4233# a_22365_3861# a_22638_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10771 a_4771_4917# a_4947_5249# a_4899_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X10772 a_17673_26159# a_17507_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10774 a_20981_17289# a_19991_16917# a_20855_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10775 _0455_ _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X10778 a_19465_16367# net18 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10780 a_21997_1685# a_21831_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10781 a_7826_9117# a_7387_8751# a_7741_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10782 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X10783 vssd1 _0420_ _0427_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10785 vssd1 a_16757_7637# _0498_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X10786 a_9125_10089# _0700_ a_9043_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X10788 a_9835_26703# ctr\[6\] a_9763_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0578 ps=0.695 w=0.42 l=0.15
X10789 vssd1 a_25271_23261# a_25439_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10790 vccd1 cal_lut\[104\] a_21034_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X10791 a_10715_21263# _0557_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10792 vssd1 a_17743_2741# _0339_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X10793 vccd1 a_6982_7093# a_6909_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10794 vssd1 a_6445_29111# net79 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X10795 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10796 a_1679_22057# _0414_ a_1461_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10798 vssd1 net41 a_14655_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10799 a_11014_22057# _0521_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X10800 a_16771_8320# cal_lut\[143\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10801 vccd1 _0442_ a_19303_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X10802 a_26339_7119# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10803 a_12061_17455# a_11895_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10804 vccd1 a_5179_14191# _0811_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10805 a_4947_24893# dbg_result[5] a_4584_24759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X10807 a_15565_8751# _0514_ a_15483_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10809 a_16079_3285# _0363_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X10810 a_3357_10383# a_2947_10615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X10811 a_25375_20407# a_25471_20407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10813 a_22685_5309# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X10814 vssd1 a_3155_9839# _0836_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X10815 a_25287_12533# a_25463_12865# a_25415_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X10816 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10817 vccd1 a_23231_3829# a_23147_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10819 _0291_ a_19619_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X10820 vssd1 a_8723_17130# _0002_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10821 a_4977_9301# a_4811_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10822 vssd1 _0377_ a_6099_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10823 vccd1 _0726_ a_9831_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X10824 a_17930_24095# a_17762_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X10827 vssd1 a_24243_19061# a_24201_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10828 _0425_ a_7631_17171# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10830 vssd1 net42 a_27167_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10831 a_21081_9839# _0104_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10832 vccd1 net40 a_13275_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10834 vssd1 _0390_ a_4487_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10836 a_11555_5853# a_10773_5487# a_11471_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10837 vccd1 a_20303_28879# a_20471_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10838 vssd1 a_12679_28010# _0007_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10839 a_19199_13647# a_18335_13653# a_18942_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10840 _0299_ a_7439_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10841 a_7826_6941# a_7553_6575# a_7741_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10842 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_1959_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X10843 a_12938_16617# _0836_ a_12856_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10844 a_9573_8585# a_8583_8213# a_9447_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10845 _0504_ a_8951_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X10846 a_4413_7497# a_3866_7241# a_4066_7396# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X10847 a_24099_4073# net33 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10849 _0190_ a_6099_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10850 a_13104_22895# a_12705_22895# a_12978_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10851 vccd1 a_14616_14709# _0872_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10852 a_6737_22671# _0432_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X10853 a_13512_13621# cal_lut\[10\] a_13732_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10854 a_9854_28879# a_9607_29257# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10855 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10856 vssd1 net1 a_10699_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X10857 a_9907_6031# a_9043_6037# a_9650_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10858 vssd1 cal_lut\[1\] a_9595_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10859 a_23943_6031# a_23763_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10860 a_27886_15645# a_27639_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X10861 a_13882_28853# a_13714_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10862 io_out[3] a_2287_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10863 a_15901_21835# _0483_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X10864 a_9671_21495# _0630_ a_9821_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X10865 vssd1 a_12263_20495# _0481_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10866 a_24485_17607# cal_lut\[74\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X10867 vccd1 a_10843_2197# _0373_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X10868 vssd1 a_14611_11079# _0563_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X10870 a_12150_26703# a_11711_26709# a_12065_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10872 vccd1 a_13838_19319# a_13714_19407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X10873 a_17042_4221# a_16727_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X10874 a_20947_21263# a_20083_21269# a_20690_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10876 a_24761_7119# _0163_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10877 a_15887_19997# a_15189_19631# a_15630_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10878 a_8289_14741# a_8123_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10879 a_2384_13353# _0411_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X10880 a_14507_3855# a_13809_3861# a_14250_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10881 a_9482_6031# a_9043_6037# a_9397_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10883 net23 a_5324_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X10884 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd _0419_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10885 vccd1 _0447_ a_13751_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X10886 a_26467_10205# a_25769_9839# a_26210_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10887 net9 a_9687_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X10888 vccd1 a_4774_27765# a_4701_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10889 vccd1 a_20931_1653# a_20847_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10890 a_2447_19087# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X10891 vccd1 _0486_ a_14829_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10892 vssd1 a_20119_5853# a_20287_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10893 a_9034_6825# cal_lut\[145\] a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10894 vssd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X10895 a_18739_12559# a_18041_12565# a_18482_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10896 a_26309_20553# a_25755_20393# a_25962_20452# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X10897 vccd1 a_22165_10357# _0635_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X10898 _0445_ a_17927_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10899 a_20390_6031# _0585_ a_20141_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10900 vccd1 _0410_ a_6463_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X10901 a_18314_12559# a_17875_12565# a_18229_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10903 temp1.dac_vout_notouch_ net14 a_11704_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X10904 vssd1 _0055_ a_23273_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X10905 vccd1 ctr\[3\] a_4816_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10906 vccd1 a_24473_9813# _0511_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X10907 a_22855_27247# a_22719_27221# a_22435_27221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10909 vccd1 a_11857_18517# _0628_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X10912 vccd1 a_16069_22923# _0487_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X10913 a_25415_12925# cal_lut\[175\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X10914 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7564_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X10915 vssd1 a_8390_23439# clknet_1_1__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10916 a_5486_9001# _0838_ a_5404_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X10917 vssd1 net9 a_9687_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10920 vccd1 _0105_ a_19225_9673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X10921 a_5376_4233# a_4977_3861# a_5250_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10923 vssd1 a_13698_23413# a_13656_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10924 a_6381_25321# _0750_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10926 a_23631_11079# _0511_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X10927 a_25842_17567# a_25674_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10928 a_15002_21263# a_14563_21269# a_14917_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10930 a_4676_25223# ctr\[7\] a_4818_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X10932 vssd1 a_5418_9269# a_5376_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X10933 _0653_ a_10607_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X10934 vssd1 a_7959_27515# dec1.i_ones vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10935 vssd1 _0725_ a_9308_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10936 cal_lut\[167\] a_27923_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10937 _0701_ a_9043_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X10938 a_23211_22351# _0863_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10939 a_7718_14303# a_7550_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X10940 a_17682_16100# a_17475_16041# a_17858_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X10941 a_12343_16617# _0519_ _0626_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10942 vssd1 _0371_ a_14379_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X10943 vccd1 a_7718_14303# a_7645_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10944 vccd1 a_24455_5639# cal_lut\[160\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10947 a_4679_19319# net21 a_5007_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10948 a_25965_14013# a_25695_13647# a_25875_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X10949 a_8251_13469# a_7387_13103# a_7994_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10951 a_4931_24135# ctr\[5\] a_5077_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X10952 a_15724_18115# cal_lut\[95\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X10953 a_15193_15431# _0491_ a_15356_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10954 vssd1 net33 a_22199_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10955 vccd1 _0508_ a_23395_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10956 a_1458_30199# a_1554_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X10957 vccd1 cal_lut\[161\] a_18475_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X10958 a_18671_9513# net35 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10959 a_20303_28879# a_19439_28885# a_20046_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X10960 _0719_ _0718_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10961 a_5545_23439# _0737_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10962 vccd1 _0481_ a_9411_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10963 vccd1 a_15519_29789# a_15687_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10965 a_27755_9117# a_27057_8751# a_27498_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10966 a_17627_9295# a_16845_9301# a_17543_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10967 a_17611_16201# a_17475_16041# a_17191_16055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X10968 a_20253_1679# _0150_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10969 ctr\[4\] a_4647_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10970 _0678_ a_10331_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X10971 vccd1 a_19167_19061# a_18698_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X10972 a_17949_28885# a_17783_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10973 a_10965_25321# _0732_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X10974 a_21936_21807# a_21537_21807# a_21810_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10975 a_3882_16911# net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10976 vccd1 a_11527_9303# net29 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10977 a_15548_19407# a_15494_19319# a_15452_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.107 ps=0.98 w=0.65 l=0.15
X10978 a_7952_8751# a_7553_8751# a_7826_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10979 a_17857_25437# a_17323_25071# a_17762_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X10980 ctr\[4\] a_4647_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10981 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X10982 a_11292_30663# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X10983 a_20522_21263# a_20249_21269# a_20437_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X10984 vccd1 _0467_ a_17507_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X10985 a_18229_12559# _0017_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10986 cal_lut\[83\] a_18355_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10987 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10988 vssd1 _0740_ a_5089_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X10989 vssd1 cal_lut\[117\] a_19433_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10990 a_12127_21959# _0671_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X10991 a_10046_8751# cal_lut\[122\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X10992 cal_lut\[45\] a_15963_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10993 cal_lut\[80\] a_9983_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10994 a_4977_3861# a_4811_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10996 a_9827_29245# a_9607_29257# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X10997 vssd1 a_14307_28853# a_14265_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10998 vccd1 cal_lut\[56\] a_22747_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11000 a_9384_29967# a_9135_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X11001 _0806_ _0804_ a_3421_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X11002 a_23201_22895# _0468_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X11003 a_10596_17705# _0663_ a_10423_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X11004 a_15354_1653# a_15186_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11005 a_24771_6031# a_24591_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11006 vccd1 a_18107_7338# _0112_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11007 cal_lut\[39\] a_10719_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11008 vccd1 a_1673_16911# a_1773_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X11009 vccd1 a_25042_13077# a_24971_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X11010 a_9858_25615# _0719_ a_9555_25847# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X11011 a_22105_18115# _0458_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X11012 a_10229_24233# _0705_ a_10083_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X11013 vccd1 a_25991_23413# a_25907_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11014 a_12202_14851# _0246_ a_12120_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11015 a_10773_14191# a_10607_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11016 vccd1 clknet_1_0__leaf_io_in[0] a_6375_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11018 vssd1 _0850_ a_25143_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X11019 vccd1 _0316_ a_6375_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X11020 vssd1 a_16991_22173# a_17159_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11021 cal_lut\[39\] a_10719_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11022 vssd1 net44 a_20083_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11023 vccd1 cal_lut\[152\] a_22471_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11024 vssd1 a_1651_14165# _0411_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X11025 a_9117_1135# a_8951_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11026 vccd1 a_10943_23671# _0717_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X11027 a_8025_21263# _0437_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X11028 a_9815_1501# a_8951_1135# a_9558_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11029 vssd1 a_17651_8181# _0450_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X11031 vccd1 a_15469_26935# _0270_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X11033 a_9678_29156# a_9471_29097# a_9854_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11035 vccd1 net46 a_17507_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11036 a_13751_16911# a_13551_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X11037 a_24853_15823# _0068_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11038 vssd1 cal_lut\[23\] a_18192_15529# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11039 net30 a_3339_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X11040 a_27710_15253# a_27503_15253# a_27886_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11041 vccd1 a_22431_13866# _0013_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11042 vssd1 a_24731_6740# _0163_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11043 a_11207_14954# _0844_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11044 _0464_ a_18151_21271# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X11045 vccd1 cal_lut\[65\] a_19100_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X11046 a_7102_21807# _0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X11047 a_9595_5737# cal_lut\[128\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X11048 cal_lut\[84\] a_20287_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11049 vccd1 a_4406_8863# a_4333_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11050 a_21384_14191# a_20985_14191# a_21258_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11051 vccd1 a_6522_8863# a_6449_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11053 _0193_ _0839_ a_5181_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11055 a_19683_2197# net31 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11056 net19 a_21095_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11057 a_23021_16617# _0475_ a_23223_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11058 a_7147_3677# a_6449_3311# a_6890_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11059 a_19244_22671# cal_lut\[65\] a_18669_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X11060 vssd1 _0453_ a_17783_21271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11061 a_2823_15823# a_2125_15829# a_2566_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11062 vssd1 a_5883_27221# a_5890_27521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11063 cal_lut\[84\] a_20287_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11064 vssd1 _0629_ a_9933_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11065 a_19625_18543# dbg_result[1] a_19525_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X11066 vssd1 _0751_ _0752_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X11067 a_15378_22895# _0645_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X11068 vssd1 _0167_ a_28057_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X11069 a_27639_15279# a_27503_15253# a_27219_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X11070 a_14471_6031# _0290_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11071 vccd1 a_15541_9985# _0550_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X11072 a_24094_14709# a_23926_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11073 a_15722_3829# a_15554_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11074 vssd1 a_21391_19899# a_21349_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11075 _0716_ _0628_ a_9503_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11076 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X11077 a_9608_6409# a_9209_6037# a_9482_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11078 vssd1 _0651_ a_11343_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11079 a_13751_16911# a_13968_17218# a_13926_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11080 a_3056_31375# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X11082 a_7980_7235# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11083 a_3891_13353# ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X11084 a_15105_8751# _0505_ a_15023_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11086 vccd1 cal_lut\[46\] a_16986_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11087 _0277_ a_11891_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11088 _0165_ a_25143_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11089 _0524_ a_19071_11584# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X11090 _0711_ a_10915_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X11091 a_25962_20452# a_25755_20393# a_26138_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X11092 cal_lut\[67\] a_22955_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11093 vssd1 net11 a_9319_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11094 a_4307_24310# _0822_ a_3848_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X11095 a_14153_20884# _0485_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11096 vssd1 a_17543_14735# a_17711_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11097 a_4563_12559# a_3781_12565# a_4479_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11098 a_18637_5487# _0443_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11099 vssd1 a_13295_13371# a_13253_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11100 a_8951_25321# _0714_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11101 a_19220_26819# cal_lut\[52\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X11102 a_22790_11471# _0451_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11103 a_11120_28853# net14 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X11104 a_24971_13103# a_24842_13377# a_24551_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11105 _0372_ a_16859_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11106 net78 a_8671_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11107 vssd1 _0481_ a_19409_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11108 vssd1 _0679_ a_10688_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X11109 a_4437_15055# _0811_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11110 vssd1 a_5031_27791# a_5199_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11111 vssd1 a_1551_19605# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11112 vccd1 cal_lut\[15\] a_22596_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X11113 a_18119_7637# net32 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11115 a_11609_10383# _0653_ a_11527_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11116 vssd1 _0307_ a_14195_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11118 a_6458_20175# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11120 a_13625_23439# a_13091_23445# a_13530_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11121 a_21872_25731# _0260_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11122 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11124 dbg_result[5] a_11366_28588# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X11125 vssd1 _0617_ a_16373_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11127 _0617_ a_16390_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X11129 vssd1 _0175_ a_26309_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X11130 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11131 a_19303_17607# _0454_ a_19537_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11132 a_20598_16885# a_20430_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11133 a_26777_6575# a_25787_6575# a_26651_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11134 vccd1 a_23351_8439# _0640_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X11135 vccd1 a_12955_25834# _0008_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11138 vccd1 _0217_ a_17047_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11139 a_9487_26481# clknet_1_1__leaf__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X11140 vccd1 a_7102_21807# clknet_0__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11142 vssd1 _0631_ a_11715_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11143 a_15722_3829# a_15554_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11144 a_6647_15823# a_6467_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11145 vssd1 clknet_1_1__leaf_io_in[0] a_10331_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11146 vssd1 a_15439_17130# _0095_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11147 vccd1 a_20046_28853# a_19973_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11148 a_6646_21041# _0435_ a_6645_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X11150 vccd1 _0453_ a_18519_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11151 vssd1 cal_lut\[14\] a_23297_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11153 vssd1 _0519_ a_11439_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X11154 a_15193_14343# _0851_ a_15356_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11155 temp1.dac_vout_notouch_ net14 a_9384_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X11156 vccd1 a_2023_19319# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11157 a_7182_2589# a_6743_2223# a_7097_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11158 a_22457_6037# a_22291_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11159 a_20203_24527# a_19421_24533# a_20119_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11160 vccd1 _0326_ a_6559_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11161 a_15645_29423# a_14655_29423# a_15519_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11162 vssd1 a_8143_14459# a_8101_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11163 _0405_ net71 a_7111_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11164 a_25003_24833# _0237_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X11165 a_10911_3677# a_10129_3311# a_10827_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11166 a_25218_5853# a_24971_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X11167 a_3965_8751# a_3799_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11168 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_2668_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X11169 temp1.dac.vdac_single.en_pupd _0801_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11170 _0195_ _0384_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11171 vssd1 _0859_ a_17599_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11172 _0724_ a_9372_24135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11173 a_20683_21972# _0241_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11174 vssd1 a_20690_18517# _0452_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11175 cal_lut\[68\] a_24519_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11176 a_8117_19407# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11177 vssd1 a_14523_16885# _0442_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X11178 a_25927_10602# _0355_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11179 a_16097_12015# cal_lut\[191\] a_16025_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11180 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_4351_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11181 a_1857_21365# clknet_1_1__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11182 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11183 vssd1 a_12898_10901# a_12827_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X11185 vssd1 _0336_ a_22659_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11186 a_21675_11293# a_20893_10927# a_21591_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11187 a_10779_28701# a_10497_28335# a_10685_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X11188 vssd1 a_7410_14709# dbg_result[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X11189 a_8017_3855# _0132_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11191 vssd1 _0420_ a_2722_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11192 a_10809_19605# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X11193 vssd1 net48 a_13551_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11194 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11195 vccd1 _0838_ a_12723_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11196 a_18475_18695# _0454_ a_18709_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11197 a_5181_16617# _0839_ _0193_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11198 a_17231_14191# cal_lut\[23\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11199 vssd1 _0762_ a_2614_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X11200 _0183_ a_11987_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11201 a_13672_5737# _0566_ a_13570_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11202 a_3965_9839# a_3799_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11203 _0506_ a_20943_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X11204 a_4333_9117# a_3799_8751# a_4238_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11205 a_1846_14735# a_1407_14741# a_1761_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R28 net62 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11206 _0017_ a_17599_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11207 vccd1 a_3695_23671# _0791_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X11208 a_23079_17607# cal_lut\[26\] a_23205_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X11209 a_25957_9839# _0169_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11211 _0056_ a_23395_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11212 a_2773_9991# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X11213 vssd1 a_20775_27412# _0053_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11214 vccd1 a_24351_14735# a_24519_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11215 vccd1 _0310_ a_10331_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11216 temp1.dac_vout_notouch_ net13 a_10416_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X11218 a_11789_3311# _0129_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11219 a_2772_23983# a_2741_24135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X11220 vccd1 a_7994_6687# a_7921_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11221 a_18272_12265# _0502_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X11222 _0716_ _0626_ a_9586_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X11223 vccd1 a_25502_21781# a_25431_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X11224 a_6427_11445# cal_lut\[190\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X11225 a_14855_12265# _0491_ _0515_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11227 a_4435_30761# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X11229 _0559_ a_18243_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11230 a_6541_7125# a_6375_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11231 vssd1 a_9559_26481# _0386_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11232 vccd1 cal_lut\[60\] a_21218_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11234 vssd1 a_25931_8725# _0350_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X11235 a_7553_13103# a_7387_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11236 a_6619_23439# _0435_ a_6527_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X11237 vccd1 net20 a_20267_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X11238 vssd1 a_18114_26271# a_18072_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11239 a_8803_15823# a_8105_15829# a_8546_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11240 a_10872_28701# a_10331_28335# a_10779_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X11241 _0732_ _0720_ a_10417_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11242 dbg_result[1] a_6674_16620# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X11243 _0498_ a_16757_7637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X11244 a_25355_24349# a_24573_23983# a_25271_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11245 _0151_ a_21463_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11246 a_4425_5487# a_4259_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11247 a_7281_27247# _0212_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11248 vccd1 _0477_ a_17231_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X11249 vccd1 net23 a_7939_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11250 vccd1 a_18355_24251# a_18271_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11252 vssd1 _0704_ _0705_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11253 a_21009_18365# cal_lut\[60\] a_20937_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11254 cal_lut\[186\] a_18355_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11257 a_4027_16144# temp_delay_last vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11258 vccd1 a_15611_1679# a_15779_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11259 a_3695_23671# _0744_ a_4040_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X11261 a_5675_13469# a_4811_13103# a_5418_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11262 a_23297_12925# a_23027_12559# a_23207_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11263 a_14155_29397# a_14331_29397# a_14283_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X11264 a_4143_17999# _0421_ a_3785_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11265 cal_lut\[120\] a_15411_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11267 a_21310_15529# _0222_ a_21228_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11268 vssd1 _0497_ a_9779_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X11269 a_1753_26133# clknet_0_temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11270 a_2887_25615# ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X11271 a_16481_27247# _0042_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11272 vssd1 _0877_ a_25235_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11273 vccd1 cal_lut\[116\] a_23117_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X11274 a_15220_29423# a_14821_29423# a_15094_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11275 a_6729_30199# ctr\[10\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X11276 _0022_ a_15575_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11277 vssd1 cal_lut\[12\] a_20308_14441# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11278 vssd1 net19 a_14441_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11279 a_5345_13469# a_4811_13103# a_5250_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11281 a_22494_10383# _0633_ a_22414_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X11282 cal_lut\[85\] a_21759_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11283 a_10969_20495# _0667_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11284 vssd1 _0838_ a_2419_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X11285 _0592_ dbg_result[5] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11286 vssd1 a_15193_15431# _0518_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X11287 vssd1 a_17895_2491# a_17853_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11288 vccd1 a_25287_12533# _0361_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X11291 vccd1 a_13698_23413# a_13625_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11292 a_10402_1679# a_10129_1685# a_10317_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11294 a_13997_15823# _0035_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11295 _0038_ a_9411_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11296 a_11189_25321# _0731_ _0749_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.305 ps=1.61 w=1 l=0.15
X11298 a_24761_25071# _0086_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11299 vssd1 net42 a_25879_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11300 vccd1 _0443_ a_22291_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X11301 vssd1 _0878_ a_14747_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11304 a_14703_21972# _0213_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11305 _0737_ _0420_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.176 ps=1.39 w=1 l=0.15
X11306 a_12856_16617# _0836_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11307 a_4678_26311# ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11308 vccd1 a_23719_12791# cal_lut\[15\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11309 a_10562_19319# _0589_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X11310 a_22625_17973# _0642_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X11311 a_5271_3677# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11312 a_21353_6575# a_21187_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11313 vccd1 _0720_ a_9678_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X11315 a_9390_14557# a_8951_14191# a_9305_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11316 vssd1 _0330_ a_22151_3073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11317 a_1937_6549# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11318 clknet_1_1__leaf_io_in[0] a_6182_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11319 _0429_ a_3615_17999# a_4143_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11320 _0216_ a_13459_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11321 _0194_ _0383_ a_6651_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11323 a_6914_28111# _0826_ a_6828_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X11324 cal_lut\[182\] a_9983_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11325 a_7829_3861# a_7663_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11327 vssd1 _0141_ a_4413_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X11328 a_21081_4399# _0114_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11329 a_19496_10089# cal_lut\[105\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X11330 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11331 vssd1 a_7716_22325# _0786_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X11332 vssd1 a_22988_4917# _0479_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X11333 a_5165_9295# _0138_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11334 a_14917_10383# _0100_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11335 a_18371_26525# a_17507_26159# a_18114_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11336 a_20390_27497# _0222_ a_20308_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11337 vssd1 a_12263_20495# _0481_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X11338 a_26677_14191# a_26130_14465# a_26330_14165# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11339 a_22523_2999# a_22619_2999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11340 a_5170_10660# a_4970_10505# a_5319_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11341 a_19862_15391# a_19694_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11342 a_14283_29423# cal_lut\[49\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X11343 a_14905_18115# dbg_result[2] a_14833_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11344 a_7308_2223# a_6909_2223# a_7182_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11345 a_18177_5487# _0462_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11346 a_12311_11079# a_12407_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11347 _0805_ a_3525_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X11348 vccd1 net34 a_26983_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11349 a_15461_7497# a_14471_7125# a_15335_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11352 a_14576_24905# a_14177_24533# a_14450_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11353 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11355 vccd1 net36 a_27167_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11356 vssd1 a_18355_25339# a_18313_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11357 a_7921_6941# a_7387_6575# a_7826_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11358 a_20733_8573# cal_lut\[166\] a_20661_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11359 a_19537_16367# cal_lut\[29\] a_19465_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11360 vssd1 a_27590_7093# a_27548_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11361 a_22388_12879# _0456_ a_21897_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X11362 vssd1 net41 a_7939_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11363 net29 a_11527_9303# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11364 a_18475_19783# _0453_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11365 a_22672_13103# a_22273_13103# a_22546_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11366 a_18041_26525# a_17507_26159# a_17946_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11368 a_15128_10761# a_14729_10389# a_15002_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11369 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11370 vssd1 a_8251_6941# a_8419_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11371 _0144_ a_6375_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11372 a_13245_10927# a_12698_11201# a_12898_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11373 a_12351_12381# a_12171_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11374 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_6835_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11375 vssd1 a_13403_25437# a_13571_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11376 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11377 vccd1 a_4484_30663# a_4435_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X11378 _0800_ a_4678_26311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11379 vccd1 a_8297_20765# a_8397_20983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X11380 a_16757_7637# _0441_ a_17003_7691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X11381 vssd1 _0659_ a_12310_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X11382 vccd1 a_12985_10615# _0276_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X11383 cal_lut\[102\] a_16975_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11384 vccd1 a_12127_21959# _0709_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X11385 _0787_ _0432_ a_5547_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11387 a_9447_8207# a_8583_8213# a_9190_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11388 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X11389 vssd1 a_13459_22359# _0841_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X11390 vssd1 _0874_ a_21279_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11391 cal_lut\[167\] a_27923_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11392 a_24573_25071# a_24407_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11393 vccd1 a_9983_1403# a_9899_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11394 vssd1 _0481_ a_10356_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X11397 cal_lut\[130\] a_12467_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11398 vccd1 a_3707_9303# net27 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11400 vccd1 a_10844_31029# net8 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X11402 vccd1 net35 a_16679_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11403 a_3877_11703# ctr\[4\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X11404 vccd1 cal_lut\[191\] a_12351_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11405 a_24573_23983# a_24407_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11406 vssd1 net27 a_4811_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11408 dbg_result[4] a_11458_27500# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X11410 _0773_ _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=2.1 w=0.65 l=0.15
X11411 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11412 vccd1 _0482_ a_15557_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X11413 _0030_ a_21279_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11414 a_10108_4373# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X11415 a_26242_13103# a_25927_13255# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X11416 vssd1 net43 a_25971_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11418 vccd1 a_14287_17999# net18 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11419 _0222_ a_20963_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11420 vccd1 _0631_ a_11799_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X11421 a_20249_3311# a_20083_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11422 a_4583_10615# a_4679_10615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11423 _0739_ _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11424 _0052_ a_19531_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11425 a_21166_25437# a_20893_25071# a_21081_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11426 vccd1 a_7347_24501# _0751_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X11427 a_24034_4221# a_23719_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X11428 a_11609_8207# _0493_ a_11693_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11429 vccd1 a_8971_15797# a_8887_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11430 a_15397_9661# cal_lut\[106\] a_15325_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11432 a_12736_14191# a_12337_14191# a_12610_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11433 vssd1 a_3479_7351# cal_lut\[142\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11434 vssd1 a_19763_28010# _0048_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11435 _0136_ a_3983_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11436 _0325_ a_4163_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11438 _0410_ ctr\[8\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X11439 a_15870_10089# _0548_ a_15790_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X11440 vssd1 a_23631_11079# _0512_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X11441 a_25355_23261# a_24573_22895# a_25271_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11442 cal_lut\[144\] a_7407_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11443 a_17935_28009# net46 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11444 vccd1 a_5418_13215# a_5345_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11445 vccd1 net58 temp1.capload\[3\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11446 vssd1 net31 a_20083_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11447 a_7559_18909# a_7111_18543# a_7465_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X11449 a_22796_11791# _0452_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X11450 vccd1 a_14031_12533# a_13947_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11451 a_9678_5737# cal_lut\[146\] a_9595_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11452 vssd1 a_11214_14303# a_11172_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11453 vssd1 _0168_ a_26677_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X11454 dbg_result[4] a_11458_27500# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X11455 vccd1 _0451_ a_9043_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X11456 a_2221_13255# ctr\[1\] a_2384_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11457 vccd1 cal_lut\[130\] a_12535_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11458 _0564_ a_14287_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11459 a_5227_26935# ctr\[7\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11460 a_4491_25654# _0828_ a_4032_25847# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X11461 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11462 _0281_ a_18055_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11463 a_25410_10901# a_25210_11201# a_25559_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11464 a_10871_27613# a_10589_27247# a_10777_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X11466 cal_lut\[90\] a_20287_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11467 a_2271_12559# a_1573_12565# a_2014_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11468 vccd1 a_19255_19631# _0462_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11469 vssd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11470 vccd1 ctr\[2\] a_5460_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11471 vccd1 _0297_ a_23671_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11473 a_6645_8573# a_6375_8207# a_6555_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11474 a_21081_10927# _0103_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11475 vccd1 _0412_ a_2010_24759# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X11476 a_10413_20719# _0677_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11477 a_15785_15279# _0467_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11479 _0773_ ctr\[5\] a_5837_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11480 _0862_ a_9131_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11481 vssd1 a_5583_6031# a_5751_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11483 a_18029_16201# a_17475_16041# a_17682_16100# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X11484 a_20775_26311# a_20871_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11485 a_9436_10927# cal_lut\[188\] a_9316_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X11486 a_15207_18543# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.109 ps=1.36 w=0.42 l=0.15
X11487 a_27491_17130# _0250_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11488 a_7393_21263# _0669_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11489 a_15722_12533# a_15554_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11490 a_17611_16201# a_17482_15945# a_17191_16055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11491 a_20325_12533# _0535_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11492 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4811_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11493 vccd1 _0229_ a_21463_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11494 _0401_ ctr\[7\] a_5722_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X11495 net43 a_22291_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X11496 a_8573_17999# _0439_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11497 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11498 vssd1 a_15193_14343# _0852_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X11500 vssd1 net26 a_13275_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11501 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5547_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11503 vssd1 a_12778_3829# a_12736_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11505 a_22247_9991# _0450_ a_22481_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11506 vssd1 net30 a_12999_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11507 _0679_ a_10975_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11508 vssd1 net47 a_22199_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11509 a_22821_8585# a_21831_8213# a_22695_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11510 vccd1 a_9613_20693# a_9643_21046# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11512 a_16734_27359# a_16566_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11514 cal_lut\[185\] a_15779_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11516 vssd1 ctr\[9\] _0410_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11517 vccd1 ctr\[9\] a_5911_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
R29 net61 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11518 a_5989_11293# a_5455_10927# a_5894_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11519 a_18313_23983# a_17323_23983# a_18187_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11521 a_19881_7663# a_19715_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11522 vccd1 cal_lut\[117\] a_23351_8439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X11523 vccd1 _0421_ _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11525 vccd1 a_11458_27500# a_11371_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X11527 vccd1 net48 a_12723_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11528 vssd1 a_10995_3579# a_10953_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11529 a_15611_1679# a_14747_1685# a_15354_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11530 cal_lut\[120\] a_15411_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11531 _0431_ a_1773_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X11533 a_11191_19659# _0666_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X11534 cal_lut\[191\] a_7407_12283# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11535 vccd1 a_3072_19637# _0747_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X11536 a_4977_13103# a_4811_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11537 a_18027_19783# _0467_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X11538 a_15561_18231# _0260_ a_15724_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11539 a_20997_24893# a_20727_24527# a_20907_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11540 vccd1 cal_lut\[25\] a_23759_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11541 _0021_ a_11987_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11542 _0560_ a_18611_20288# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11543 _0341_ a_25143_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X11544 a_4310_8439# a_4406_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X11545 vssd1 a_18671_9513# a_18678_9417# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11546 vccd1 a_18114_26271# a_18041_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11547 a_17135_25615# a_16955_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11548 vssd1 a_7350_2335# a_7308_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11549 a_5667_6031# a_4885_6037# a_5583_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11551 a_19402_25589# a_19234_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11552 cal_lut\[74\] a_28199_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11553 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11554 a_21441_11791# cal_lut\[158\] a_21003_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11555 a_22185_23439# _0060_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11556 a_25389_5487# a_24842_5761# a_25042_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X11558 _0864_ a_11707_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11560 a_17651_8181# _0445_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X11561 vccd1 a_1407_15823# net7 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11562 _0746_ _0414_ a_2887_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.36 ps=2.72 w=1 l=0.15
X11563 vssd1 net46 a_17507_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11564 _0033_ a_25235_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11565 vssd1 a_24455_5639# cal_lut\[160\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11566 vssd1 _0837_ a_1867_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11567 _0427_ _0420_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11568 vccd1 _0728_ a_7853_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11569 a_15877_5309# _0452_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X11570 vssd1 _0234_ a_20359_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11571 a_4265_20175# _0447_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11572 vssd1 a_15354_1653# a_15312_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11573 _0522_ a_19807_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11576 _0460_ a_20451_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X11577 a_18145_10749# a_17875_10383# a_18055_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11578 vssd1 net46 a_19439_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11579 vssd1 a_9595_26703# a_10043_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0683 ps=0.745 w=0.42 l=0.15
X11582 vssd1 a_4583_10615# cal_lut\[189\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11584 vccd1 _0290_ a_19163_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X11585 a_7741_8751# _0120_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11587 a_9607_29257# a_9478_29001# a_9187_29111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X11588 vccd1 a_13751_16911# _0477_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X11589 _0811_ a_5179_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X11590 vssd1 a_20303_28879# a_20471_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11591 _0425_ a_7631_17171# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11592 cal_lut\[95\] a_15687_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11593 a_2287_22325# clknet_1_1__leaf_io_in[0] a_2569_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X11594 a_22194_19631# a_21879_19783# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X11595 vccd1 cal_lut\[81\] a_12202_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11596 vssd1 a_25375_20407# cal_lut\[34\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11597 a_12134_7093# a_11966_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11598 vccd1 _0705_ a_7101_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X11599 vccd1 a_15170_21237# a_15097_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11600 vccd1 net21 _0771_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11601 cal_lut\[23\] a_17711_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11602 vssd1 a_15871_2741# a_15829_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11603 cal_lut\[95\] a_15687_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11604 cal_lut\[54\] a_21299_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11605 vccd1 a_4676_25223# _0828_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11606 a_14167_19783# _0442_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X11608 a_17578_6941# a_17139_6575# a_17493_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11609 vssd1 a_9555_25847# _0721_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X11610 a_9547_3073# _0363_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X11611 a_10773_5487# a_10607_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11612 a_7323_7119# a_6541_7125# a_7239_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11613 vccd1 a_16550_11039# a_16477_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11614 a_25397_8751# a_24407_8751# a_25271_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11615 a_16761_24527# cal_lut\[46\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X11616 a_19383_16911# a_18685_16917# a_19126_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11617 a_13422_9269# a_13254_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11618 a_26444_16367# a_26045_16367# a_26318_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11619 vssd1 a_5170_10660# a_5099_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X11620 vccd1 _0425_ a_12263_20495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X11621 vssd1 _0610_ a_16574_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X11622 a_27123_15431# a_27219_15253# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11623 vccd1 a_6982_17973# a_6916_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X11624 a_17814_14441# _0851_ a_17732_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11625 _0305_ a_11247_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11626 _0872_ a_14616_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X11627 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11628 vccd1 a_25842_17567# a_25769_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11629 a_5675_9295# a_4811_9301# a_5418_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11630 net38 a_16731_9813# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11632 vccd1 a_1464_23957# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X11633 vssd1 a_17283_28853# _0217_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X11634 _0847_ a_12443_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11637 a_19303_18695# a_19667_18517# a_19625_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11638 a_13445_23439# _0009_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11639 a_21971_13879# _0505_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11640 a_19057_26935# cal_lut\[52\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X11642 vccd1 a_9471_29097# a_9478_29001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11643 vssd1 _0404_ a_6732_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X11644 a_12391_7119# a_11693_7125# a_12134_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11645 vccd1 a_14103_17455# _0447_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11646 _0478_ a_22843_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X11647 a_13882_28853# a_13714_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11648 a_13073_21269# a_12907_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11650 a_20203_5853# a_19421_5487# a_20119_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11651 vccd1 _0461_ a_19255_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X11652 _0669_ _0662_ a_10137_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X11653 _0358_ a_27071_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11654 a_23757_11177# _0506_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X11655 a_9595_16367# _0692_ a_9749_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11657 a_21721_18909# dbg_result[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X11658 _0098_ a_12263_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11659 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5087_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X11660 a_6537_19605# clknet_0__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11661 vccd1 a_13139_7351# _0570_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X11662 vccd1 _0414_ a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11663 vccd1 a_4277_23957# a_4307_24310# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11665 vccd1 _0812_ a_4988_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X11666 vssd1 a_2722_20175# _0424_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11667 a_27149_18005# a_26983_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11668 _0871_ a_18100_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X11669 a_8335_16733# a_7553_16367# a_8251_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11670 vssd1 a_26819_6843# a_26777_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11671 vssd1 net1 a_2235_9303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11672 a_12351_12559# _0650_ a_12245_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.19 ps=1.38 w=1 l=0.15
X11673 _0861_ a_7751_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11674 vccd1 a_10570_1653# a_10497_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11675 _0883_ a_11891_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X11676 cal_lut\[40\] a_13939_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11677 vccd1 io_in[3] a_1407_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11678 a_12709_27247# _0007_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11679 a_19057_26935# _0222_ a_19220_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11680 a_2317_16911# net5 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11681 vssd1 a_23351_7338# _0109_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11682 a_28031_10205# a_27167_9839# a_27774_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11683 _0191_ a_12815_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11684 a_18693_20541# _0464_ a_18611_20288# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11685 a_22875_17249# _0460_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X11686 vssd1 a_22523_5175# _0687_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11687 vssd1 a_7994_13215# a_7952_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11688 _0466_ a_17999_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X11689 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11690 vssd1 _0838_ a_4167_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X11692 a_10497_3677# a_9963_3311# a_10402_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11694 cal_lut\[40\] a_13939_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11695 vccd1 cal_lut\[47\] a_18751_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X11696 vccd1 a_9385_4373# _0503_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X11697 a_9551_2388# _0368_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11698 a_9853_11477# a_9687_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11699 vccd1 _0376_ a_5639_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11700 _0301_ a_14651_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11701 vccd1 dec1.i_ones a_9223_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X11702 a_14686_13353# _0851_ a_14604_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11704 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11705 a_24268_10703# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X11706 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4811_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11707 a_5461_27069# ctr\[8\] a_5389_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11708 _0686_ a_22291_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X11709 a_1458_30199# a_1554_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X11710 a_15603_23439# a_14821_23445# a_15519_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11711 a_4624_15823# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11713 a_7853_25615# _0748_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11714 a_4520_20175# _0760_ a_4265_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X11715 vssd1 a_21591_4765# a_21759_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11716 a_8485_23145# _0728_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X11717 _0626_ _0519_ a_12343_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11718 vssd1 a_1407_4399# net1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11719 a_25585_8213# a_25419_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11720 _0189_ a_5639_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11721 vssd1 a_13571_23163# a_13529_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11722 vccd1 _0483_ a_16035_18112# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X11723 a_24823_15444# _0244_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11724 vssd1 _0385_ _0196_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11725 vccd1 a_5307_29789# a_5475_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11726 vccd1 a_15163_9527# _0562_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X11727 a_6072_31055# a_5823_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X11729 a_9559_26481# _0592_ a_9487_26481# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.0672 ps=0.85 w=0.64 l=0.15
X11732 a_15005_2773# a_14839_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11733 vccd1 a_13415_20884# _0039_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11734 vccd1 _0316_ a_3983_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X11735 vccd1 cal_lut\[41\] a_16158_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11736 a_3072_19637# _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11737 _0508_ a_19308_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X11738 vccd1 a_7439_4373# _0299_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X11739 vccd1 net46 a_19439_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11740 a_8975_18793# _0439_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11741 a_12265_24233# _0708_ _0712_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11742 vssd1 a_20683_21972# _0065_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11744 vccd1 a_4479_12559# a_4647_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11745 a_23391_21263# a_23211_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11746 a_17191_16055# a_17482_15945# a_17433_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X11747 a_14082_3855# a_13643_3861# a_13997_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11748 vccd1 cal_lut\[107\] a_17871_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11749 vssd1 net7 a_1932_17271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
R30 vssd1 net65 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11751 a_18291_9527# a_18387_9527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11752 vssd1 a_17159_27515# a_17117_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11753 a_26042_10205# a_25603_9839# a_25957_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11754 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X11755 vssd1 a_8251_16733# a_8419_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11756 a_3851_15253# _0839_ a_4407_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X11757 vssd1 net33 a_22291_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11758 vssd1 a_4479_12559# a_4647_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11760 a_4215_7485# a_3995_7497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X11762 vssd1 net26 a_9595_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X11763 vssd1 a_18187_24349# a_18355_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11764 _0856_ a_23207_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11765 a_9956_31375# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X11766 vssd1 _0226_ a_17415_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11767 a_16681_16617# _0617_ a_16585_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11768 vccd1 _0854_ a_20635_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11769 a_27245_8751# _0166_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11770 a_12429_17821# a_11895_17455# a_12334_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11772 a_10953_7497# a_9963_7125# a_10827_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11773 vccd1 cal_lut\[57\] a_23391_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11775 vccd1 net24 a_6375_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11777 vssd1 _0483_ a_16097_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11778 vssd1 a_20325_12533# _0538_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X11779 a_26609_7485# a_26339_7119# a_26519_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11780 vssd1 a_4679_19319# _0742_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X11781 a_14337_8779# _0472_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X11782 a_2247_27791# _0817_ a_1735_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X11783 vssd1 a_1651_14165# _0411_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11784 cal_lut\[156\] a_18723_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11785 vccd1 a_9615_8181# a_9531_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11786 vssd1 _0882_ a_9411_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11787 vssd1 a_10083_24135# _0713_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X11788 a_10746_10615# _0696_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X11789 a_4744_22057# _0747_ a_4283_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
X11790 a_1639_15444# _0388_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11791 vccd1 a_28199_15797# a_28115_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11792 a_17095_5639# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11793 vssd1 net30 a_10607_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11795 a_16035_15279# cal_lut\[35\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11797 vssd1 _0401_ a_4897_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X11798 a_27337_7119# _0162_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11799 vssd1 a_20287_11195# a_20245_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11800 a_6799_28853# ctr\[9\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11801 vccd1 _0425_ a_4805_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X11802 vssd1 _0406_ a_8951_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11803 vssd1 _0543_ _0555_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11804 a_17704_6575# a_17305_6575# a_17578_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11805 vccd1 a_7073_25589# _0792_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11807 vccd1 a_21591_10205# a_21759_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11808 _0766_ a_8478_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X11809 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_3128_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X11810 a_25064_16201# a_24665_15829# a_24938_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11811 a_16925_8573# cal_lut\[143\] a_16853_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11812 a_18555_3677# a_17857_3311# a_18298_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11813 a_18383_5175# _0462_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X11814 net27 a_3707_9303# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11815 _0870_ a_24863_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11817 a_4816_16617# _0382_ a_5181_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11818 a_4789_9839# a_3799_9839# a_4663_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11819 a_15285_17455# _0095_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11820 a_21591_25437# a_20893_25071# a_21334_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11821 vccd1 a_4313_17429# _0790_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11822 _0154_ a_19439_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11823 a_20090_19453# a_19715_19087# a_19999_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.064 ps=0.725 w=0.42 l=0.15
X11825 a_27590_7093# a_27422_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11826 vssd1 a_13422_9269# a_13380_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11827 a_7733_10761# a_6743_10389# a_7607_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11828 _0855_ a_21735_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11829 vccd1 a_22843_9295# _0451_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11830 a_19605_28885# a_19439_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11831 vccd1 a_20119_24527# a_20287_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11832 vssd1 _0712_ a_9750_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
X11833 a_7631_17171# dbg_result[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X11834 a_27330_9117# a_26891_8751# a_27245_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11835 ctr\[8\] a_5199_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11836 a_3990_19631# _0421_ a_4180_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11837 vssd1 _0643_ a_22383_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11838 vccd1 a_5583_14735# a_5751_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11840 vccd1 a_18907_12533# a_18823_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11842 a_23683_27081# a_23547_26921# a_23263_26935# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X11843 vssd1 a_20119_24527# a_20287_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11844 a_6982_14709# a_6823_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X11845 a_23804_8323# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11846 vccd1 _0392_ a_3799_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11848 a_8229_25071# _0713_ a_8419_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11851 a_7704_8323# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11852 vssd1 a_25455_17999# a_25623_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11853 a_1761_14735# _0199_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11854 a_27731_14025# a_27595_13865# a_27311_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X11855 a_28157_11849# a_27167_11477# a_28031_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11856 _0882_ a_8947_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X11857 a_20832_28169# a_20433_27797# a_20706_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11858 a_3995_18793# _0426_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11859 vccd1 _0476_ a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X11861 vssd1 a_1963_21365# _0772_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11862 vccd1 cal_lut\[66\] a_21310_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11863 vccd1 _0450_ a_10699_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11864 vssd1 a_7618_26935# _0409_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X11865 a_10685_28335# _0197_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X11866 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11867 _0213_ a_14604_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X11868 vssd1 _0461_ a_19255_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11869 a_25783_14735# a_25603_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11870 a_21353_6575# a_21187_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11871 _0201_ a_3799_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11872 a_16955_19087# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X11873 vssd1 a_2750_14303# a_2708_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11874 a_7741_10927# _0037_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11875 a_13714_4943# a_13441_4949# a_13629_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11878 vssd1 a_25014_24095# a_24972_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X11879 vccd1 a_1743_18259# _0422_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11880 a_11765_17973# net4 a_12269_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X11882 a_4479_12559# a_3615_12565# a_4222_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11883 a_17762_24349# a_17489_23983# a_17677_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11884 vccd1 a_17095_16055# cal_lut\[78\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11885 a_13525_20175# _0425_ a_13722_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11888 a_10881_10499# _0515_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X11889 _0212_ a_6914_28111# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11890 vccd1 net21 a_4154_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X11891 a_7839_32463# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X11892 vssd1 _0227_ a_19531_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11893 vccd1 _0675_ a_10603_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X11894 a_18659_10615# _0514_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11895 vssd1 net35 a_17875_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11896 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8024_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X11897 vccd1 _0748_ a_7939_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X11898 a_20815_6941# a_20635_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11899 a_12846_7913# _0572_ a_12597_7809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X11903 _0237_ a_12723_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X11904 vccd1 cal_lut\[116\] a_23426_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11905 cal_lut\[128\] a_10075_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11906 vccd1 _0741_ a_4995_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11907 a_21954_20291# _0222_ a_21872_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11909 a_8286_4943# a_8013_4949# a_8201_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11910 a_14331_29397# _0216_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X11911 vssd1 a_3339_9295# net30 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11912 vssd1 _0398_ a_4437_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X11913 vccd1 _0380_ a_7102_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11914 io_out[1] a_1551_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11915 vccd1 _0329_ a_9963_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X11916 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6072_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X11917 a_4149_12559# a_3615_12565# a_4054_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X11918 _0654_ a_11527_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X11920 net74 a_6003_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X11921 a_12035_26324# _0846_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11922 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11923 a_22431_7338# _0343_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11924 _0532_ a_19807_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X11925 a_4180_19631# a_3799_19631# _0737_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11926 vccd1 a_10699_4399# _0850_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11928 vssd1 a_18815_28853# a_18773_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11929 vccd1 _0789_ a_4129_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X11930 vccd1 a_17599_6039# _0514_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11931 vssd1 a_9091_29111# ctr\[12\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11932 a_6087_16733# a_5639_16367# a_5993_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X11935 vssd1 _0755_ _0827_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X11936 a_17168_13647# _0597_ a_17066_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11937 vccd1 cal_lut\[184\] a_13672_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X11938 a_20039_18695# _0485_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X11939 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9956_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X11941 vssd1 a_21851_14459# a_21809_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11942 vssd1 a_8999_7828# _0121_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X11943 a_11142_24233# _0681_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X11944 a_15335_7119# a_14471_7125# a_15078_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11945 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11946 a_17907_10955# _0445_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X11947 a_4988_27497# _0401_ _0207_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X11948 a_21537_21807# a_21371_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11949 a_15606_11177# _0260_ a_15524_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11951 vssd1 a_24683_14191# _0352_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11952 vccd1 clknet_1_1__leaf_net67 net70 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11953 vssd1 a_4167_16367# _0839_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X11954 a_19333_9991# _0283_ a_19496_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11955 a_5433_29423# a_4443_29423# a_5307_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11956 vccd1 a_18482_12533# a_18409_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X11957 a_10781_8573# _0450_ a_10699_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X11958 a_18763_20871# _0453_ a_18937_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X11959 a_14208_4233# a_13809_3861# a_14082_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11960 vssd1 a_19303_2375# cal_lut\[155\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11961 vccd1 io_in[4] a_1407_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11962 vccd1 cal_lut\[53\] a_20390_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11963 a_21717_9839# a_20727_9839# a_21591_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11964 a_11868_30761# a_11619_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X11965 vccd1 clknet_0_io_in[0] a_6182_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11966 vssd1 a_15903_3285# _0366_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X11967 a_26168_9839# a_25769_9839# a_26042_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11968 a_9179_28309# _0839_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.178 ps=1.4 w=0.42 l=0.15
X11969 cal_lut\[166\] a_26451_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11970 io_out[0] a_2023_19319# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11971 a_9037_11837# a_8767_11471# a_8947_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X11973 a_20119_24527# a_19255_24533# a_19862_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11974 a_17168_12559# _0456_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X11975 a_8543_30485# temp1.dac.parallel_cells\[4\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X11976 vssd1 _0414_ a_1867_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11977 a_5115_27791# a_4333_27797# a_5031_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11978 a_23351_21959# _0443_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X11979 a_5583_14735# a_4719_14741# a_5326_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X11980 a_12153_2223# a_11987_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11981 a_16127_5056# cal_lut\[179\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11982 cal_lut\[136\] a_7131_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11983 a_23167_26935# a_23263_26935# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11984 a_7676_14191# a_7277_14191# a_7550_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11985 vccd1 a_17291_29397# a_17298_29697# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11986 a_4917_26165# _0410_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.13 ps=1.11 w=0.42 l=0.15
X11987 a_7097_2223# _0186_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X11989 a_17095_10004# _0286_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X11990 vccd1 _0631_ _0665_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11991 a_24945_17999# _0074_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X11992 vssd1 a_15812_9269# net35 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X11993 vccd1 cal_lut\[53\] a_20039_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X11994 a_27215_13879# a_27311_13879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11995 _0603_ a_16035_6144# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X11997 a_1863_24233# _0791_ a_1464_23957# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11998 vssd1 a_13714_19407# _0495_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X11999 vccd1 a_7410_17973# dbg_result[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12000 _0029_ a_19991_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12001 a_12893_22895# _0081_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12002 a_3885_21583# _0427_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X12003 a_24030_20452# a_23830_20297# a_24179_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12005 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12006 _0574_ a_13091_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X12007 a_23155_6031# a_22457_6037# a_22898_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12008 a_3325_8903# _0838_ a_3488_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12009 vccd1 a_15887_19997# a_16055_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12010 a_5253_14735# a_4719_14741# a_5158_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12011 vssd1 a_17746_6687# a_17704_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12012 vssd1 _0602_ a_16737_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X12013 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X12014 a_15101_1679# _0184_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12015 a_17421_13103# cal_lut\[173\] a_17349_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12016 vccd1 a_2439_12533# ctr\[1\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12017 a_19878_26703# a_19439_26709# a_19793_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12018 vssd1 _0729_ a_10347_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X12019 a_20249_21269# a_20083_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12020 a_25603_14735# _0352_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12021 vssd1 a_5418_13215# a_5376_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12022 a_6909_2223# a_6743_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12023 _0456_ a_18597_13077# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X12024 vccd1 a_19333_13255# _0860_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X12025 vccd1 a_16219_25623# net47 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12026 vssd1 a_23355_23671# _0471_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X12027 vssd1 a_2439_12533# ctr\[1\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12028 _0785_ _0434_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12029 a_10051_3855# a_9871_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12030 a_19583_2741# cal_lut\[154\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X12032 a_14967_1501# a_14269_1135# a_14710_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12033 a_5894_11293# a_5455_10927# a_5809_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12035 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd a_3128_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X12036 a_13809_3861# a_13643_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12038 a_14265_5321# a_13275_4949# a_14139_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12039 vccd1 a_5843_9269# a_5759_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12040 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4068_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X12042 a_6090_27221# a_5890_27521# a_6239_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12043 a_10160_16201# a_9761_15829# a_10034_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12044 a_8059_14557# a_7277_14191# a_7975_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12045 a_4789_8751# a_3799_8751# a_4663_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12046 vssd1 net28 a_7387_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12047 vccd1 _0834_ a_4811_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X12048 cal_lut\[66\] a_21115_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12049 _0521_ a_8645_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12050 a_6905_8751# a_5915_8751# a_6779_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12051 vccd1 a_13512_13621# _0576_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X12052 a_15715_5175# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12053 a_27456_8751# a_27057_8751# a_27330_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12054 a_10417_25935# _0715_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12055 vssd1 net31 a_20727_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12056 a_25743_14343# a_25839_14165# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X12058 vssd1 net23 a_6743_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12059 a_7239_14735# a_6541_14741# a_6982_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X12061 _0514_ a_17599_6039# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X12062 vssd1 _0839_ _0197_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12063 net69 clknet_1_1__leaf_net67 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12065 vccd1 a_9678_29156# a_9607_29257# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X12066 a_15879_28879# a_15097_28885# a_15795_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12067 a_9423_18793# _0520_ _0680_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12070 a_15623_26324# _0219_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12071 a_27774_15797# a_27606_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12072 vccd1 a_26330_14165# a_26259_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X12073 a_20621_27791# _0053_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12074 a_23079_17607# _0479_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X12076 vccd1 cal_lut\[173\] a_27531_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12077 _0423_ _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12078 vssd1 a_15561_18231# _0274_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X12079 a_26045_16367# a_25879_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12080 a_23450_7775# a_23282_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12082 vssd1 _0814_ a_8001_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12084 vccd1 a_15370_19407# _0467_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12086 a_20112_12265# _0522_ a_20010_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X12087 vccd1 _0418_ a_2887_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12088 vccd1 _0486_ a_14185_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X12089 a_22779_23439# a_21997_23445# a_22695_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12090 a_23443_20407# a_23539_20407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X12091 a_19303_18695# dbg_result[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X12092 vccd1 cal_lut\[148\] a_13139_7351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X12093 vccd1 a_4461_25913# a_4491_25654# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12094 a_23481_23759# _0463_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X12095 a_17302_2589# a_16863_2223# a_17217_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12096 a_15354_1653# a_15186_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12097 cal_lut\[109\] a_22863_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12098 a_21334_25183# a_21166_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12099 a_9949_15823# _0003_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12100 vccd1 a_3175_14459# a_3091_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12101 vssd1 a_16911_29575# cal_lut\[44\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12102 a_20308_14441# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12103 vccd1 a_15531_4564# _0178_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12104 a_15979_3855# a_15281_3861# a_15722_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12105 _0287_ a_17871_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12106 a_5377_16143# clknet_1_0__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12107 vccd1 net9 a_9595_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X12108 a_15857_15279# cal_lut\[36\] a_15785_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12109 a_22695_8207# a_21831_8213# a_22438_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12110 vssd1 net36 a_27167_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12111 vssd1 _0492_ a_10504_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X12112 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_6644_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X12113 a_13905_26703# _0092_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12114 a_16225_8751# cal_lut\[120\] a_16153_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12116 a_7365_12015# a_6375_12015# a_7239_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12118 a_16679_3677# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12119 vssd1 cal_lut\[160\] a_24861_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12120 vssd1 _0492_ a_11965_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X12121 a_10635_13469# a_9853_13103# a_10551_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12122 a_22431_13866# _0855_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12123 a_10108_4373# _0850_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X12124 vccd1 _0418_ a_2366_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X12125 _0235_ a_21136_23145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X12126 _0376_ a_5083_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12127 a_8645_17999# _0433_ a_8573_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X12128 a_25014_7093# a_24846_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12129 vssd1 a_20407_16519# _0540_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X12132 clknet_1_0__leaf_io_in[0] a_5341_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X12133 net80 a_16311_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12134 a_20690_3423# a_20522_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12136 dbg_result[0] a_7410_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X12137 a_7733_6409# a_6743_6037# a_7607_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12141 a_19609_28335# _0089_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12142 vccd1 _0728_ a_7289_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X12143 cal_lut\[181\] a_8971_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12144 a_1471_19319# _0422_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X12145 vccd1 net39 a_17415_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X12146 a_22041_16189# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12147 a_11742_5059# _0299_ a_11660_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12150 vccd1 a_15909_7809# _0546_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X12151 a_15611_1679# a_14913_1685# a_15354_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12152 vssd1 net34 a_24407_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12153 vccd1 a_1461_21781# _0763_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12154 temp1.capload\[13\].cap.Y net53 a_1861_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12155 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12156 _0061_ a_23671_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12157 a_3299_19061# _0744_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X12158 vccd1 a_21970_18231# _0490_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X12159 vssd1 net44 a_19991_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12160 a_27333_11477# a_27167_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12162 a_6546_26159# _0390_ a_6377_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X12163 a_21537_21807# a_21371_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12164 _0854_ a_20308_14441# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X12167 vssd1 a_26210_9951# a_26168_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12168 clknet_1_0__leaf_net67 a_3869_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12169 a_19694_5853# a_19421_5487# a_19609_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12170 vccd1 _0369_ a_10055_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12171 _0390_ a_2419_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X12174 vccd1 a_5399_8029# a_5567_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12175 vssd1 a_25439_9019# a_25397_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12176 a_8571_22895# _0748_ _0775_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X12178 a_9033_12559# cal_lut\[19\] a_8951_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12181 a_26693_21807# _0063_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12182 vccd1 a_5326_14709# a_5253_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12183 _0684_ a_21831_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X12184 vssd1 cal_lut\[88\] a_17417_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X12185 vccd1 cal_lut\[28\] a_18475_19783# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X12186 a_16986_25321# _0872_ a_16904_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12187 vssd1 net15 a_12160_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X12188 vccd1 net55 temp1.capload\[15\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12189 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12190 a_17888_25071# a_17489_25071# a_17762_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12191 a_25042_19605# a_24842_19905# a_25191_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12192 vccd1 cal_lut\[174\] a_25875_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12195 vccd1 clknet_0_temp1.i_precharge_n a_3882_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12197 a_14283_25437# a_14103_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12198 vssd1 a_27774_17567# a_27732_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12199 vssd1 a_14507_3855# a_14675_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12200 a_12621_5309# _0441_ a_12539_5056# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12201 vssd1 a_16807_11293# a_16975_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12202 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7012_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X12203 a_25011_14709# cal_lut\[68\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X12204 a_21538_26525# a_21291_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X12205 vccd1 _0759_ a_4892_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X12208 a_6863_29789# a_6081_29423# a_6779_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12211 a_7350_6005# a_7182_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12213 vccd1 net47 a_24407_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12214 vssd1 _0432_ a_5167_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X12215 a_13816_5487# cal_lut\[184\] a_13241_5633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X12216 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12217 a_13863_12559# a_13165_12565# a_13606_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12218 vssd1 net47 a_24407_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12219 _0347_ a_26519_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12220 a_26835_18909# a_25971_18543# a_26578_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12222 a_1765_30761# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12223 vccd1 a_21023_16885# a_20939_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12224 a_12258_20407# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X12225 vccd1 _0481_ a_12079_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X12226 vssd1 a_21115_21237# a_21073_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12227 a_7368_15113# a_6375_14741# a_7239_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X12228 vccd1 a_20451_23439# _0460_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X12229 vccd1 cal_lut\[166\] a_20499_8439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X12230 a_16355_29397# _0216_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X12231 vssd1 _0834_ a_4811_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12232 a_7381_28111# _0814_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12233 vssd1 a_27498_8863# a_27456_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12234 vccd1 a_4583_10615# cal_lut\[189\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12235 vccd1 _0252_ a_26063_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12236 vccd1 cal_lut\[11\] a_17814_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12237 cal_lut\[183\] a_10995_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12238 vccd1 a_2327_22895# _0418_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12239 vccd1 cal_lut\[143\] a_6187_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12240 a_20046_26677# a_19878_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12241 vssd1 _0747_ a_4997_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12242 vccd1 a_19793_21959# _0240_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X12243 vssd1 a_26946_21919# a_26904_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12244 a_18763_20871# _0485_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X12245 vccd1 a_20779_15253# _0851_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12247 _0804_ net22 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12248 a_10229_18793# net4 _0590_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12249 vssd1 a_17682_16100# a_17611_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X12250 vccd1 a_4647_12533# ctr\[4\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12251 _0429_ _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X12253 vssd1 a_1639_15444# _0199_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12254 a_3852_14165# _0411_ a_4075_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X12255 cal_lut\[136\] a_7131_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12256 vssd1 a_17935_28009# a_17942_27913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12257 a_13169_9295# _0099_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12258 a_6729_12559# _0018_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12259 vssd1 a_4647_12533# ctr\[4\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12261 a_9360_30663# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X12262 a_15745_25071# _0045_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12263 vccd1 _0422_ _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12264 vccd1 a_13882_4917# a_13809_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12265 a_14703_25236# _0272_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12266 vccd1 a_2060_30199# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X12267 a_7366_27613# a_6927_27247# a_7281_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12268 a_17428_2223# a_17029_2223# a_17302_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12269 cal_lut\[19\] a_7407_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12270 vccd1 net31 a_19255_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12271 vccd1 ctr\[8\] a_5227_26935# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X12273 a_16361_23777# _0481_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X12274 a_7936_22671# _0775_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X12275 vssd1 a_20119_28701# a_20287_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12276 vssd1 _0630_ a_10372_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12277 a_12361_21807# _0665_ a_12289_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12278 a_17410_16189# a_17095_16055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X12280 vssd1 _0392_ a_3799_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12281 a_7101_23439# _0437_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X12283 a_6963_5853# a_6265_5487# a_6706_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12284 cal_lut\[19\] a_7407_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12285 _0874_ a_20860_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X12286 clknet_0_io_in[0] a_6458_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12287 vccd1 _0840_ a_7387_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12288 vccd1 a_14733_15431# _0879_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X12289 a_17845_29423# a_17298_29697# a_17498_29397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X12290 vccd1 a_11287_27613# a_11458_27500# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X12291 a_10247_21583# _0630_ _0631_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X12292 a_24482_12559# a_24235_12937# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X12295 _0149_ a_16311_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12296 vccd1 a_8454_4917# a_8381_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12297 a_16025_12015# _0445_ a_15943_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12298 a_15285_28879# _0044_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12299 vssd1 a_20775_26311# cal_lut\[88\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12301 vccd1 _0663_ a_10596_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X12302 a_18765_20541# cal_lut\[58\] a_18693_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12303 _0662_ _0519_ a_9769_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X12304 _0201_ a_3799_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12305 vccd1 a_15727_21959# _0484_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X12307 a_6522_8863# a_6354_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12308 _0390_ a_2419_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X12310 vssd1 a_1407_10383# net4 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12311 a_21113_26525# a_20775_26311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X12312 a_12249_17455# _0005_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12313 vccd1 _0345_ a_25879_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12315 a_9692_4175# _0502_ a_9201_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12316 a_9763_27069# clknet_1_1__leaf__0380_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0567 ps=0.69 w=0.42 l=0.15
X12318 vccd1 cal_lut\[16\] a_14686_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12319 vccd1 net40 a_11711_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12320 cal_lut\[188\] a_7775_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12321 vccd1 dbg_result[3] a_15115_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=2.12 as=0.109 ps=1.36 w=0.42 l=0.15
X12322 a_26410_18909# a_26137_18543# a_26325_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12323 a_5227_26935# ctr\[7\] a_5461_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12324 a_23765_23759# _0466_ a_23355_23671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X12325 a_23513_8573# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12326 vssd1 net29 a_12815_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12327 a_27491_11092# _0357_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12328 cal_lut\[85\] a_21759_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12329 vccd1 _0706_ _0714_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12330 net25 a_9595_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X12332 a_22733_25437# a_22199_25071# a_22638_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12333 a_15105_22717# _0531_ a_15023_22464# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12334 a_26514_13077# a_26314_13377# a_26663_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12335 a_11874_3677# a_11435_3311# a_11789_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12336 a_4663_10205# a_3799_9839# a_4406_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12337 a_19071_11584# cal_lut\[186\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12338 a_5077_23983# _0429_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X12339 a_4435_32143# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X12340 vssd1 _0217_ a_17047_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12341 vccd1 _0334_ a_19439_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12342 vccd1 a_15503_7093# a_15419_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12343 a_24846_25437# a_24407_25071# a_24761_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12344 vssd1 a_6637_5175# _0318_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X12347 vccd1 a_12575_26703# a_12743_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12348 a_4069_25071# _0802_ a_3851_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X12349 a_22821_23817# a_21831_23445# a_22695_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12350 a_14917_21263# _0040_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12351 _0434_ _0421_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12352 vssd1 net34 a_17783_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12353 a_27621_13103# a_27351_13469# a_27531_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X12355 a_5451_10205# a_5271_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12356 vccd1 _0216_ a_21739_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X12357 a_25125_23445# a_24959_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12358 a_12171_12381# _0836_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12359 vccd1 _0447_ a_6391_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12360 vssd1 a_7239_12381# a_7407_12283# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12361 a_22103_3133# cal_lut\[153\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X12364 a_26141_6575# _0161_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12365 vccd1 a_8419_29691# a_8335_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12366 cal_lut\[179\] a_16147_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12367 vssd1 a_28199_11445# a_28157_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12368 _0395_ _0808_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12369 a_18961_25621# a_18795_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12370 vssd1 _0326_ a_6559_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12371 a_4333_10205# a_3799_9839# a_4238_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12373 a_14151_5652# _0300_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12374 a_22273_13103# a_22107_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12375 _0177_ a_16955_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12376 _0499_ a_9678_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X12377 vccd1 cal_lut\[188\] a_5451_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12378 a_25678_22173# a_25431_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X12379 a_15557_25071# a_15391_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12380 a_15128_21641# a_14729_21269# a_15002_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12382 a_11597_5487# a_10607_5487# a_11471_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12383 cal_lut\[163\] a_28015_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12385 vccd1 a_14875_24527# a_15043_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12386 vccd1 a_25271_7119# a_25439_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12387 vssd1 a_4831_10107# a_4789_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12388 vssd1 a_12035_26324# _0006_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12389 _0734_ _0724_ a_7755_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12390 vssd1 a_14155_3285# _0313_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X12391 a_3607_25935# clknet_1_1__leaf_temp1.i_precharge_n temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X12393 a_2099_18695# a_2371_18523# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12394 a_3607_20291# _0421_ a_3525_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12395 vssd1 a_20775_18231# _0526_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X12396 a_16753_16617# _0621_ a_16681_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12397 a_8562_14735# a_8123_14741# a_8477_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12399 _0272_ a_14283_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12400 _0032_ a_24591_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12401 cal_lut\[23\] a_17711_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12402 vccd1 _0465_ a_19071_11584# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X12403 vssd1 a_14875_24527# a_15043_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12404 vssd1 _0381_ _0192_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12405 _0183_ a_11987_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12406 a_9221_10089# _0699_ a_9125_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X12407 a_10325_7663# a_10055_8029# a_10235_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X12408 a_10677_11849# a_9687_11477# a_10551_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12409 vssd1 a_18027_19783# _0468_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X12410 vccd1 a_24499_9295# net36 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12412 _0477_ a_13751_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.331 ps=1.71 w=1 l=0.15
X12413 a_13592_7235# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12414 vccd1 cal_lut\[54\] a_21218_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12415 vssd1 _0310_ a_10331_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12416 vccd1 _0477_ a_16035_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X12417 vccd1 a_15519_23439# a_15687_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12418 a_24827_24501# cal_lut\[62\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X12419 a_26578_18655# a_26410_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12420 a_1773_22467# _0410_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X12421 a_15446_2741# a_15278_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12422 vssd1 a_14583_26677# a_14541_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12424 a_19862_24501# a_19694_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12425 a_2288_17973# net7 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X12426 vssd1 a_19583_2741# _0338_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X12427 vssd1 a_21978_21919# a_21936_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12428 vccd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12429 vssd1 a_15519_23439# a_15687_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12431 vssd1 _0637_ a_22441_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X12432 a_5460_15823# _0381_ a_5825_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12433 a_5871_10004# _0321_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12435 vccd1 _0235_ a_21279_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12436 a_9613_20693# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X12438 vssd1 a_4032_25847# _0829_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X12439 vccd1 a_1464_23957# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12440 a_6463_22057# _0431_ a_6245_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12442 a_10521_21263# _0627_ _0631_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12443 a_14277_13647# _0501_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X12444 vssd1 _0483_ a_9068_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X12445 vccd1 a_13403_25437# a_13571_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12446 a_7716_22325# _0434_ a_7936_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12447 a_12337_14191# a_12171_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12448 a_5353_28585# _0812_ _0402_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12449 a_12263_20495# _0447_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X12450 a_19915_19087# a_20132_19394# a_20090_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12451 a_14250_15797# a_14082_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12452 vccd1 a_27123_15431# cal_lut\[168\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12453 a_21073_21641# a_20083_21269# a_20947_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12454 a_19525_18543# _0442_ a_19437_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X12455 _0334_ a_18975_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12456 a_4713_21583# _0759_ a_4495_21495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X12457 vccd1 _0863_ a_24683_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X12458 a_17493_6575# _0112_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12459 vccd1 _0279_ a_14287_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12460 a_19694_24527# a_19421_24533# a_19609_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12461 a_27437_14191# a_27167_14557# a_27347_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X12462 vssd1 _0411_ _0428_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12463 a_27606_15823# a_27333_15829# a_27521_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12464 _0060_ a_21279_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12465 a_6587_16733# a_5805_16367# a_6503_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X12466 vccd1 a_2805_30265# a_2835_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12467 a_12163_29967# net14 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X12468 a_2209_25589# ctr\[3\] a_2462_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X12470 vssd1 _0752_ a_7389_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X12471 a_6611_22583# ctr\[12\] a_6737_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X12472 a_9385_4373# _0502_ a_9542_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12474 vccd1 net33 a_22843_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12475 vssd1 a_5399_8029# a_5567_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12476 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12477 vssd1 _0260_ a_13997_28023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12478 vccd1 a_19890_2197# a_19819_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X12479 a_8381_4943# a_7847_4949# a_8286_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12480 vccd1 a_22895_16519# _0689_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X12481 a_14082_15823# a_13809_15829# a_13997_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12482 a_14818_5853# a_14379_5487# a_14733_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12483 a_4593_8439# net24 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X12484 vssd1 a_21371_17455# net42 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X12485 vssd1 net30 a_11527_9303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12486 a_24306_12836# a_24099_12777# a_24482_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X12487 a_12575_26703# a_11711_26709# a_12318_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12488 a_2931_22325# _0744_ a_3362_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X12490 vssd1 a_17470_2335# a_17428_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12491 vccd1 net19 a_14287_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X12492 vccd1 clknet_0_io_in[0] a_5341_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12493 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12495 vssd1 a_8879_4917# a_8837_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12496 vccd1 a_20325_12533# _0538_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X12498 a_14979_24148# _0273_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12499 a_18187_1679# a_17323_1685# a_17930_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12500 vssd1 a_15715_5175# _0566_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X12501 a_10280_5059# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12503 vccd1 net47 a_24959_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12504 vssd1 a_10202_15797# a_10160_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12505 a_25783_6031# a_25603_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12506 a_7826_11293# a_7553_10927# a_7741_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12507 a_1735_27765# _0817_ a_1944_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X12508 vccd1 a_22863_8181# a_22779_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12509 a_1863_24233# _0414_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12510 vssd1 _0704_ a_9053_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X12511 _0572_ a_12079_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X12512 a_22806_25183# a_22638_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12513 _0424_ a_2722_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12514 a_24235_12937# a_24099_12777# a_23815_12791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X12515 a_12245_26703# a_11711_26709# a_12150_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12516 a_14156_11989# dbg_result[4] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X12517 vccd1 a_13771_21263# a_13939_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12518 a_17135_19087# a_16955_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12521 vccd1 _0237_ a_25235_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X12522 a_23841_14735# _0067_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12523 vccd1 a_13144_22325# _0863_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12524 vssd1 clknet_0__0380_ a_6537_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12525 a_22466_19605# a_22266_19905# a_22615_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12526 a_19789_11293# a_19255_10927# a_19694_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12527 vccd1 a_22806_25183# a_22733_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12528 a_22690_21263# _0638_ a_22441_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X12529 a_5100_7663# a_4701_7663# a_4974_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12530 a_19820_28335# a_19421_28335# a_19694_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12531 _0760_ a_4283_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X12532 vccd1 a_4484_32375# a_4435_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X12533 vssd1 clknet_1_1__leaf__0380_ a_7478_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X12535 a_21166_4765# a_20893_4399# a_21081_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12536 a_4624_15823# a_4351_15823# _0387_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12537 a_5644_12533# ctr\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.123 ps=1.07 w=0.42 l=0.15
X12538 _0197_ _0386_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12540 _0081_ a_12723_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12541 vssd1 a_21759_10107# a_21717_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12542 a_23021_16617# _0473_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X12543 vssd1 net29 a_9687_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12544 vccd1 a_21759_25339# a_21675_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12545 vssd1 a_10385_23413# _0681_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12546 a_18455_18337# _0464_ a_18369_18337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X12548 a_21166_11293# a_20727_10927# a_21081_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12550 vccd1 a_7527_15444# _0036_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12551 a_20223_15073# _0477_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X12552 vccd1 _0514_ a_14855_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12553 a_23723_25045# a_23899_25045# a_23851_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X12554 a_6611_22583# _0429_ a_6939_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12555 vccd1 _0363_ a_9411_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X12556 a_16097_7485# cal_lut\[138\] a_16025_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12557 a_13165_12565# a_12999_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12559 a_20267_9839# cal_lut\[108\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12560 vssd1 a_26911_16635# a_26869_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12561 vccd1 a_23811_4564# _0115_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12562 a_12000_3311# a_11601_3311# a_11874_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12563 vccd1 _0505_ a_15851_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12564 a_7741_29423# _0210_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12565 vssd1 a_14618_24501# a_14576_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X12566 a_15519_23439# a_14655_23445# a_15262_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12567 a_25839_14165# a_26123_14165# a_26058_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X12568 vssd1 a_3299_19061# _0745_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12569 a_21235_9514# _0284_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12570 vccd1 a_4406_9951# a_4333_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12572 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12573 vccd1 cal_lut\[30\] a_20942_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12575 vssd1 a_1921_11989# _0200_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12576 a_5323_4917# a_5499_5249# a_5451_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X12577 a_16574_17455# _0611_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X12578 vccd1 net1 a_3155_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X12579 _0196_ _0385_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12580 vssd1 cal_lut\[27\] a_24953_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12581 vccd1 a_26417_18231# _0247_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X12582 vssd1 cal_lut\[71\] a_26748_17705# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12583 a_7527_15444# _0880_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12584 a_25271_25437# a_24407_25071# a_25014_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12585 vccd1 _0857_ a_23763_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12586 a_11439_16367# _0625_ a_11302_16519# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X12587 a_14542_8029# a_14269_7663# a_14457_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12588 vccd1 cal_lut\[2\] a_8303_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12589 a_18269_8573# net19 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12590 vssd1 _0440_ a_17599_6039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12591 vccd1 cal_lut\[101\] a_15606_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12592 a_9131_2589# a_8951_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12593 a_13679_9295# a_12815_9301# a_13422_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12594 a_19694_24527# a_19255_24533# a_19609_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12595 _0757_ _0756_ a_3891_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12596 vccd1 a_19862_5599# a_19789_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12597 a_9542_4649# _0451_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X12598 vssd1 _0836_ a_6603_11777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12599 a_4789_11703# a_4885_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X12600 _0712_ _0708_ a_12265_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12601 a_15189_23439# a_14655_23445# a_15094_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12602 vccd1 cal_lut\[75\] a_25634_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X12604 a_5416_23413# _0820_ a_5545_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X12605 a_20569_16367# net18 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12606 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X12608 a_7255_20871# _0429_ a_7583_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12609 a_12502_17567# a_12334_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12610 a_18869_13647# a_18335_13653# a_18774_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12611 a_14139_28879# a_13441_28885# a_13882_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12612 ctr\[3\] a_3175_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12615 a_14151_4564# _0313_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12616 a_5554_19958# _0737_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X12617 a_15207_18543# dbg_result[1] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X12618 a_11579_3829# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X12619 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_6835_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12620 a_16692_27247# a_16293_27247# a_16566_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12621 _0061_ a_23671_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12622 _0839_ a_4167_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X12623 a_11671_2741# cal_lut\[147\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X12624 a_8478_19631# _0755_ a_8309_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X12625 vssd1 a_12691_10901# a_12698_11201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12626 _0528_ a_20267_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X12627 vssd1 a_4831_9019# a_4789_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12628 a_4963_10601# net27 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12629 a_7182_10383# a_6743_10389# a_7097_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12630 a_7366_27613# a_7093_27247# a_7281_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12631 vssd1 a_6947_9019# a_6905_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12632 vssd1 a_10827_3677# a_10995_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12633 vssd1 a_11195_28701# a_11366_28588# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X12634 vccd1 dbg_result[3] a_20690_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X12635 vssd1 a_8971_15797# a_8929_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12636 a_19807_14191# cal_lut\[12\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12637 a_8565_28879# a_8329_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X12638 cal_lut\[74\] a_28199_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12639 a_10294_11445# a_10126_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12640 a_10691_29423# net13 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X12641 vssd1 net81 a_16155_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X12642 a_14345_9269# _0564_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X12643 net5 a_1407_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12644 dec1.i_ones a_7959_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12646 vccd1 _0678_ a_10975_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12647 vssd1 a_12723_23439# net40 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12648 vccd1 _0454_ a_16035_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12649 vccd1 clknet_1_1__leaf_io_in[0] _0415_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12650 vssd1 a_2419_21807# _0414_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X12651 a_22201_18115# _0471_ a_22105_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X12652 a_27491_17130# _0250_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12653 a_26045_16367# a_25879_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12654 a_11609_8207# _0649_ a_11527_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12655 temp1.capload\[12\].cap.Y net52 a_1769_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12657 a_3128_31055# a_2879_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X12658 a_25891_20553# a_25762_20297# a_25471_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X12659 a_15009_29423# _0050_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12660 a_23377_19093# a_23211_19093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12661 _0555_ _0546_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X12662 vssd1 _0809_ a_4259_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12664 a_17187_13255# _0445_ a_17421_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12665 a_15933_8573# _0505_ a_15851_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12666 vccd1 a_12212_30199# a_12163_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X12667 a_7755_25321# _0721_ a_8055_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12668 a_25271_23261# a_24573_22895# a_25014_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12669 vccd1 cal_lut\[148\] a_13639_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12670 a_14541_27081# a_13551_26709# a_14415_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12671 vccd1 _0420_ _0737_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12673 a_2137_20719# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12674 vssd1 a_5583_14735# a_5751_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12675 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12676 vssd1 a_22843_9295# _0451_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12677 vccd1 _0448_ a_15023_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12678 vccd1 a_26026_8181# a_25953_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12679 a_7553_29423# a_7387_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12680 a_12265_24233# _0706_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12681 a_3983_8029# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12682 vssd1 _0483_ a_10761_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12684 vssd1 net44 a_18519_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12685 a_17762_1679# a_17323_1685# a_17677_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12687 a_15297_22895# _0486_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X12688 vssd1 cal_lut\[39\] a_11981_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12689 cal_lut\[48\] a_19827_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12690 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12691 a_14913_13653# a_14747_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12693 _0136_ a_3983_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12694 a_26307_13077# net37 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12695 vssd1 a_27003_18811# a_26961_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12696 a_12594_2335# a_12426_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12699 a_17065_3855# a_16727_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X12700 a_12299_3677# a_11601_3311# a_12042_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12701 vssd1 net36 a_25603_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12702 vccd1 a_22903_21959# _0463_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X12703 cal_lut\[48\] a_19827_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12704 a_23263_26935# a_23554_26825# a_23505_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X12705 vccd1 _0841_ a_9043_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X12706 a_14944_5487# a_14545_5487# a_14818_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12707 _0801_ _0800_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12708 a_12959_15253# a_13135_15253# a_13087_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X12710 _0509_ a_23151_10955# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X12711 _0472_ _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12712 a_9815_14557# a_9117_14191# a_9558_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12714 a_2804_20175# a_2750_20407# a_2722_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X12715 a_25271_7119# a_24407_7125# a_25014_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12716 a_27311_13879# a_27602_13769# a_27553_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X12717 vssd1 a_9201_3829# _0700_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X12718 a_12594_2335# a_12426_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12719 a_27245_8751# _0166_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12720 vssd1 cal_lut\[15\] a_23849_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12721 vccd1 a_12318_26677# a_12245_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12722 a_14243_16532# _0879_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12723 vccd1 net32 a_19715_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12724 _0633_ a_21831_9408# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X12725 a_20069_9295# _0107_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X12727 a_10975_20969# _0676_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12728 a_11521_13103# cal_lut\[21\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X12730 a_9595_5737# _0498_ a_9678_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X12731 a_8105_15829# a_7939_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12733 vccd1 a_12962_27359# a_12889_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12734 vccd1 a_23627_19796# _0026_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12735 vssd1 _0297_ a_23671_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12737 _0465_ a_21721_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.143 ps=1.33 w=1 l=0.15
X12738 _0588_ a_10832_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X12739 a_7553_6575# a_7387_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12740 net34 a_17415_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X12741 a_2489_8181# temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12742 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12743 vccd1 _0467_ a_12079_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X12744 vssd1 _0851_ a_19333_13255# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12745 _0185_ a_17231_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12747 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X12748 a_14156_11989# dbg_result[4] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X12749 vccd1 _0717_ _0718_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12750 vccd1 net25 a_12079_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12751 vccd1 net25 a_9963_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12752 a_1677_7663# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12753 vssd1 a_15904_25589# net45 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X12755 vssd1 _0229_ a_21463_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X12756 a_23627_19796# _0869_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12757 vccd1 a_19551_16885# a_19467_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12758 vssd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12759 vccd1 a_6427_11445# _0377_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X12760 _0438_ a_13459_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12761 _0344_ a_23943_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X12762 _0699_ a_9034_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X12763 a_7369_28879# a_7133_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X12764 vssd1 a_16187_23671# _0482_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X12765 a_18130_3677# a_17691_3311# a_18045_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12766 _0370_ a_11707_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X12767 a_24635_8513# _0341_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X12768 a_4912_8439# net39 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X12770 vssd1 a_11458_27500# dbg_result[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X12771 vccd1 a_17094_20407# _0587_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X12772 vssd1 a_7410_14709# a_7368_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X12773 vssd1 _0693_ a_9963_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12774 _0020_ a_9595_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12775 a_2377_28500# _0832_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12776 vssd1 _0635_ a_22383_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X12777 a_2582_14557# a_2309_14191# a_2497_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12778 temp1.dac_vout_notouch_ net14 a_11796_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X12779 vssd1 _0414_ _0801_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X12781 vssd1 net36 a_26891_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12782 vssd1 a_14031_12533# a_13989_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12783 a_25014_25183# a_24846_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12784 vssd1 a_14770_18517# _0472_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12785 a_7323_17999# a_6541_18005# a_7239_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X12786 vssd1 a_23231_25339# a_23189_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12787 vssd1 _0839_ _0194_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12788 vccd1 a_20963_15797# _0222_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12789 a_19287_21835# _0454_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X12790 _0297_ a_23344_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X12791 a_12233_7663# cal_lut\[142\] a_12161_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12792 net73 a_7475_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X12793 vssd1 net31 a_19899_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12794 vccd1 a_10839_15444# net12 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12796 vssd1 a_6244_25045# _0807_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X12797 a_26183_17821# a_25401_17455# a_26099_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12798 a_3759_21495# net21 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X12799 _0242_ a_21228_15529# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X12800 a_15680_12937# a_15281_12565# a_15554_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12801 vccd1 a_25014_25183# a_24941_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12802 vssd1 a_3685_22325# clknet_1_1__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X12803 a_23539_20407# a_23830_20297# a_23781_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X12804 vccd1 a_8951_31599# net10 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12805 a_14185_27497# cal_lut\[50\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X12807 a_1951_27023# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X12808 a_5412_19783# ctr\[2\] a_5554_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X12809 a_13087_15279# cal_lut\[96\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X12810 a_12092_7497# a_11693_7125# a_11966_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12811 a_27491_11092# _0357_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12812 a_18560_27497# _0260_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12813 _0381_ clknet_1_0__leaf__0380_ a_5639_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12814 a_22291_22895# _0466_ a_22469_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X12815 vccd1 net41 a_11895_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12817 vccd1 a_28031_12559# a_28199_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12818 vccd1 a_18475_18695# _0605_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X12819 _0099_ a_12723_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12821 a_26827_16733# a_26045_16367# a_26743_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12822 vccd1 a_26123_14165# a_26130_14465# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12823 a_18639_3677# a_17857_3311# a_18555_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12824 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12826 vssd1 a_22619_15253# net37 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X12827 vccd1 _0350_ a_25143_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12829 a_2700_25935# _0800_ a_2209_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12830 vccd1 _0450_ a_23395_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12831 _0720_ dec1.i_ones vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12832 vccd1 a_14307_28853# a_14223_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12833 vccd1 _0476_ a_9411_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12834 a_19889_22895# _0459_ a_19807_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12835 a_25156_18377# a_24757_18005# a_25030_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12836 a_2949_16201# a_1959_15829# a_2823_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12837 a_20775_5639# _0441_ a_21009_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12838 a_13441_28885# a_13275_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12839 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12840 vccd1 _0453_ a_18979_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12842 a_11506_15645# a_11067_15279# a_11421_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12843 _0668_ _0628_ a_11067_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12849 vssd1 _0591_ a_10247_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.127 ps=1.04 w=0.65 l=0.15
X12850 a_4899_5309# cal_lut\[137\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X12851 vccd1 a_27215_13879# cal_lut\[174\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12852 a_6449_3311# a_6283_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12853 cal_lut\[144\] a_7407_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12854 vccd1 a_12691_10901# a_12698_11201# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12855 vccd1 a_5143_11445# a_4885_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X12856 vccd1 _0445_ a_17507_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12857 a_9301_23145# _0704_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X12858 _0237_ a_12723_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X12859 _0519_ a_13052_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X12861 _0494_ a_10046_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X12862 a_22133_14013# _0474_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12864 _0535_ a_19255_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X12865 a_20421_9839# cal_lut\[108\] a_20349_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12866 vccd1 _0813_ a_5915_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12867 a_5553_25321# ctr\[7\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12869 a_21767_14557# a_20985_14191# a_21683_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12871 vccd1 a_10975_20969# _0679_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12872 a_3862_23439# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X12873 a_2417_17027# net6 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X12874 a_10129_15823# a_9595_15829# a_10034_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12875 a_22259_19605# net43 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12876 a_4988_32463# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X12877 vssd1 net23 a_6283_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12878 a_18482_12533# a_18314_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X12879 vssd1 a_18369_18337# _0475_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X12881 vccd1 _0817_ a_1765_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X12882 a_12472_5487# cal_lut\[129\] a_12352_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X12883 net47 a_16219_25623# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X12884 a_8397_24847# _0714_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X12885 a_11516_16617# _0609_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X12886 a_17888_2057# a_17489_1685# a_17762_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12887 a_11693_7125# a_11527_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12888 cal_lut\[100\] a_13847_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12889 a_20598_16885# a_20430_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12890 vccd1 a_6508_32375# a_6459_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X12891 vccd1 a_8383_22583# _0777_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X12893 a_6428_24501# _0437_ a_6820_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X12894 a_10635_11471# a_9853_11477# a_10551_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12895 _0228_ a_20308_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X12896 a_8024_31599# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X12897 vssd1 _0836_ a_3288_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12899 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12900 _0426_ _0422_ a_3425_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12901 a_11895_16617# _0625_ _0626_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12902 _0330_ a_12223_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12903 vccd1 a_25743_14343# cal_lut\[169\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12905 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12907 a_17871_3133# cal_lut\[155\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X12908 _0680_ _0520_ a_9423_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12909 a_20855_16911# a_20157_16917# a_20598_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12910 a_22523_2999# a_22619_2999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X12911 a_15370_17821# a_14931_17455# a_15285_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12912 _0081_ a_12723_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12913 a_3785_17999# _0422_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12914 _0012_ a_20635_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12915 a_20430_16911# a_20157_16917# a_20345_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X12916 a_5897_28335# a_5661_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X12918 vccd1 a_18015_5639# _0598_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X12919 vssd1 net9 a_9595_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12920 vssd1 net27 a_7387_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12921 net35 a_15812_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X12922 _0467_ a_15370_19407# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X12923 vccd1 a_18355_1653# a_18271_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12924 a_13301_7485# net17 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X12925 vssd1 a_15370_19407# _0467_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X12926 vccd1 _0465_ a_18645_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X12927 vccd1 a_23079_17607# _0480_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X12928 a_2049_21623# a_1857_21365# a_1963_21365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X12929 vccd1 a_23443_20407# cal_lut\[58\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12930 a_23155_6031# a_22291_6037# a_22898_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12931 a_20654_12559# _0536_ a_20574_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12933 a_7251_1898# _0373_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12934 vccd1 a_25927_10602# _0169_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X12936 a_24122_17188# a_23915_17129# a_24298_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X12937 a_15632_20291# cal_lut\[34\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X12938 vssd1 _0580_ a_17197_19777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X12939 a_7350_6005# a_7182_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12940 a_12127_21959# _0521_ a_12361_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12941 a_2524_16201# a_2125_15829# a_2398_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12942 vssd1 _0751_ a_6244_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X12943 vssd1 a_11587_8725# a_11594_9025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X12944 _0552_ a_16955_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X12945 _0740_ _0738_ a_4709_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X12946 vssd1 a_16727_4087# cal_lut\[178\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12947 vssd1 a_10719_11445# a_10677_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12948 _0191_ a_12815_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12949 a_8299_32463# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X12952 a_17217_2223# _0149_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X12953 vssd1 a_1743_18259# _0422_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12954 vccd1 a_21334_4511# a_21261_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12955 a_18878_9572# a_18678_9417# a_19027_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X12956 cal_lut\[171\] a_28199_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12958 clknet_0_temp1.i_precharge_n a_2778_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12959 a_7239_12381# a_6375_12015# a_6982_12127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12960 a_24051_17289# a_23915_17129# a_23631_17143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X12961 vccd1 a_25439_9019# a_25355_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12962 vssd1 net30 a_3707_9303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12963 _0697_ a_8758_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X12964 a_7826_11293# a_7387_10927# a_7741_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12965 a_14979_24148# _0273_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12966 a_18256_3311# a_17857_3311# a_18130_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12967 vssd1 cal_lut\[169\] a_25597_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12968 vccd1 a_22695_27791# a_22863_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12969 vssd1 _0461_ a_18765_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12970 vssd1 a_25594_5220# a_25523_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X12971 _0277_ a_11891_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X12972 vccd1 net9 a_9687_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X12973 a_2961_7663# net60 temp1.capload\[5\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12975 vssd1 io_in[0] a_6458_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12976 vssd1 _0260_ a_15469_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12977 a_14542_1501# a_14103_1135# a_14457_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12978 a_11969_3677# a_11435_3311# a_11874_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X12979 vssd1 a_11639_5755# a_11597_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12980 _0523_ a_19623_23552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X12981 a_7206_19087# a_7157_19319# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X12982 _0258_ a_12120_14851# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X12983 a_8546_1653# a_8378_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12984 vccd1 cal_lut\[72\] a_22983_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X12986 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12987 vssd1 cal_lut\[86\] a_23765_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X12988 cal_lut\[71\] a_28015_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12989 a_15177_22717# cal_lut\[93\] a_15105_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12990 vssd1 _0468_ a_23016_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X12991 a_28031_15823# a_27333_15829# a_27774_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12992 a_17029_2223# a_16863_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12994 _0088_ a_17231_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12995 vccd1 a_14710_7775# a_14637_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12996 vssd1 _0590_ a_10562_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X12997 a_6779_9117# a_5915_8751# a_6522_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X12998 a_24455_13255# a_24551_13077# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12999 a_19421_28335# a_19255_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13000 vssd1 net6 a_3155_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X13001 _0779_ ctr\[5\] a_5998_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X13002 _0090_ a_17875_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13003 _0747_ a_3072_19637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X13004 vssd1 _0504_ a_9779_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X13005 vccd1 a_13847_9269# a_13763_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13006 cal_lut\[119\] a_14307_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13007 vssd1 a_20046_26677# a_20004_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13008 vssd1 a_19977_14709# _0501_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X13010 a_25769_9839# a_25603_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13011 a_16550_11039# a_16382_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13012 vccd1 net36 a_27167_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13013 a_11796_30287# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13016 a_19793_21959# cal_lut\[64\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X13017 vssd1 _0876_ a_24591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13020 vccd1 a_2563_23957# _0824_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X13021 a_20372_22729# a_19973_22357# a_20246_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13022 a_6541_14741# a_6375_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13023 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4351_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13024 net76 a_6739_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X13025 vssd1 a_23110_3044# a_23039_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13026 a_7277_14191# a_7111_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13027 vccd1 a_9595_3311# net25 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13028 a_15637_8751# cal_lut\[126\] a_15565_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13029 a_17853_18377# a_16863_18005# a_17727_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13030 vccd1 _0487_ a_13649_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13031 vccd1 a_10746_10615# _0702_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X13032 a_26309_12015# a_25762_12289# a_25962_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X13033 a_8929_16201# a_7939_15829# a_8803_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13034 vccd1 dbg_result[3] a_14905_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X13035 a_2504_29423# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13037 a_21081_25071# _0084_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13038 a_22757_5309# cal_lut\[115\] a_22685_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13039 vccd1 a_28031_11471# a_28199_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13040 a_11292_30663# net8 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X13042 a_20303_26703# a_19605_26709# a_20046_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13043 a_3679_20291# _0422_ a_3607_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13044 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13045 a_20119_4765# a_19421_4399# a_19862_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13046 a_24679_22351# a_24499_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13047 vssd1 _0426_ _0427_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13048 a_23763_6031# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13049 a_9293_10089# _0698_ a_9221_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13050 a_2564_25045# _0806_ a_3246_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13051 a_10659_7637# net39 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X13052 a_21511_26159# a_21291_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X13053 _0802_ a_4984_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X13054 a_11759_4564# _0311_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13055 _0662_ _0433_ a_9687_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13056 a_12610_3855# a_12337_3861# a_12525_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13057 a_19694_11293# a_19255_10927# a_19609_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13058 a_24770_19631# a_24455_19783# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13059 vccd1 net18 a_22875_17249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13061 _0357_ a_27163_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X13062 vccd1 a_20451_23439# _0460_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13063 vccd1 _0451_ a_23763_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X13064 vssd1 _0341_ a_27211_8513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13065 a_25597_10749# a_25327_10383# a_25507_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X13066 a_6779_29789# a_5915_29423# a_6522_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13067 vccd1 a_19333_24135# _0261_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13068 a_18751_23671# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13069 vssd1 net31 a_17323_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13070 a_22185_1679# _0151_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13071 a_10126_13469# a_9853_13103# a_10041_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13072 a_17107_4073# net31 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13073 a_11671_2741# a_11847_3073# a_11799_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X13075 a_16293_27247# a_16127_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13076 a_3112_19783# _0420_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X13079 a_15991_8903# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X13080 _0210_ a_7557_28640# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X13081 vccd1 _0732_ a_10659_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X13082 vssd1 _0492_ a_10401_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X13083 a_14167_19783# _0442_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X13085 a_27024_17027# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13086 a_12955_3476# _0312_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13087 vccd1 a_23355_10615# _0696_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X13088 a_19255_3677# _0330_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13089 a_6449_29789# a_5915_29423# a_6354_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13090 a_17243_4233# a_17107_4073# a_16823_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X13091 vssd1 _0749_ a_7716_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X13092 a_8477_14735# _0078_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13093 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X13094 vccd1 a_18171_6843# a_18087_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13095 vccd1 net30 a_6007_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13096 cal_lut\[55\] a_22863_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13097 a_3981_14191# ctr\[2\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X13099 a_21810_16733# a_21371_16367# a_21725_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13100 a_14523_6549# cal_lut\[125\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X13101 a_8351_11777# _0863_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X13102 _0175_ a_25051_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13103 a_6429_28309# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X13104 vccd1 a_17105_10357# _0624_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X13105 vssd1 a_1736_18517# _0744_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X13106 a_4811_17705# _0446_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13107 a_24867_16733# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13108 _0851_ a_20779_15253# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13109 vssd1 a_8730_14709# a_8688_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13110 a_3338_27247# _0830_ a_2839_27221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X13111 a_21261_4765# a_20727_4399# a_21166_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13112 vssd1 a_13367_10391# _0260_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X13113 vssd1 a_10551_13469# a_10719_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13114 vccd1 a_6611_22583# _0788_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X13115 cal_lut\[124\] a_12559_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13116 a_5911_22057# _0429_ a_5693_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13117 _0110_ a_19807_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13118 a_2485_22351# net22 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13121 vccd1 cal_lut\[138\] a_5486_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X13122 vccd1 a_7239_12559# a_7407_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13123 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6835_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X13125 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13126 vssd1 _0177_ a_17661_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X13127 _0103_ a_20175_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13129 a_15921_29257# a_14931_28885# a_15795_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13130 a_22553_3855# _0115_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13131 vccd1 a_2489_8181# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13132 vssd1 a_10938_28471# a_10876_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X13133 a_23481_10383# _0506_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X13134 _0173_ a_27903_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13136 a_5555_24233# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X13137 a_5508_24501# _0431_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X13138 vccd1 net62 temp1.capload\[7\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13139 vssd1 a_7239_12559# a_7407_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13141 a_2447_19087# _0411_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13142 a_8335_9117# a_7553_8751# a_8251_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13143 a_10777_27247# _0196_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13144 a_17831_24746# _0220_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13145 a_19225_9673# a_18671_9513# a_18878_9572# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X13146 _0174_ a_26063_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13149 a_19999_19453# dbg_result[1] a_19915_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0567 ps=0.69 w=0.42 l=0.15
X13150 a_24630_10089# cal_lut\[170\] a_24473_9813# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13151 vssd1 a_23231_3829# a_23189_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13152 a_16949_3311# a_16679_3677# a_16859_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X13153 vssd1 a_18298_3423# a_18256_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13154 vccd1 a_16907_1985# a_16731_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13155 a_14223_4943# a_13441_4949# a_14139_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13156 vccd1 a_12597_7809# _0573_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X13157 vssd1 a_12575_26703# a_12743_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13158 vccd1 cal_lut\[31\] a_22649_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X13162 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13163 vssd1 clknet_1_1__leaf__0380_ a_9595_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X13164 a_14668_1135# a_14269_1135# a_14542_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13165 cal_lut\[190\] a_6487_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13166 vssd1 a_5751_14709# ctr\[6\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13167 vssd1 a_14131_13879# _0575_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X13168 a_16679_24527# _0484_ a_16761_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X13169 vccd1 a_22625_17973# _0643_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X13170 a_24591_6031# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13172 _0714_ _0706_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13173 a_9613_20693# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X13175 a_18698_19319# dbg_result[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X13178 _0784_ _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=2.1 w=0.65 l=0.15
X13179 a_10121_19631# _0667_ a_10037_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X13180 a_16823_4087# a_17107_4073# a_17042_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X13181 vccd1 _0505_ a_22291_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13182 a_23547_26921# net47 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13184 a_4068_31375# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13185 _0298_ a_19343_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X13186 a_12343_16617# cal_lut\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13188 a_7012_32463# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13189 clknet_1_1__leaf__0380_ a_8390_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13190 a_15289_18543# _0446_ a_15207_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X13191 a_12863_14954# _0275_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13192 _0825_ a_1735_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13193 a_24915_21959# a_25011_21781# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X13194 vssd1 _0439_ a_8979_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13195 a_6391_16911# clknet_1_0__leaf__0380_ _0382_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13196 ctr\[6\] a_5751_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13197 vccd1 a_7607_6031# a_7775_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13198 _0321_ a_5404_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13199 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6375_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13200 vccd1 cal_lut\[82\] a_17129_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X13201 vssd1 _0316_ a_6879_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13203 a_15725_15797# _0540_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13204 a_13161_4233# a_12171_3861# a_13035_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13205 vccd1 clknet_1_0__leaf_io_in[0] a_2143_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13206 vssd1 a_17927_4917# _0445_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X13208 vssd1 _0724_ a_7165_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.266 pd=2.12 as=0.091 ps=0.93 w=0.65 l=0.15
X13209 a_23926_14735# a_23653_14741# a_23841_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13210 vccd1 net45 a_18795_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13211 a_10570_1653# a_10402_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13212 a_4701_7663# a_4535_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13213 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_1407_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13214 a_6916_14735# a_6375_14741# a_6823_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X13216 vssd1 net36 a_22107_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13217 a_22277_14735# _0066_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
R31 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd_66.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X13218 a_17489_25071# a_17323_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13219 vssd1 a_20931_1653# a_20889_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13221 a_8001_29245# ctr\[11\] a_7929_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13222 vccd1 cal_lut\[33\] a_22872_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X13223 a_9312_30287# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13225 vccd1 _0421_ a_2742_18082# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X13226 a_15354_13621# a_15186_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13227 a_10129_3311# a_9963_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13228 a_6538_5853# a_6099_5487# a_6453_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13229 vssd1 _0421_ a_2099_18695# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13230 a_7618_26935# ctr\[12\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X13231 a_7921_26819# ctr\[12\] a_7849_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13232 a_4091_15529# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X13233 a_20141_6005# _0585_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X13234 vccd1 _0271_ a_13275_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13235 _0029_ a_19991_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13236 a_15524_11177# _0260_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13237 a_24551_13077# a_24835_13077# a_24770_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X13238 a_10454_22057# _0669_ a_10372_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13239 _0877_ a_24771_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X13241 vccd1 a_23899_25045# a_23723_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13242 a_23016_21583# cal_lut\[33\] a_22441_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X13244 _0289_ a_23804_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13245 a_3325_8903# cal_lut\[140\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X13246 _0449_ a_17907_10955# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X13247 a_9933_19061# _0628_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X13248 vccd1 a_16727_21482# _0041_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13249 a_17628_19881# _0579_ a_17526_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X13250 vccd1 a_22926_27221# a_22855_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X13252 _0099_ a_12723_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13253 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_6467_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X13254 a_7939_22895# _0724_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13255 a_27422_17999# a_26983_18005# a_27337_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13257 a_20513_20719# cal_lut\[54\] a_20441_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13258 a_7239_12559# a_6375_12565# a_6982_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13259 vssd1 a_24915_21959# cal_lut\[33\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13260 vssd1 a_5871_10004# _0138_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13261 a_22273_18115# _0480_ a_22201_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13262 vccd1 a_14795_5162# _0119_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13263 vccd1 _0285_ a_18795_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13264 a_5319_10749# a_5099_10761# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X13265 _0485_ _0447_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13266 vccd1 a_16147_3829# a_16063_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13267 a_2397_12937# a_1407_12565# a_2271_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13268 a_7891_5461# _0316_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X13269 vssd1 a_9678_29156# a_9607_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13270 a_5599_27221# a_5890_27521# a_5841_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X13271 a_16727_21482# _0214_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13272 a_8979_18543# _0433_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X13273 a_5165_3855# _0134_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13275 vssd1 a_25271_9117# a_25439_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13276 a_13459_2589# _0330_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13277 vccd1 _0221_ a_18519_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13278 a_8392_19631# _0765_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13279 _0151_ a_21463_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13281 a_24057_3855# a_23719_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X13282 a_13403_25437# a_12705_25071# a_13146_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13283 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X13284 a_22365_3861# a_22199_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13285 a_7553_6575# a_7387_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13286 _0282_ a_20032_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13287 vccd1 a_6428_24501# _0793_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X13288 vccd1 _0722_ _0765_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13289 vccd1 net20 a_17907_10955# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13290 vssd1 a_25042_19605# a_24971_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13291 vssd1 _0467_ a_16189_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13292 a_15177_8751# cal_lut\[132\] a_15105_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13293 _0047_ a_18519_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13294 vccd1 _0863_ a_11711_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X13295 a_9815_14557# a_8951_14191# a_9558_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13296 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_4435_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X13297 a_9406_29245# a_9091_29111# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13298 a_9223_24527# _0727_ a_9005_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13299 a_12162_5487# cal_lut\[183\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X13301 vssd1 cal_lut\[26\] a_23573_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13302 vccd1 a_22059_1109# a_21883_1109# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13303 a_15519_29789# a_14821_29423# a_15262_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13304 clknet_1_1__leaf_io_in[0] a_6182_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13305 vccd1 a_5341_17429# clknet_1_0__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13306 clknet_0_net67 a_3882_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13307 a_7452_31055# a_7203_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X13308 a_22895_16519# _0688_ a_23223_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13310 vccd1 a_8171_3476# _0132_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13311 _0280_ a_15524_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13312 a_9936_30761# a_9687_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X13313 vccd1 cal_lut\[14\] a_23207_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13314 vccd1 a_22633_11445# _0457_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X13315 a_8111_21583# _0627_ _0794_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X13316 vccd1 cal_lut\[65\] a_20298_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X13317 net42 a_21371_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13318 vccd1 a_23323_6005# a_23239_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13319 vccd1 cal_lut\[11\] a_17168_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X13321 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13322 vssd1 a_17415_7119# net34 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13323 vssd1 a_17841_12161# _0608_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X13324 _0229_ a_21136_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X13325 vccd1 _0500_ a_9033_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13326 a_9485_14557# a_8951_14191# a_9390_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13327 a_11343_13103# _0501_ a_11521_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X13328 a_14733_5487# _0119_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13329 vccd1 a_5412_19783# _0738_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X13330 a_17312_13967# cal_lut\[11\] a_16737_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X13331 vssd1 a_9021_29575# net71 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X13332 vssd1 cal_lut\[139\] a_6645_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13333 a_26551_10205# a_25769_9839# a_26467_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13334 a_8348_32375# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13335 vssd1 cal_lut\[103\] a_20032_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13336 vccd1 a_2099_18695# _0743_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X13337 vccd1 cal_lut\[110\] a_23757_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X13339 vssd1 _0679_ a_11756_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X13340 vccd1 a_12502_17567# a_12429_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13341 a_4277_23957# _0759_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X13342 a_15830_25437# a_15391_25071# a_15745_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13343 a_22079_5263# _0476_ a_21889_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X13344 cal_lut\[166\] a_26451_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13345 a_13514_21237# a_13346_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13346 a_7994_11039# a_7826_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13347 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13350 vssd1 ctr\[1\] a_4472_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13351 vssd1 net41 a_11895_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13352 a_2092_31287# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13353 vssd1 a_14710_1247# a_14668_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13354 a_6645_21583# _0432_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X13355 vssd1 _0589_ a_11067_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13356 vssd1 _0510_ a_23936_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X13358 a_10028_31055# a_9779_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X13360 vccd1 a_17401_24759# _0215_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13361 vssd1 _0427_ a_4616_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X13362 vccd1 a_9190_8181# a_9117_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13365 vccd1 _0505_ a_20267_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13366 a_21997_18543# dbg_result[2] a_21897_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13367 vccd1 a_6947_9019# a_6863_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13368 a_12445_10499# _0652_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X13369 a_22054_12559# _0476_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X13370 a_27517_17999# a_26983_18005# a_27422_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13371 a_14507_15823# a_13809_15829# a_14250_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13372 vccd1 a_10857_21781# _0675_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X13373 a_11609_10383# _0496_ a_11693_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13374 vccd1 _0316_ a_5271_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X13375 a_23481_10383# _0509_ a_23683_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13376 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13377 a_19609_24527# _0083_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13378 vccd1 _0664_ a_10413_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13379 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13380 a_17470_17973# a_17302_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13381 vccd1 a_10501_13879# _0257_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13382 _0368_ a_9131_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X13383 a_17841_12161# _0607_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X13384 a_26748_17705# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13385 _0308_ a_7980_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X13386 a_20154_9295# a_19715_9301# a_20069_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13387 a_11797_21379# a_11609_21379# a_11715_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13388 a_13968_17218# _0446_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13389 a_15703_2767# a_15005_2773# a_15446_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13390 a_20801_27791# a_20267_27797# a_20706_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13391 vccd1 _0032_ a_25849_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X13392 vssd1 _0489_ a_21970_18231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X13394 a_23573_18543# a_23303_18909# a_23483_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X13395 a_19509_17289# a_18519_16917# a_19383_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13396 vssd1 net25 a_15115_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13397 vccd1 a_27710_15253# a_27639_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X13399 vssd1 a_25962_20452# a_25891_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13400 vssd1 _0369_ a_10055_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13401 vccd1 a_5687_4564# _0134_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13402 vssd1 cal_lut\[170\] a_27253_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13403 a_7653_23439# _0728_ _0776_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X13404 vccd1 a_6927_16911# net48 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13405 a_2750_14303# a_2582_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13406 _0500_ a_16803_22689# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X13407 a_7583_20969# _0767_ a_7381_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13408 vccd1 a_12679_28010# _0007_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13409 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13410 vssd1 a_21023_16885# a_20981_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13411 vssd1 net8 a_10691_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X13414 a_17381_15425# _0551_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13415 vssd1 a_3007_14557# a_3175_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13416 a_6664_5487# a_6265_5487# a_6538_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13417 vssd1 _0746_ a_2700_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X13418 a_6445_10927# a_5455_10927# a_6319_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13419 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13420 a_6428_24501# _0750_ a_6648_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13421 vccd1 a_7410_17973# dbg_result[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13422 a_16911_29575# a_17007_29397# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13424 vccd1 net24 a_4259_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13425 vssd1 a_26514_13077# a_26443_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13427 vccd1 a_23723_25045# _0264_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X13428 vssd1 a_2419_21807# _0414_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13429 vccd1 net26 a_11527_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13430 vccd1 clknet_1_0__leaf__0380_ a_4816_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13431 vssd1 a_18659_10615# _0623_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X13432 vccd1 a_4963_10601# a_4970_10505# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13433 _0705_ _0704_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13434 vssd1 a_20690_18517# _0452_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.213 pd=1.3 as=0.0878 ps=0.92 w=0.65 l=0.15
X13436 a_4797_29423# _0208_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13437 vccd1 _0531_ a_19807_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13439 vssd1 _0840_ a_7387_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13442 vccd1 a_7791_27613# a_7959_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13444 a_13656_23817# a_13257_23445# a_13530_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13445 _0725_ _0712_ a_9301_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X13446 a_9779_11177# _0499_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13447 vssd1 _0701_ a_10746_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X13448 a_5779_8426# _0324_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13449 a_5099_10761# a_4963_10601# a_4679_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X13450 _0415_ clknet_1_1__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13451 vccd1 net40 a_14931_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13452 a_3695_23671# _0784_ a_3862_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X13453 _0248_ a_26748_17705# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13454 a_2014_12533# a_1846_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13457 cal_lut\[145\] a_7775_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13458 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13459 vssd1 _0746_ a_2137_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X13461 vccd1 a_11605_16055# _0844_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13462 a_15511_10383# a_14729_10389# a_15427_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13463 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_7452_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X13464 vccd1 clknet_1_1__leaf_io_in[0] a_7387_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13465 a_12533_26159# a_12263_26525# a_12443_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X13467 a_10603_23439# _0680_ a_10385_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13468 net20 a_14747_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X13469 vccd1 net45 a_21831_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13470 vccd1 a_14705_17620# net15 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13471 a_6909_6037# a_6743_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13472 a_7365_7497# a_6375_7125# a_7239_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13473 vssd1 _0715_ a_9967_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X13474 vccd1 a_6729_30199# _0404_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13475 a_4998_26165# ctr\[7\] a_4917_26165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X13476 a_21978_16479# a_21810_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13477 a_22530_14709# a_22362_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13478 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13479 vccd1 a_19659_25615# a_19827_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13480 vccd1 net29 a_14747_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13482 vssd1 a_19683_2197# a_19690_2497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13483 vccd1 a_4947_5249# a_4771_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13484 _0378_ a_12351_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X13485 vccd1 a_18763_20871# _0486_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
R32 temp1.capload\[9\].cap_64.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X13486 a_15538_28853# a_15370_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13487 vccd1 a_3575_15797# _0379_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X13488 vccd1 a_9558_14303# a_9485_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13489 a_17434_10383# _0622_ a_17354_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13490 cal_lut\[77\] a_17895_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13492 vccd1 _0446_ a_14103_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13494 vssd1 a_19659_25615# a_19827_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13495 vssd1 _0252_ a_26063_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13496 vssd1 a_23811_15431# _0656_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X13497 a_3149_22351# _0424_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X13499 a_3882_16911# net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X13500 _0023_ a_18611_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13501 vssd1 _0330_ a_19759_3073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13502 a_14703_25236# _0272_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13503 a_26536_18543# a_26137_18543# a_26410_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13504 cal_lut\[181\] a_8971_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13505 vssd1 net41 a_13643_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13506 a_16996_7235# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13508 a_4143_17999# a_3615_17999# _0429_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13509 a_7895_12778# _0861_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13510 a_20966_19743# a_20798_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13511 a_8803_1679# a_7939_1685# a_8546_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13512 a_21735_13469# a_21555_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13513 vccd1 _0676_ a_10975_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13514 a_25755_20393# net43 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13515 vccd1 a_22219_6843# a_22135_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13516 a_13146_25183# a_12978_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13518 _0547_ a_15483_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X13519 a_19421_28335# a_19255_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13520 a_19465_22895# _0465_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X13521 cal_lut\[31\] a_22403_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13522 a_22185_27791# _0054_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13523 a_19333_13255# cal_lut\[18\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X13524 vssd1 net19 a_21157_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13525 vssd1 a_5508_24501# _0796_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X13526 vccd1 _0753_ a_3891_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X13527 a_4609_29423# a_4443_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13528 a_4040_23759# _0789_ a_3850_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X13529 a_15243_5853# a_14379_5487# a_14986_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13530 vccd1 a_3877_11703# _0396_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13531 a_17475_16041# net44 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13532 a_1651_14165# ctr\[0\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X13533 a_1493_9615# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13534 a_16255_25437# a_15391_25071# a_15998_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13535 a_5418_13215# a_5250_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13536 vssd1 _0345_ a_25879_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13537 vccd1 a_27211_8513# a_27035_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13538 vssd1 a_7715_5461# _0328_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X13539 a_1573_12565# a_1407_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13540 a_17463_4221# a_17243_4233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X13541 vssd1 _0498_ a_11965_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X13542 vccd1 a_2419_21807# _0414_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X13543 dbg_result[0] a_7410_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X13544 vccd1 a_10551_11471# a_10719_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13545 _0446_ a_12815_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13546 a_3048_27247# a_3017_27399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X13547 a_3435_19407# _0424_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X13548 vccd1 a_14156_11989# _0440_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13549 vssd1 a_5675_13469# a_5843_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13550 vssd1 a_8546_1653# a_8504_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13551 a_14269_7663# a_14103_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13552 a_18222_28879# a_17783_28885# a_18137_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13553 vccd1 a_10075_6005# a_9991_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13554 vccd1 dbg_result[2] a_13459_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X13556 a_9871_3855# _0316_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13557 vccd1 a_20874_27765# a_20801_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13558 a_22954_17999# _0641_ a_22874_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13560 vssd1 _0500_ a_11781_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X13561 a_3067_22671# _0773_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X13562 vssd1 _0334_ a_19439_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13563 a_3848_24135# _0822_ a_3990_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X13564 vccd1 io_in[6] a_1407_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13565 _0568_ a_12539_5056# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X13566 a_4174_25981# _0759_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X13567 vssd1 _0751_ a_6428_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X13568 vccd1 _0264_ a_23763_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13569 a_21905_22173# a_21371_21807# a_21810_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13570 a_18045_3311# _0155_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13571 vccd1 a_4931_24135# _0798_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X13573 a_12705_22895# a_12539_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13574 vssd1 _0483_ a_15177_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13577 vssd1 a_13387_27515# a_13345_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13578 vccd1 _0742_ a_3299_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X13579 vccd1 a_14675_15797# a_14591_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13580 a_18249_5487# cal_lut\[155\] a_18177_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13581 a_18515_6031# a_18335_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13582 a_18170_12265# _0606_ a_18090_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13583 vssd1 a_9831_24501# _0727_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13584 a_6184_16367# a_5805_16367# a_6087_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X13585 a_13855_21263# a_13073_21269# a_13771_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13586 a_20280_9673# a_19881_9301# a_20154_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13587 a_26099_17821# a_25235_17455# a_25842_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13588 _0400_ a_5864_26819# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13589 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13590 a_6729_12015# _0190_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13591 vssd1 net26 a_14103_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13592 a_2043_31375# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X13593 a_22764_25071# a_22365_25071# a_22638_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13595 vccd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13596 net10 a_8951_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X13597 a_4897_20969# _0768_ a_5099_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13598 a_7826_29789# a_7387_29423# a_7741_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13599 a_19623_23552# cal_lut\[48\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13600 a_14151_5652# _0300_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13601 vssd1 a_22466_19605# a_22395_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X13602 a_21717_25071# a_20727_25071# a_21591_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13603 vssd1 a_21591_10205# a_21759_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13604 vssd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13605 a_5639_16911# _0425_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13606 a_11527_1679# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13607 a_3995_7497# a_3866_7241# a_3575_7351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X13608 a_13643_1679# _0363_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13609 a_9650_6005# a_9482_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13610 net33 a_23211_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X13611 a_16293_27247# a_16127_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13612 a_17857_3311# a_17691_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13613 vssd1 a_5843_9269# a_5801_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13614 a_12898_10901# a_12698_11201# a_13047_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X13615 a_20325_12533# _0537_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X13616 vccd1 _0853_ a_18151_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13617 vssd1 a_6706_5599# a_6664_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13618 net37 a_22619_15253# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13620 _0652_ a_11343_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X13621 vccd1 a_18187_24349# a_18355_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13622 a_9585_17999# _0516_ _0517_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X13623 a_20119_4765# a_19255_4399# a_19862_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13624 a_20893_4399# a_20727_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13625 a_2309_11791# ctr\[2\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13627 a_14369_22895# _0460_ a_14287_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13628 vssd1 net40 a_13275_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13629 a_10827_1679# a_9963_1685# a_10570_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13630 a_2447_19087# _0423_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13631 a_17191_16055# a_17475_16041# a_17410_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X13632 _0263_ a_21872_24643# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13633 vssd1 net10 a_7203_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13634 a_24099_4073# net33 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13635 _0311_ a_11660_5059# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13636 vssd1 a_13939_21237# a_13897_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13637 vssd1 net31 a_17691_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13638 vssd1 a_2947_10615# ctr\[2\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13639 vssd1 net48 a_16219_25623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13640 _0671_ a_11715_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
X13641 _0558_ a_18979_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X13642 a_18942_13621# a_18774_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13643 a_9568_31849# a_9319_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X13644 a_23147_25437# a_22365_25071# a_23063_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13646 a_3759_21495# _0446_ a_3885_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X13647 vccd1 _0481_ a_19623_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X13649 cal_lut\[104\] a_21759_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13651 a_8251_16733# a_7553_16367# a_7994_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13653 a_24653_12937# a_24099_12777# a_24306_12836# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X13654 vssd1 a_21115_3579# a_21073_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13655 vccd1 cal_lut\[119\] a_14651_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13656 a_11965_10703# cal_lut\[147\] a_11527_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13657 a_13629_28879# _0049_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13658 vccd1 _0465_ a_19807_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X13659 vccd1 a_22431_7338# _0158_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13660 a_10497_28335# a_10331_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13661 a_18187_24349# a_17489_23983# a_17930_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13662 vccd1 a_2317_16911# a_2417_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X13663 a_24235_4233# a_24099_4073# a_23815_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X13664 vccd1 net80 a_21095_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13665 cal_lut\[187\] a_7775_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13666 vccd1 a_8447_7338# _0126_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13667 a_15163_9527# _0440_ a_15397_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13669 _0015_ a_23763_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13670 vssd1 _0090_ a_18489_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X13671 _0462_ a_19255_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X13672 a_17095_5639# _0495_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X13673 a_1937_6549# clknet_0_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13674 vccd1 net54 temp1.capload\[14\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13675 clknet_1_0__leaf_net67 a_3869_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X13676 vccd1 a_11120_28853# net13 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13677 a_16404_17705# cal_lut\[101\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X13678 vccd1 a_2695_14013# _0808_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X13679 vccd1 a_15715_30186# _0044_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13680 vssd1 _0446_ _0448_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X13681 vssd1 a_10570_1653# a_10528_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13682 cal_lut\[107\] a_17711_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13683 vccd1 _0811_ a_5639_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X13685 a_25014_23007# a_24846_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13687 vccd1 net42 a_21371_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13688 a_9823_15041# _0237_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X13690 vssd1 a_19333_9991# _0285_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X13691 vssd1 cal_lut\[100\] a_14465_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13692 cal_lut\[7\] a_12743_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13693 io_out[4] a_1464_23957# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13694 vssd1 _0285_ a_18795_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13695 a_20690_21237# a_20522_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13696 _0375_ a_5451_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X13697 a_3288_11177# _0391_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13700 _0626_ _0625_ a_11895_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13701 a_18317_28879# a_17783_28885# a_18222_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13702 a_19973_26703# a_19439_26709# a_19878_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13703 _0453_ dbg_result[4] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13704 vccd1 _0472_ a_14287_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X13705 a_24351_14735# a_23653_14741# a_24094_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13706 _0184_ a_14379_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13707 vssd1 a_8454_4917# a_8412_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13708 vccd1 a_2376_30199# _0833_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X13709 _0446_ a_12815_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13710 a_4339_19407# _0428_ _0430_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X13711 vssd1 _0116_ a_24653_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X13712 vssd1 a_16373_13077# _0609_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X13714 a_18326_7637# a_18119_7637# a_18502_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X13715 a_9437_28157# _0815_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X13716 a_15377_19631# _0034_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13717 vccd1 cal_lut\[115\] a_22523_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X13718 a_19862_11039# a_19694_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13719 vccd1 a_7959_27515# a_7875_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13720 vssd1 cal_lut\[59\] a_19940_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13721 a_6464_25071# _0792_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X13722 vccd1 a_26651_6941# a_26819_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13723 a_14776_9295# _0492_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X13724 a_2778_24527# temp1.i_precharge_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13726 a_10083_24135# _0681_ a_10229_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X13727 a_13073_21269# a_12907_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13728 vccd1 a_8146_18796# dbg_result[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13729 vssd1 _0467_ a_12472_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X13730 vccd1 a_9179_28309# _0211_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.153 ps=1.3 w=1 l=0.15
X13731 a_10522_19958# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X13732 _0657_ a_21003_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X13733 a_5921_23145# _0776_ _0818_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X13734 vssd1 _0513_ a_9929_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X13735 a_7895_11690# _0881_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13736 _0599_ a_16035_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X13737 a_15998_25183# a_15830_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13738 a_22060_12879# _0452_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X13739 a_17691_27613# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13740 _0206_ a_6546_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X13741 a_20907_24527# a_20727_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13742 a_6847_21263# _0779_ a_6645_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13743 vssd1 a_28031_17821# a_28199_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13745 a_17033_14735# _0022_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13746 vccd1 a_21978_21919# a_21905_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13747 vccd1 a_7005_4551# _0315_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13748 a_17226_29423# a_16911_29575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13749 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13750 a_13537_15431# cal_lut\[78\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X13751 vssd1 a_17323_7663# _0505_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X13752 vssd1 a_2439_12533# a_2397_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13753 a_14604_13353# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13754 a_4003_30006# _0800_ a_3931_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X13755 a_25566_23413# a_25398_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13757 a_9956_31599# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X13758 a_5173_29199# a_4981_28940# _0208_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X13759 vccd1 a_22887_6549# a_22711_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X13760 _0392_ a_3288_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13761 a_17949_28885# a_17783_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13762 a_17302_17999# a_16863_18005# a_17217_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13763 a_22903_2985# net33 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13764 vccd1 a_12134_7093# a_12061_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13767 vssd1 _0453_ a_18519_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X13768 vssd1 _0502_ a_13816_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X13769 vssd1 a_4995_17999# net21 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13773 a_18291_9527# a_18387_9527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X13774 vssd1 a_27847_17999# a_28015_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13775 a_25743_5309# a_25523_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X13777 a_26690_13469# a_26443_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X13778 a_21954_25731# _0260_ a_21872_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13779 vssd1 a_20287_15547# a_20245_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13780 a_25463_12865# _0352_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X13781 vccd1 a_17875_16367# net44 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X13782 a_20985_14191# a_20819_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13784 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13785 vssd1 a_24455_13255# cal_lut\[16\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13787 a_25398_23439# a_25125_23445# a_25313_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13788 a_14457_1135# _0148_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13790 a_10126_11471# a_9853_11477# a_10041_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13792 a_8951_12559# _0501_ a_9033_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X13793 vssd1 a_27203_22173# a_27371_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13794 vccd1 a_21391_19899# a_21307_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13796 _0771_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13797 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_2504_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X13798 a_13052_15797# _0518_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13800 a_8268_24501# dec1.i_ones a_8491_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X13801 a_18611_20288# cal_lut\[58\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13802 a_15949_5309# cal_lut\[178\] a_15877_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13804 vssd1 a_21131_27791# a_21299_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13805 a_9547_20719# _0592_ a_9184_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X13806 a_21235_9514# _0284_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13807 vccd1 net42 a_24499_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13808 _0542_ a_15023_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X13809 _0223_ a_19664_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X13810 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13811 a_4678_26311# _0410_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.151 ps=1.35 w=0.42 l=0.15
X13812 a_11950_17999# _0574_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X13813 vssd1 clknet_1_0__leaf_io_in[0] a_6375_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13814 a_16250_9411# _0283_ a_16168_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13815 a_15189_19631# a_15023_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13816 a_25042_19605# a_24835_19605# a_25218_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X13817 a_16054_15823# _0541_ a_15974_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13820 vssd1 _0260_ a_15561_18231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13821 a_12426_2589# a_12153_2223# a_12341_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13822 a_6637_5175# cal_lut\[135\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X13823 a_15051_8029# a_14269_7663# a_14967_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13824 vssd1 a_6522_29535# a_6480_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13825 a_23811_27412# _0230_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13826 a_7733_2223# a_6743_2223# a_7607_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13827 vssd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13828 vccd1 a_13295_13371# a_13211_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13829 a_22886_11791# cal_lut\[176\] a_22796_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X13831 a_13303_27613# a_12521_27247# a_13219_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13832 vssd1 _0775_ a_8533_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X13833 vccd1 a_25363_15823# a_25531_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13834 a_20617_3677# a_20083_3311# a_20522_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13835 temp1.capload\[9\].cap.Y net64 a_1585_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13836 a_12245_12559# _0648_ a_12161_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X13837 vccd1 _0055_ a_23273_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X13839 a_27774_11445# a_27606_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13841 vssd1 _0159_ a_25389_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X13842 vccd1 a_16911_29575# cal_lut\[44\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13843 _0858_ a_14604_13353# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13844 vccd1 io_in[7] a_1407_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X13845 a_22971_13469# a_22107_13103# a_22714_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13846 _0427_ _0426_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13847 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5823_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X13848 _0595_ a_17231_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X13849 vccd1 a_5142_7775# a_5069_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13850 net5 a_1407_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13851 cal_lut\[32\] a_25439_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13852 a_6729_14735# _0192_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X13853 _0317_ a_5451_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X13854 vssd1 _0485_ a_20513_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13855 vccd1 _0461_ a_18611_20288# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X13857 vccd1 a_2221_13255# _0412_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X13859 a_16986_12559# _0603_ a_16737_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X13860 a_11030_27383# a_10871_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X13861 a_2778_24527# temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X13862 vssd1 _0436_ a_7111_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X13863 a_25523_5321# a_25394_5065# a_25103_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X13865 a_22641_13469# a_22107_13103# a_22546_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13866 vccd1 net45 a_16127_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13867 a_18502_8029# a_18255_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X13869 vccd1 a_6429_28309# _0209_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X13870 a_4245_14796# _0390_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X13871 vccd1 cal_lut\[15\] a_23759_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13872 net1 a_1407_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X13873 _0269_ a_17871_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X13874 vssd1 a_8711_4943# a_8879_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13877 a_27219_15253# a_27503_15253# a_27438_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X13878 a_8102_3855# a_7663_3861# a_8017_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13879 _0451_ a_22843_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13880 cal_lut\[49\] a_20471_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13881 vccd1 _0077_ a_18029_16201# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X13882 a_10783_30761# net13 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X13883 vccd1 ctr\[7\] a_4678_26311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X13884 vssd1 cal_lut\[61\] a_23389_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13885 vssd1 a_17095_10004# _0106_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13886 a_24206_20175# a_23959_20553# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X13887 a_20663_9295# a_19881_9301# a_20579_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13888 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13889 vssd1 cal_lut\[119\] a_14741_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13890 a_3362_22671# _0782_ a_3067_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X13891 vssd1 a_19551_16885# a_19509_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13893 a_10380_19783# dbg_result[5] a_10522_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X13894 _0195_ _0839_ a_5825_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13895 a_5599_27221# a_5883_27221# a_5818_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X13896 a_25398_23439# a_24959_23445# a_25313_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13897 vccd1 _0446_ a_4811_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13898 _0744_ a_1736_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X13900 a_27337_17999# _0070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X13901 vccd1 net16 a_12075_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X13902 a_7994_16479# a_7826_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13903 a_14243_16532# _0879_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13904 a_22988_4917# _0476_ a_23211_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X13905 _0434_ net7 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13907 a_7072_15797# net48 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X13908 _0393_ _0808_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13909 vccd1 a_8971_1653# a_8887_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13910 vssd1 _0443_ a_22445_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13911 a_17555_19319# _0474_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X13913 vssd1 a_23627_19796# _0026_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13914 vssd1 a_27590_17973# a_27548_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13915 a_15727_21959# _0464_ a_15901_21835# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X13916 a_17170_12265# _0851_ a_17088_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X13917 a_10784_23983# _0707_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X13918 a_7523_24833# _0724_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X13919 _0185_ a_17231_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13920 vccd1 a_15262_29535# a_15189_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X13922 ctr\[11\] a_8419_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13923 vccd1 _0865_ a_15575_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13924 a_12061_7119# a_11527_7125# a_11966_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13925 a_24630_10089# _0451_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X13926 vccd1 dec1.i_ones a_8951_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.18 ps=1.36 w=1 l=0.15
X13927 _0513_ a_9779_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X13928 vccd1 _0419_ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13929 vccd1 _0755_ a_5915_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X13930 vccd1 a_15411_5755# a_15327_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13931 a_10402_7119# a_10129_7125# a_10317_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X13932 vccd1 a_9687_29423# net9 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13935 _0050_ a_14747_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X13937 a_23627_19796# _0869_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13938 vssd1 net38 a_24499_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X13939 vccd1 _0411_ a_2447_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13940 vssd1 _0329_ a_9963_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13941 vccd1 temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13942 a_2518_30333# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X13943 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13944 vssd1 _0268_ a_18979_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X13946 a_25651_21807# a_25431_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X13947 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13948 vccd1 a_12959_15253# _0275_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X13949 a_25363_15823# a_24499_15829# a_25106_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X13951 a_26514_13077# a_26307_13077# a_26690_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X13953 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13954 a_2377_28500# _0832_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13955 temp1.capload\[2\].cap.Y net57 a_2413_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13956 _0089_ a_18979_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13958 a_14917_10383# _0100_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13959 vccd1 a_6319_11293# a_6487_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13960 ctr\[6\] a_5751_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13961 vssd1 a_23323_6005# a_23281_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13962 a_26309_12015# a_25755_11989# a_25962_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X13963 vssd1 a_11366_28588# a_11324_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X13964 _0371_ a_13823_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X13965 vccd1 _0351_ a_26615_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X13966 a_9235_25071# _0713_ a_9431_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13967 a_17029_18005# a_16863_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13968 a_20141_6005# _0583_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13969 vssd1 _0432_ _0767_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X13970 vssd1 a_17875_4399# _0290_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X13971 vssd1 a_12042_3423# a_12000_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X13972 a_25033_15823# a_24499_15829# a_24938_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X13973 a_26443_13103# a_26307_13077# a_26023_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X13974 vccd1 a_14655_18115# _0491_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X13975 vccd1 net7 _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13976 vccd1 _0167_ a_28057_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X13977 a_23389_23983# a_23119_24349# a_23299_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X13978 _0481_ a_12263_20495# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.327 ps=1.65 w=1 l=0.15
X13979 cal_lut\[131\] a_13203_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13980 _0611_ a_16035_18112# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X13981 a_26409_8585# a_25419_8213# a_26283_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13982 a_13989_12937# a_12999_12565# a_13863_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13983 _0020_ a_9595_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13984 vssd1 a_5507_22325# _0789_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13985 vccd1 a_3685_22325# clknet_1_1__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13986 vccd1 cal_lut\[5\] a_12343_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13987 a_8293_1679# _0180_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X13988 a_11869_21379# _0664_ a_11797_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X13989 a_25389_13103# a_24842_13377# a_25042_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X13990 a_22913_15113# a_21923_14741# a_22787_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13991 a_7994_29535# a_7826_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13992 a_25552_18793# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X13993 temp1.dac_vout_notouch_ net14 a_9312_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X13994 a_25011_14709# a_25187_15041# a_25139_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X13996 a_9033_12559# cal_lut\[79\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X13997 a_18597_13077# _0454_ a_18843_13131# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X13998 a_8335_13469# a_7553_13103# a_8251_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13999 a_23851_25071# cal_lut\[86\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X14001 vccd1 a_20417_13249# _0529_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14002 vccd1 net11 a_9319_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X14005 a_20387_28879# a_19605_28885# a_20303_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14006 vccd1 a_20287_4667# a_20203_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14007 a_14825_7119# _0125_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14008 a_19977_14709# _0477_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X14010 a_14821_29423# a_14655_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14011 vccd1 a_3882_22895# clknet_1_0__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X14012 cal_lut\[97\] a_13203_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14014 vssd1 a_11471_5853# a_11639_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14016 a_27521_15823# _0071_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14017 a_20203_15645# a_19421_15279# a_20119_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14018 a_17286_14709# a_17118_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14019 a_10570_3423# a_10402_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14020 vssd1 _0571_ a_12597_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X14021 a_15787_2767# a_15005_2773# a_15703_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14022 _0205_ a_4245_14796# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X14023 vccd1 a_10995_1653# a_10911_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14024 a_7994_6687# a_7826_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14025 a_9861_11177# _0512_ a_9779_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X14026 a_5060_32143# a_4811_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X14027 vccd1 a_19439_21263# _0459_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14029 a_19862_5599# a_19694_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14030 vssd1 _0839_ _0195_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X14031 vccd1 a_28015_7093# a_27931_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14032 vssd1 a_15469_20407# _0878_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X14033 vssd1 a_21971_13879# _0533_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14034 vccd1 a_22714_13215# a_22641_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14036 a_7097_2223# _0186_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14037 vssd1 _0481_ a_16925_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14038 vssd1 cal_lut\[130\] a_12625_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14039 vccd1 a_19763_28010# _0048_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14040 _0432_ a_6375_19095# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X14041 a_7994_6687# a_7826_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14042 cal_lut\[38\] a_8419_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14043 a_6453_5487# _0135_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14044 a_12443_26525# a_12263_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14045 vssd1 a_13146_23007# a_13104_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14047 a_7921_29789# a_7387_29423# a_7826_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14048 _0230_ a_21919_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X14050 vccd1 a_22695_1679# a_22863_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14052 a_1773_17027# net5 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X14053 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14054 vssd1 net23 a_7939_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14055 a_7097_10383# _0187_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14056 vssd1 a_18645_12043# _0502_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X14057 a_9761_15829# a_9595_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14059 vccd1 a_10832_30663# a_10783_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X14061 a_9221_14013# a_8951_13647# a_9131_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X14063 vssd1 _0614_ a_16390_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X14064 a_19402_25589# a_19234_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14065 a_7239_7119# a_6375_7125# a_6982_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14066 a_10413_20969# _0673_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X14067 a_24030_20452# a_23823_20393# a_24206_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X14068 cal_lut\[42\] a_17159_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14070 a_20249_21269# a_20083_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14071 vccd1 a_8730_14709# a_8657_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14072 vssd1 _0433_ a_8979_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14074 vssd1 a_4277_23957# a_4211_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X14075 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14076 _0252_ a_25552_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X14077 a_4395_25981# ctr\[1\] a_4032_25847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X14078 a_12276_27081# a_11877_26709# a_12150_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14079 a_8228_4233# a_7829_3861# a_8102_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14080 a_24358_10703# cal_lut\[163\] a_24268_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X14082 vccd1 _0339_ a_17415_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14084 a_25953_6575# a_25787_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14085 a_16991_22173# a_16127_21807# a_16734_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14088 a_18054_7663# a_17739_7815# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X14089 _0622_ a_16771_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X14090 a_19234_25615# a_18961_25621# a_19149_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14091 a_20296_13647# _0530_ a_20194_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X14092 vssd1 _0260_ a_12985_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14093 a_22567_26703# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14094 a_12127_21959# _0521_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14098 vssd1 a_6537_19605# clknet_1_0__leaf__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14099 a_2805_30265# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X14101 a_4128_20149# net21 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X14102 a_10317_1679# _0182_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14103 a_18440_12937# a_18041_12565# a_18314_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14104 a_23223_16617# cal_lut\[73\] a_23021_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14105 a_9364_4175# _0495_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X14106 _0737_ a_3799_19631# a_4180_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14107 vssd1 a_15722_12533# a_15680_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14108 a_3496_29967# a_3247_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X14109 a_16949_29245# a_16679_28879# a_16859_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X14111 _0708_ a_10784_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14112 a_16661_22173# a_16127_21807# a_16566_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14113 a_23299_14557# a_23119_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14115 a_8937_8207# _0121_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14116 vccd1 a_28199_12533# a_28115_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14117 vccd1 a_23063_3855# a_23231_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14118 a_8201_4943# _0145_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14120 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14121 a_19421_4399# a_19255_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14123 a_2552_31287# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X14126 _0407_ _0815_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14127 a_5093_23483# _0747_ a_4584_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X14128 clknet_1_1__leaf_net67 a_3685_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14129 a_12345_20495# a_12258_20407# a_12263_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
X14130 vssd1 cal_lut\[22\] a_14696_14441# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14131 a_24455_4221# a_24235_4233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X14132 _0336_ a_22471_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14133 a_26467_10205# a_25603_9839# a_26210_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14134 a_19537_22895# cal_lut\[89\] a_19465_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14135 a_10521_18793# _0589_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X14136 a_17996_13647# _0593_ a_17894_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X14137 vssd1 _0462_ a_22997_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14138 a_6277_24233# _0431_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X14139 a_15378_22895# cal_lut\[51\] a_15297_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X14140 a_1765_17455# net7 a_1683_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14143 _0485_ a_13942_20149# a_13722_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14144 vccd1 _0591_ a_9503_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X14145 a_9371_2741# cal_lut\[180\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X14146 a_7829_3861# a_7663_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14147 vssd1 _0718_ _0719_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14148 a_22395_19631# a_22259_19605# a_21975_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X14149 a_21825_18543# a_21555_18909# a_21721_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14150 vccd1 a_25106_15797# a_25033_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14151 a_11601_15645# a_11067_15279# a_11506_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14152 vccd1 _0363_ a_16679_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14153 vccd1 _0773_ a_4217_30006# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X14154 a_4951_7338# _0325_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14155 vccd1 _0630_ a_9671_21495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X14156 a_4484_32375# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X14157 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X14158 a_26137_10205# a_25603_9839# a_26042_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14159 a_5031_27791# a_4167_27797# a_4774_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14161 a_3115_10615# a_3406_10505# a_3357_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X14163 a_22077_21629# cal_lut\[87\] a_22005_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14164 vssd1 cal_lut\[134\] a_5541_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14165 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_3128_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14166 a_15473_27497# _0488_ a_15391_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14168 a_9190_8181# a_9022_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14169 a_23650_19087# a_23211_19093# a_23565_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14170 a_16493_17455# _0492_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X14171 a_10570_1653# a_10402_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14172 a_7281_27247# _0212_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14173 a_16635_26324# _0215_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14175 a_12686_1653# a_12518_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14176 vssd1 net20 a_21985_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14177 vccd1 _0817_ a_4351_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14178 a_10853_8573# cal_lut\[135\] a_10781_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14180 a_1464_23957# _0791_ a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14181 _0090_ a_17875_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14182 vssd1 a_10809_19605# a_10743_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X14183 a_9217_17999# cal_lut\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X14184 _0302_ a_7704_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X14185 a_4154_25321# _0799_ a_3851_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X14186 a_25007_5175# a_25103_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14187 a_8062_7235# _0299_ a_7980_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14188 _0278_ a_12259_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14189 _0241_ a_20216_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X14190 vssd1 a_19303_16519# _0606_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14192 vccd1 _0425_ a_13091_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X14193 clknet_0__0380_ a_7102_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14194 vssd1 _0550_ _0555_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X14195 a_5499_5249# _0316_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X14196 a_13606_12533# a_13438_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14197 a_22457_23145# cal_lut\[55\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14199 vccd1 _0347_ a_26799_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14201 vccd1 _0666_ _0670_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X14202 a_7718_18679# a_7559_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14204 a_27333_11477# a_27167_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14205 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_5060_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14206 a_17470_17973# a_17302_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14207 vssd1 a_13019_2491# a_12977_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14208 a_2224_12015# _0412_ a_1921_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X14210 a_8546_15797# a_8378_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14211 vccd1 a_12594_2335# a_12521_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14212 a_27163_10383# a_26983_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14213 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14215 _0441_ a_17560_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X14216 a_2209_25589# _0800_ a_2366_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X14217 a_10497_28335# a_10331_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14218 cal_lut\[137\] a_5291_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14219 vccd1 _0792_ a_6565_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14220 vccd1 a_24306_4132# a_24235_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X14224 a_11439_16367# cal_lut\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14225 vssd1 a_10075_6005# a_10033_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14226 a_15812_9269# net38 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X14227 vccd1 a_7994_29535# a_7921_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14228 a_20414_22325# a_20246_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14229 a_18137_28879# _0051_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14230 vssd1 a_7895_11690# _0037_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14231 vccd1 _0490_ a_9585_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
R33 vssd1 net60 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X14232 _0487_ a_16069_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X14233 vssd1 net42 a_21371_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14234 _0246_ a_24407_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X14237 _0207_ a_4705_27552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X14238 cal_lut\[154\] a_21759_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14239 a_8378_15823# a_8105_15829# a_8293_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14240 a_2689_7663# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14241 vccd1 cal_lut\[172\] a_14151_11079# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X14242 a_7239_12381# a_6541_12015# a_6982_12127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14243 cal_lut\[187\] a_7775_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14244 a_10827_1679# a_10129_1685# a_10570_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14245 a_19421_5487# a_19255_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14247 a_9126_10927# cal_lut\[38\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X14248 vssd1 _0801_ temp1.dac.vdac_single.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14249 vccd1 net41 a_12907_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14251 a_12943_1679# a_12245_1685# a_12686_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14253 vssd1 a_18390_28853# a_18348_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14254 a_3882_22895# clknet_0_temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14255 a_5089_19407# _0430_ a_4679_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X14256 vssd1 _0556_ _0557_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X14257 _0452_ a_20690_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14258 vssd1 a_1471_19319# _0423_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X14260 a_4351_31055# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14261 vssd1 a_7775_2491# a_7733_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14262 a_14710_7775# a_14542_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14263 _0577_ a_16679_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X14265 a_20246_22351# a_19973_22357# a_20161_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14266 vssd1 a_21426_14303# a_21384_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14267 a_19337_7663# _0505_ a_19255_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14269 a_2614_19631# _0762_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14271 a_25191_5487# a_24971_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X14272 a_7376_25935# _0722_ a_7073_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X14273 a_14686_20969# _0872_ a_14604_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14274 a_21591_2589# a_20893_2223# a_21334_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14275 a_18673_7663# a_18126_7937# a_18326_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X14276 _0198_ a_3851_15253# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14277 vssd1 a_11458_27500# a_11416_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X14278 vccd1 a_5675_3855# a_5843_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14279 a_2936_10089# net3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X14280 a_23754_26980# a_23554_26825# a_23903_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X14281 vssd1 a_4593_8439# a_4406_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X14282 a_8758_10383# cal_lut\[37\] a_8675_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14283 a_14875_24527# a_14011_24533# a_14618_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14284 a_24835_19605# net43 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14286 _0445_ a_17927_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14287 _0231_ a_22747_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X14288 vccd1 a_3759_21495# _0782_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X14289 a_8749_8213# a_8583_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14290 a_12535_4765# a_12355_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14291 a_12955_3476# _0312_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14292 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X14293 a_18795_1679# _0330_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14294 vccd1 _0445_ a_16035_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14295 a_15829_27247# cal_lut\[44\] a_15391_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14296 vssd1 a_22339_27399# cal_lut\[56\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14297 a_15427_10383# a_14563_10389# a_15170_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14298 a_13363_24349# a_13183_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14299 a_15522_23145# _0644_ a_15208_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X14301 temp1.dac_vout_notouch_ net66 a_3496_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14302 vccd1 a_16734_21919# a_16661_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14303 a_22638_3855# a_22365_3861# a_22553_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14304 a_15278_2767# a_14839_2773# a_15193_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14305 a_9650_6005# a_9482_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14306 a_3869_11989# clknet_0_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14308 a_11579_25045# _0708_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X14309 _0175_ a_25051_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14310 vccd1 a_2947_10615# ctr\[2\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14312 a_14545_24527# a_14011_24533# a_14450_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14313 vssd1 a_18383_5175# _0541_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14314 a_10416_30511# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X14315 a_16859_3677# a_16679_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14316 vccd1 dbg_result[2] a_15370_19407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X14317 _0236_ a_23299_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14318 a_22054_12559# cal_lut\[13\] a_21897_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14319 a_20579_8029# a_19881_7663# a_20322_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14320 a_15097_10383# a_14563_10389# a_15002_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14321 a_26259_14191# a_26130_14465# a_25839_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X14322 a_28031_10205# a_27333_9839# a_27774_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14323 a_25690_20541# a_25375_20407# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X14324 a_9423_18793# _0517_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X14325 vssd1 net30 a_6007_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14327 a_15538_28853# a_15370_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14328 a_22821_28169# a_21831_27797# a_22695_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14329 a_2900_20175# _0422_ a_2804_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X14330 a_5759_13469# a_4977_13103# a_5675_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14331 a_15991_8903# _0514_ a_16225_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X14332 a_9360_30663# net10 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X14333 a_4253_19087# _0427_ _0430_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14335 _0149_ a_16311_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14336 vccd1 a_25755_20393# a_25762_20297# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14337 vccd1 _0839_ a_6651_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14338 vccd1 a_11674_15391# a_11601_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14339 vssd1 cal_lut\[129\] a_11660_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14340 vccd1 a_10570_7093# a_10497_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14341 vccd1 cal_lut\[98\] a_10360_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X14342 _0584_ a_20175_5056# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X14343 a_20893_9839# a_20727_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14344 _0062_ a_24683_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14345 vccd1 net37 a_21923_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14346 vccd1 a_28199_11445# a_28115_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14347 _0835_ a_4187_28918# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X14348 a_24941_25437# a_24407_25071# a_24846_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14349 vccd1 _0750_ a_5921_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14350 vssd1 a_28199_15797# a_28157_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14351 a_15662_19407# _0442_ a_15548_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.137 ps=1.07 w=0.65 l=0.15
X14352 a_22438_23413# a_22270_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14353 vccd1 a_19333_9991# _0285_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X14354 vssd1 _0814_ a_6729_30199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14355 vssd1 _0271_ a_13275_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14356 vccd1 a_2419_21807# _0414_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14358 a_9209_6037# a_9043_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14359 clknet_0_temp1.dcdel_capnode_notouch_ a_2489_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14360 a_13714_28879# a_13275_28885# a_13629_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14361 vccd1 a_23055_23047# _0470_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X14362 a_25387_5161# net33 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14363 vccd1 net26 a_14379_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14364 vccd1 _0441_ a_14287_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14366 a_15354_13621# a_15186_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14367 a_15370_28879# a_15097_28885# a_15285_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14370 cal_lut\[41\] a_15595_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14371 vssd1 a_17475_16041# a_17482_15945# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14372 a_13783_24148# _0849_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14373 a_14737_18115# _0442_ a_14655_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X14375 vccd1 dbg_result[5] _0592_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14377 vccd1 _0467_ a_12539_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X14378 vccd1 clknet_1_0__leaf_io_in[0] a_1407_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14379 vccd1 a_6458_20175# clknet_0_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14380 a_7826_16733# a_7553_16367# a_7741_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14381 a_6266_27613# a_6019_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X14382 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14384 a_22270_23439# a_21997_23445# a_22185_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14385 a_16117_6397# _0445_ a_16035_6144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14386 _0440_ a_14156_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X14387 _0174_ a_26063_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14388 _0418_ a_2327_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14389 vssd1 a_14795_5162# _0119_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14390 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14391 vssd1 _0475_ a_17956_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X14392 a_12521_2589# a_11987_2223# a_12426_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14394 a_15186_13647# a_14913_13653# a_15101_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14395 a_21334_4511# a_21166_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14396 a_5073_6031# _0137_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14397 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X14398 vccd1 a_10202_15797# a_10129_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14399 vssd1 a_23719_12791# cal_lut\[15\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14400 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14401 _0363_ a_11579_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14402 vssd1 a_15991_8903# _0548_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14404 a_11151_29673# net13 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X14405 vssd1 a_9190_8181# a_9148_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14406 a_23719_12791# a_23815_12791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14407 a_9142_19958# _0433_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X14409 vssd1 net48 a_17875_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X14410 a_21334_4511# a_21166_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14411 a_13144_22325# _0838_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X14412 vssd1 cal_lut\[77\] a_17456_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14413 vccd1 a_7888_32375# a_7839_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X14416 a_25397_22895# a_24407_22895# a_25271_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14417 vccd1 a_15135_1403# a_15051_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14418 a_6651_18793# _0383_ _0194_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14419 net41 a_7072_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X14420 _0384_ clknet_1_0__leaf__0380_ a_4811_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14421 a_24953_19453# a_24683_19087# a_24863_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X14422 vssd1 _0351_ a_26615_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14423 a_12079_9295# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14424 vccd1 net10 a_7663_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X14425 a_14913_1685# a_14747_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14426 a_17118_14735# a_16845_14741# a_17033_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14427 cal_lut\[21\] a_10719_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14428 a_20746_13353# _0527_ a_20666_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X14429 a_1972_15113# a_1573_14741# a_1846_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14430 a_23815_12791# a_24099_12777# a_24034_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X14431 vssd1 net8 a_11151_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X14432 vssd1 net45 a_16127_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14433 a_18455_26525# a_17673_26159# a_18371_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14434 a_21905_16733# a_21371_16367# a_21810_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14435 a_14633_4233# a_13643_3861# a_14507_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14437 vssd1 _0608_ a_16373_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X14438 vccd1 a_4167_16367# _0839_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14439 a_12693_5309# cal_lut\[136\] a_12621_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14440 vssd1 net10 a_7011_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X14441 vccd1 a_10380_19783# _0667_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X14443 a_20249_9295# a_19715_9301# a_20154_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14444 a_7534_27359# a_7366_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14445 a_19496_25321# cal_lut\[47\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X14446 vssd1 a_7256_21237# _0778_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X14447 vssd1 _0417_ a_1764_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X14449 a_17217_17999# _0076_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14450 a_14369_8573# _0441_ a_14287_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14451 vccd1 a_16983_23047# _0578_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X14452 vccd1 a_16727_4087# cal_lut\[178\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14453 vssd1 a_27123_15431# cal_lut\[168\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14454 vccd1 a_1651_14165# _0411_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14456 vccd1 _0418_ a_2447_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14458 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_5547_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X14459 vccd1 net25 a_12171_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14460 cal_lut\[124\] a_12559_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14461 vssd1 a_17470_17973# a_17428_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14462 a_21009_15101# cal_lut\[66\] a_20937_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14463 vssd1 _0548_ a_15541_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X14464 cal_lut\[60\] a_21391_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14465 a_18501_13653# a_18335_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14466 _0630_ a_9933_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X14467 a_10697_19203# _0628_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X14468 vccd1 a_25594_5220# a_25523_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X14469 vccd1 a_12310_10615# _0660_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X14470 a_25042_5461# a_24842_5761# a_25191_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X14471 cal_lut\[9\] a_13571_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14472 a_18085_22923# _0464_ a_17999_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X14473 _0401_ net74 a_5639_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14474 vccd1 _0665_ a_11014_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X14475 a_18709_18543# cal_lut\[59\] a_18637_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14476 vssd1 cal_lut\[152\] a_22561_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14477 vccd1 a_7407_7093# a_7323_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14478 vccd1 a_13955_23439# a_14123_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14479 a_12463_20495# _0438_ a_12345_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.143 ps=1.09 w=0.65 l=0.15
X14480 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4068_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X14481 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_1951_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X14482 cal_lut\[7\] a_12743_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14483 a_15693_23983# _0481_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X14484 vssd1 a_2023_19319# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14485 a_20690_18517# a_20543_18543# a_21331_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X14486 _0593_ a_16771_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14487 vccd1 a_3007_14557# a_3175_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14488 a_12702_13469# a_12429_13103# a_12617_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14489 vccd1 _0216_ a_23119_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14491 cal_lut\[92\] a_15687_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14492 vccd1 net39 a_3339_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X14493 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_10239_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X14494 a_15511_21263# a_14729_21269# a_15427_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14495 vccd1 a_6503_16733# a_6674_16620# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X14496 vccd1 _0713_ a_8397_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X14497 vccd1 a_14618_24501# a_14545_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14498 io_out[4] a_1464_23957# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X14499 vssd1 a_13955_23439# a_14123_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14500 a_10372_22057# _0669_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14501 a_4882_29789# a_4443_29423# a_4797_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14502 vssd1 net25 a_11435_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14503 a_7840_31375# net10 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X14504 a_22695_23439# a_21997_23445# a_22438_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14506 a_21878_17143# _0684_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X14508 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14509 vccd1 a_8146_18796# a_8059_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X14510 a_16891_11293# a_16109_10927# a_16807_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14511 vssd1 a_9471_29097# a_9478_29001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14512 a_1461_21781# _0414_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X14513 _0448_ _0438_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X14514 vccd1 _0352_ a_26891_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14515 vssd1 net45 a_15391_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14516 a_15404_3145# a_15005_2773# a_15278_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14517 a_25191_13103# a_24971_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X14518 vssd1 a_5617_15431# net77 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X14519 a_10857_21781# _0521_ a_11110_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X14520 vccd1 cal_lut\[178\] a_15715_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X14521 a_28031_12559# a_27333_12565# a_27774_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14522 a_14155_3285# a_14331_3285# a_14283_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X14523 vccd1 a_14155_29397# _0224_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X14524 a_22790_11471# _0452_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X14525 a_21218_23145# _0222_ a_21136_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14526 a_2747_18517# _0423_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X14527 a_26137_18543# a_25971_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14529 cal_lut\[137\] a_5291_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14530 vccd1 a_12955_3476# _0130_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14531 vssd1 a_18371_26525# a_18539_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14532 vssd1 a_8171_3476# _0132_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14533 a_18606_9661# a_18291_9527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X14534 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_2879_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X14537 _0304_ a_10235_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X14538 vssd1 _0330_ a_22059_1109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14539 _0497_ a_9126_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X14540 vssd1 a_7255_20871# _0768_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X14541 vssd1 a_4128_20149# _0761_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X14542 ctr\[10\] a_6947_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14543 _0429_ _0421_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14544 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14545 a_19570_20969# _0558_ a_19256_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X14546 a_13291_18909# _0438_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X14547 a_9563_28487# ctr\[12\] a_9737_28363# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X14548 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_1959_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X14549 a_22872_21263# _0468_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X14551 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14552 dbg_result[2] a_8146_18796# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X14553 vccd1 cal_lut\[17\] a_17170_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X14554 _0734_ _0724_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.0878 ps=0.92 w=0.65 l=0.15
X14555 vccd1 _0421_ _0434_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14556 vssd1 a_7607_6031# a_7775_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14557 a_2777_14013# ctr\[0\] a_2695_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X14558 vccd1 a_4487_13077# _0204_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.153 ps=1.3 w=1 l=0.15
X14559 _0691_ a_16679_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X14560 a_19711_3133# cal_lut\[154\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X14561 a_10126_11471# a_9687_11477# a_10041_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14562 vssd1 net47 a_24959_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14563 vssd1 cal_lut\[181\] a_9692_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X14564 a_7715_5461# cal_lut\[145\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X14565 a_6090_27221# a_5883_27221# a_6266_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X14566 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14567 _0425_ a_7631_17171# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14568 cal_lut\[54\] a_21299_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14569 a_15632_26819# cal_lut\[91\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X14570 a_27311_13879# a_27595_13865# a_27530_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X14572 a_9516_14191# a_9117_14191# a_9390_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14574 a_23585_8573# cal_lut\[117\] a_23513_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14575 a_6645_21263# _0778_ a_6847_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14577 _0362_ a_25047_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14579 a_15005_2773# a_14839_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14580 vssd1 a_14163_8903# _0493_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X14581 vccd1 a_11200_29575# a_11151_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X14582 a_25931_8725# a_26107_8725# a_26059_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X14583 a_11014_22057# _0671_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X14584 a_7381_20719# _0432_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X14585 a_9000_19783# _0447_ a_9142_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X14586 vssd1 _0438_ a_13551_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X14587 a_6019_27247# a_5883_27221# a_5599_27221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X14589 a_4713_23805# _0797_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X14590 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14592 a_24065_18543# net18 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X14594 a_5517_10761# a_4963_10601# a_5170_10660# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X14595 vssd1 _0457_ a_21003_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14596 a_13165_12565# a_12999_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14597 vssd1 _0459_ a_20451_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
R34 temp1.capload\[15\].cap_55.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X14598 vssd1 io_in[4] a_1407_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X14599 a_6363_23983# _0720_ _0797_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X14600 a_22365_25071# a_22199_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14601 vssd1 a_25566_23413# a_25524_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14602 vssd1 _0777_ a_7256_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X14603 cal_lut\[150\] a_17895_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14604 vccd1 _0292_ a_18519_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14605 a_12815_26525# _0841_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14606 a_18111_25589# net47 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X14607 a_7741_29423# _0210_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14608 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14609 a_9371_2741# a_9547_3073# a_9499_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X14610 vssd1 _0784_ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14611 vccd1 _0711_ _0714_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14612 a_23355_23671# _0470_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X14613 vccd1 a_10197_25223# _0733_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X14614 a_6548_21807# _0410_ a_6245_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X14615 a_14703_21972# _0213_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14616 vccd1 dbg_result[3] a_12815_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X14617 _0056_ a_23395_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14618 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14619 vccd1 a_21978_16479# a_21905_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14620 vssd1 _0839_ a_9179_28309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14621 vssd1 a_22714_13215# a_22672_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14622 vssd1 a_25363_15823# a_25531_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14624 vccd1 cal_lut\[50\] a_14375_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14625 vccd1 a_14151_11079# _0567_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X14626 a_24835_13077# net36 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14627 a_3113_22923# _0410_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X14628 vssd1 _0508_ a_23237_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X14629 a_12978_25437# a_12705_25071# a_12893_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14630 a_16991_22173# a_16293_21807# a_16734_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14631 vccd1 a_22438_1653# a_22365_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14632 vccd1 clknet_0_net67 a_3685_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14633 _0444_ a_20943_6369# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X14634 _0326_ a_6187_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14635 a_4818_25398# _0747_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X14636 vccd1 _0453_ a_18027_19783# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X14637 a_14829_27247# cal_lut\[7\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X14638 dbg_delay clknet_1_0__leaf_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14639 a_17858_15823# a_17611_16201# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X14640 a_5508_24501# _0793_ a_5728_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14641 _0658_ a_23395_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14642 a_17117_21807# a_16127_21807# a_16991_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14643 vssd1 _0424_ a_4811_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14645 _0693_ a_9411_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14646 a_3081_28309# _0419_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X14647 a_13219_27613# a_12355_27247# a_12962_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14648 a_17956_15279# cal_lut\[78\] a_17381_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X14649 a_21031_3677# a_20249_3311# a_20947_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14650 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14651 a_15959_18793# _0491_ _0492_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14653 vccd1 a_8879_4917# a_8795_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14654 a_25953_6575# a_25787_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14655 temp1.capload\[15\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14657 vssd1 dbg_result[1] a_19057_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X14659 a_24793_13469# a_24455_13255# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X14660 a_16955_25615# _0266_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14662 a_9929_10357# _0494_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X14663 vccd1 _0420_ a_3679_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X14665 a_4963_10601# net27 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14667 vssd1 a_12950_16988# _0455_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X14668 vccd1 a_13882_28853# a_13809_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14669 a_10129_7125# a_9963_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14671 a_16069_22923# _0464_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X14672 vssd1 clknet_0_io_in[0] a_5341_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X14673 a_7347_24501# a_7523_24833# a_7475_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X14675 vccd1 a_10562_19319# _0666_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X14676 a_19605_28885# a_19439_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14677 vccd1 net47 a_21831_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14678 vccd1 net61 temp1.capload\[6\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14679 a_4583_10615# a_4679_10615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14680 net6 a_1407_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14681 vccd1 a_7131_5755# a_7047_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14682 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X14684 cal_lut\[49\] a_20471_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14685 vccd1 a_15262_27765# a_15189_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14686 _0086_ a_23763_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14687 _0875_ a_23391_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14688 a_25137_11837# a_24867_11471# a_25047_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X14689 clknet_1_0__leaf_temp1.i_precharge_n a_3882_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14690 a_6246_16503# a_6087_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14691 vssd1 a_12778_14303# a_12736_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14692 a_15009_29423# _0050_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14693 a_25603_6031# _0341_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X14694 a_21215_27791# a_20433_27797# a_21131_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14695 a_21081_25071# _0084_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14697 vssd1 a_14705_17620# net15 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14698 vccd1 a_8390_23439# clknet_1_1__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14699 vccd1 a_22806_3829# a_22733_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14700 a_21334_11039# a_21166_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14701 a_3081_28309# _0419_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X14702 a_16209_5309# _0514_ a_16127_5056# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14704 vssd1 _0616_ a_16390_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X14705 a_24455_13255# a_24551_13077# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14706 a_27521_9839# _0170_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14707 _0101_ a_16035_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14708 a_22438_27765# a_22270_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14709 _0531_ a_17783_21271# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X14710 vccd1 a_12851_2589# a_13019_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14711 vccd1 a_7631_17171# _0425_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X14712 a_25757_10927# a_25203_10901# a_25410_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X14713 _0625_ a_16373_16341# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X14714 vssd1 a_19862_4511# a_19820_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14715 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10416_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X14716 _0000_ a_1867_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14718 a_17538_16617# _0246_ a_17456_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X14719 vssd1 a_24075_19087# a_24243_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14721 vccd1 a_16731_9813# net38 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X14722 a_21978_21919# a_21810_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14723 vccd1 a_13241_5633# _0569_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14724 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_2149_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14725 a_28157_16201# a_27167_15829# a_28031_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14726 vssd1 a_20947_3677# a_21115_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14727 vssd1 clknet_0_io_in[0] a_6182_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14728 vccd1 cal_lut\[100\] a_14375_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14729 vccd1 a_5050_29535# a_4977_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14730 clknet_1_0__leaf_io_in[0] a_5341_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14731 _0306_ a_13592_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X14732 vssd1 _0222_ a_19057_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14733 vssd1 a_11471_14557# a_11639_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14737 a_9471_29097# clknet_1_1__leaf_io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14738 vccd1 ctr\[6\] a_5093_23483# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X14739 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X14740 a_5451_5309# cal_lut\[136\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X14741 vccd1 _0668_ _0670_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14742 vssd1 a_14675_15797# a_14633_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14743 vssd1 _0699_ a_9043_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X14744 vccd1 a_8251_29789# a_8419_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14745 a_17853_2223# a_16863_2223# a_17727_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14746 vssd1 a_25439_25339# a_25397_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14747 _0591_ _0590_ a_10521_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14748 a_5871_19958# _0736_ a_5412_19783# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X14749 a_15462_19997# a_15023_19631# a_15377_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14750 _0668_ _0590_ a_11149_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X14751 a_13508_18517# dbg_result[1] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X14753 a_25471_20407# a_25755_20393# a_25690_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X14754 clknet_1_0__leaf__0380_ a_6537_19605# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14755 a_19421_24533# a_19255_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14757 vssd1 _0495_ a_16097_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14758 temp1.dac_vout_notouch_ net14 a_9936_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14759 a_1656_26703# a_1407_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X14760 a_1837_17455# net5 a_1765_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14761 a_7895_12778# _0861_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14762 a_1863_24233# net22 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=2.79 as=0.135 ps=1.27 w=1 l=0.15
X14764 a_7475_24893# _0728_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X14765 a_14273_15431# cal_lut\[36\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X14766 _0424_ a_2722_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14768 a_14415_26703# a_13717_26709# a_14158_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14770 vccd1 clknet_1_1__leaf_io_in[0] a_10423_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14771 a_15285_17455# _0095_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14772 a_27606_12559# a_27333_12565# a_27521_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14773 vssd1 a_12723_21807# _0237_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X14774 a_21897_18543# dbg_result[1] a_21825_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X14775 a_4313_17429# _0741_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X14777 a_20429_27081# a_19439_26709# a_20303_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14778 vccd1 cal_lut\[89\] a_19303_23047# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X14779 cal_lut\[182\] a_9983_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14780 a_13796_19407# a_13459_19087# a_13714_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14781 a_15097_28885# a_14931_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14782 vccd1 a_9555_25847# _0721_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X14783 a_5687_4564# _0317_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14784 vssd1 a_3882_16911# clknet_0_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14785 a_22365_1679# a_21831_1685# a_22270_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14786 vssd1 _0465_ a_22077_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14787 a_5915_20175# ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X14788 a_26138_20175# a_25891_20553# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X14789 _0712_ a_11896_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X14790 vssd1 _0446_ a_13459_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X14791 a_6814_12381# a_6541_12015# a_6729_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14792 vssd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14794 a_1769_6351# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14796 a_1753_26133# clknet_0_temp1.i_precharge_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14797 a_2709_19407# _0423_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X14799 vccd1 _0056_ a_24101_27081# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X14800 vccd1 _0316_ a_6007_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14801 a_20690_18517# dbg_result[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.327 ps=1.65 w=1 l=0.15
X14802 _0520_ _0519_ a_9217_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X14803 _0545_ a_15851_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14804 a_11207_8903# a_11303_8725# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14805 a_26023_13077# a_26314_13377# a_26265_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X14806 a_13783_24148# _0849_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14807 vssd1 _0487_ a_17312_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X14809 _0491_ a_14655_18115# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X14810 vccd1 a_25455_17999# a_25623_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14811 a_2271_14735# a_1407_14741# a_2014_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14812 vccd1 _0173_ a_28149_14025# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X14813 vccd1 ctr\[7\] a_5946_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X14814 vccd1 cal_lut\[178\] a_15479_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14815 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_4528_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X14817 a_11195_28701# a_10331_28335# a_10938_28471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14819 a_23535_17143# a_23631_17143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14820 a_11046_5853# a_10773_5487# a_10961_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14821 ctr\[9\] a_5475_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14822 a_9821_21583# _0557_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X14823 a_22695_27791# a_21831_27797# a_22438_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14824 vccd1 ctr\[3\] a_4798_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X14825 _0602_ a_16127_20288# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14827 a_14637_7125# a_14471_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14828 a_7665_20719# _0766_ a_7255_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X14829 vssd1 _0853_ a_18151_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14831 vccd1 _0291_ a_19807_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14832 vccd1 _0672_ _0710_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X14834 a_4997_23805# a_4714_23483# a_4584_23671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14835 a_18823_12559# a_18041_12565# a_18739_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14836 a_9429_28879# a_9091_29111# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X14837 a_15163_9527# net20 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X14839 vssd1 a_9275_28023# _0816_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14840 a_19605_26709# a_19439_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14841 vssd1 _0797_ a_5365_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X14842 vccd1 a_5418_3829# a_5345_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X14843 vssd1 a_20451_23439# _0460_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X14844 a_8485_23145# _0724_ _0775_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14846 _0594_ a_17507_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14847 vccd1 a_6982_14709# a_6916_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X14848 a_20119_15645# a_19255_15279# a_19862_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14849 vssd1 a_24835_5461# a_24842_5761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14850 vssd1 a_17187_13255# _0601_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14852 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14853 a_23849_16367# a_23579_16733# a_23759_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X14854 a_22747_26703# a_22567_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14855 a_22365_27791# a_21831_27797# a_22270_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14856 vccd1 a_19308_17973# _0508_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X14857 vssd1 a_7631_17171# _0425_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X14858 cal_lut\[130\] a_12467_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14859 a_3420_12879# _0395_ a_3117_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X14860 _0459_ a_19439_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X14861 a_19881_13353# _0529_ a_19797_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X14862 cal_lut\[2\] a_8419_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14863 a_25891_12015# a_25755_11989# a_25471_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X14864 vssd1 a_7102_21807# clknet_0__0380_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14865 a_22733_3855# a_22199_3861# a_22638_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X14866 a_5525_7663# a_4535_7663# a_5399_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14867 vssd1 _0813_ a_5915_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14868 _0706_ a_10607_24640# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X14869 vssd1 a_26486_16479# a_26444_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14870 a_9126_11177# _0496_ a_9126_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X14871 a_3335_12559# _0396_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14872 vssd1 a_23818_19061# a_23776_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14873 a_9190_8181# a_9022_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14874 cal_lut\[158\] a_22219_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14875 vccd1 a_8251_11293# a_8419_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14876 a_22319_22173# a_21537_21807# a_22235_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14877 vssd1 a_25743_14343# cal_lut\[169\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14879 vssd1 a_26635_10107# a_26593_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14881 a_7194_28335# _0814_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X14882 temp1.capload\[4\].cap.Y net59 a_1953_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14885 vccd1 a_6537_19605# clknet_1_0__leaf__0380_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14886 a_3479_7351# a_3575_7351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14887 a_15469_12559# _0016_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X14889 a_22438_8181# a_22270_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14890 vccd1 cal_lut\[40\] a_14686_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X14891 a_9953_19631# _0669_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14892 vccd1 net41 a_9595_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14893 a_10699_8751# cal_lut\[141\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14895 _0618_ a_18611_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X14896 a_2668_30761# a_2419_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X14897 a_5050_29535# a_4882_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14898 vccd1 net38 a_16679_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14899 vssd1 a_24459_8181# _0349_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X14900 a_5809_10927# _0189_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14901 vccd1 a_13203_14459# a_13119_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14902 vssd1 a_10108_4373# _0316_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X14903 a_2009_30676# _0831_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14905 _0329_ a_10051_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14906 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd _0746_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14907 vccd1 net40 a_12539_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14908 vssd1 net23 a_8583_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14909 vccd1 _0306_ a_13183_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X14910 vccd1 a_3656_25847# a_3607_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X14911 vccd1 _0421_ _0737_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14912 vccd1 a_12525_18231# _0846_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X14913 vccd1 a_3882_16911# clknet_0_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14914 vccd1 _0341_ a_23855_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14915 cal_lut\[123\] a_10995_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14916 a_14967_8029# a_14103_7663# a_14710_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14918 a_17229_20291# _0577_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X14919 a_23063_3855# a_22365_3861# a_22806_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14920 vccd1 clknet_0_temp1.dcdel_capnode_notouch_ a_1937_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14921 a_14313_10927# _0474_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X14922 net45 a_15904_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X14923 vssd1 a_7607_10383# a_7775_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14924 vccd1 a_2722_20175# _0424_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X14925 vssd1 net80 a_21095_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14926 vccd1 a_8419_6843# a_8335_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14927 a_12870_13215# a_12702_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14928 vssd1 _0838_ a_12723_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X14929 a_13751_17277# _0425_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X14930 a_20506_1653# a_20338_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14932 vccd1 a_21591_25437# a_21759_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14933 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd a_2024_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14934 a_12985_10615# cal_lut\[97\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X14935 vccd1 a_14415_26703# a_14583_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14936 a_23151_10955# _0460_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X14937 vccd1 a_17841_12161# _0608_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14938 vccd1 net40 a_14655_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14939 vccd1 _0665_ a_12127_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X14940 vssd1 a_21721_18909# _0465_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X14941 a_10129_9295# cal_lut\[97\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14943 vssd1 a_6779_9117# a_6947_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14944 a_12065_26703# _0006_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14945 a_7291_10205# a_7111_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14946 a_10029_11177# _0499_ a_9957_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X14947 vssd1 _0719_ a_9773_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X14948 a_10423_26703# _0839_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14949 vccd1 _0679_ _0682_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14950 clknet_0_net67 a_3882_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14951 vccd1 a_2933_14709# _0202_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X14952 a_7251_1898# _0373_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14953 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ a_1937_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14954 a_11207_8903# a_11303_8725# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X14956 a_1860_17271# a_1673_16911# a_1773_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X14957 vssd1 a_8546_15797# a_8504_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14958 vssd1 a_15623_15431# _0549_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X14959 a_12778_3829# a_12610_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14960 a_4771_4917# cal_lut\[137\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X14961 vccd1 _0836_ a_4903_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X14962 a_4180_19631# _0421_ a_3990_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14963 a_22383_18793# _0639_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X14965 vccd1 _0666_ _0676_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14966 a_14131_13879# cal_lut\[16\] a_14277_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14967 a_19325_14025# a_18335_13653# a_19199_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14968 a_25455_17999# a_24591_18005# a_25198_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14969 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd a_1656_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X14970 a_8419_25071# _0713_ a_8229_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14971 vccd1 net8 a_10975_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X14973 cal_lut\[75\] a_25623_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14974 vssd1 a_5278_12533# net72 vssd1 sky130_fd_pr__nfet_01v8 ad=0.186 pd=1.26 as=0.208 ps=1.83 w=0.42 l=0.15
X14975 a_13403_23261# a_12539_22895# a_13146_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X14976 vssd1 _0420_ a_3995_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X14978 vccd1 cal_lut\[187\] a_7291_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14979 vssd1 a_15078_7093# a_15036_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X14980 vssd1 a_14153_20884# net17 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X14981 _0842_ a_8303_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X14983 vssd1 a_27923_9019# a_27881_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14984 _0850_ a_10699_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X14985 a_17118_9295# a_16845_9301# a_17033_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X14986 _0125_ a_14195_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X14987 a_14696_14441# _0851_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14988 a_19819_2223# a_19683_2197# a_19399_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X14989 a_27521_17455# _0073_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X14990 a_22503_24135# cal_lut\[61\] a_22649_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14992 a_11674_15391# a_11506_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X14993 vssd1 cal_lut\[177\] a_16949_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14994 a_10875_31599# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X14995 vssd1 _0482_ a_17025_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X14996 vssd1 net23 a_9043_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X14997 _0353_ a_27347_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X14998 a_10551_13469# a_9853_13103# a_10294_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14999 a_13722_20175# _0425_ a_13525_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15000 a_17217_2223# _0149_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15001 a_13073_23261# a_12539_22895# a_12978_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15002 a_20763_1679# a_20065_1685# a_20506_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15003 a_26743_16733# a_25879_16367# a_26486_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15004 a_25322_5309# a_25007_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X15005 a_14917_21263# _0040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X15006 a_21997_8213# a_21831_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15007 a_23653_14741# a_23487_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15008 a_23344_4649# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15009 a_9454_4175# cal_lut\[133\] a_9364_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X15010 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_1407_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X15011 vssd1 a_8251_13469# a_8419_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15012 a_9673_23047# _0716_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X15013 a_11950_18319# _0587_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X15014 a_17291_29397# net45 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15015 a_23886_8323# _0283_ a_23804_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15016 a_6519_21495# ctr\[11\] a_6645_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X15018 a_27606_11471# a_27333_11477# a_27521_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15019 vssd1 a_4584_23671# _0822_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X15020 a_11067_19407# _0590_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X15021 vccd1 a_7111_17455# _0437_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15022 a_21878_17143# _0689_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X15023 a_7786_8323# _0299_ a_7704_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15024 a_6445_29111# a_6541_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X15025 a_19694_15645# a_19255_15279# a_19609_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15026 a_5345_3855# a_4811_3861# a_5250_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15027 vssd1 _0431_ a_6375_19095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X15028 a_5389_27069# _0811_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X15029 a_19149_25615# _0047_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X15030 _0239_ a_25415_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X15031 vccd1 _0453_ a_18243_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15032 a_12541_10499# _0654_ a_12445_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15036 _0772_ a_1963_21365# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X15037 vccd1 a_2014_14709# a_1941_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15038 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15039 a_17630_15529# _0553_ a_17381_15425# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X15040 vccd1 a_4310_8439# a_4259_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X15041 clknet_1_0__leaf__0380_ a_6537_19605# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15042 _0249_ a_26012_15939# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X15043 a_12778_3829# a_12610_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15044 a_25042_5461# a_24835_5461# a_25218_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X15045 vssd1 _0465_ a_19961_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15046 clknet_0_io_in[0] a_6458_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X15047 a_17470_2335# a_17302_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15048 vccd1 a_22438_27765# a_22365_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15049 vccd1 net24 a_4719_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15050 vssd1 a_21879_16055# _0551_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X15051 vssd1 net36 a_27167_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15052 a_5264_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X15054 a_13529_25071# a_12539_25071# a_13403_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15055 vccd1 _0707_ a_11142_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15057 _0865_ a_14696_14441# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X15058 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ a_1477_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15059 a_10232_30287# net8 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X15060 _0448_ a_14167_19783# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X15061 vssd1 _0438_ _0439_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15062 vccd1 a_23719_4087# cal_lut\[117\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15064 a_23811_27412# _0230_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15065 _0399_ _0811_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15066 a_7071_25045# _0734_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X15067 a_16158_21379# _0872_ a_16076_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15068 a_15538_17567# a_15370_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15070 vccd1 a_4771_20871# _0770_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X15072 vssd1 a_7315_3579# a_7273_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15073 a_2823_15823# a_1959_15829# a_2566_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15074 vccd1 a_19303_2375# cal_lut\[155\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15075 vccd1 a_20683_21972# _0065_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15076 a_14415_26703# a_13551_26709# a_14158_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15077 a_14565_13967# _0456_ a_14131_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X15078 a_5801_13103# a_4811_13103# a_5675_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15079 vssd1 net20 a_20421_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15080 a_19333_25223# _0872_ a_19496_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X15081 a_23200_18319# cal_lut\[75\] a_22625_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X15082 vccd1 a_7350_10357# a_7277_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15084 a_17772_19631# cal_lut\[34\] a_17197_19777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X15085 a_5667_14735# a_4885_14741# a_5583_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15086 a_14910_7119# a_14471_7125# a_14825_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15087 vssd1 net11 a_9779_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X15088 a_27215_13879# a_27311_13879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15089 vssd1 _0330_ a_16907_1985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X15090 vccd1 net45 a_19255_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15091 a_6519_21495# _0429_ a_6847_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15092 _0557_ _0556_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=2.1 w=0.65 l=0.15
X15093 vssd1 _0231_ a_23395_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15094 a_2493_15823# a_1959_15829# a_2398_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15095 vssd1 ctr\[8\] a_5661_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15097 a_20039_18695# _0459_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15098 temp1.capload\[13\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15099 a_24262_10383# _0476_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X15101 a_19609_28335# _0089_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15102 a_14085_26703# a_13551_26709# a_13990_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15104 _0085_ a_22291_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X15105 vccd1 a_22983_15431# _0537_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X15106 cal_lut\[97\] a_13203_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15107 a_18645_12043# _0440_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X15108 a_15765_23983# cal_lut\[45\] a_15693_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15109 vccd1 net24 a_6099_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15110 a_11025_10955# _0495_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X15112 vssd1 a_24835_19605# a_24842_19905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15113 a_3869_11989# clknet_0_net67 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15114 vccd1 _0408_ a_6745_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15115 cal_lut\[35\] a_16055_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15116 vssd1 net15 a_12895_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0894 ps=0.925 w=0.65 l=0.15
X15117 vccd1 _0323_ a_2971_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15118 temp1.capload\[11\].cap.Y clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15119 a_6814_12559# a_6541_12565# a_6729_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15120 a_16761_26703# _0690_ a_16679_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15121 vccd1 a_25011_14709# _0244_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X15122 a_18325_19453# _0453_ a_18243_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15123 vssd1 a_22438_8181# a_22396_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X15124 a_17249_29789# a_16911_29575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X15126 a_11799_3133# cal_lut\[147\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X15127 a_8251_9117# a_7553_8751# a_7994_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15128 a_5418_9269# a_5250_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15129 a_4115_28918# a_3933_28918# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15130 cal_lut\[119\] a_14307_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15131 _0324_ a_5359_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X15132 _0774_ a_7939_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X15133 vccd1 a_9000_19783# _0704_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X15134 a_13373_7485# cal_lut\[148\] a_13301_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15135 a_12517_7497# a_11527_7125# a_12391_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15136 vssd1 _0591_ _0785_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15137 vccd1 _0330_ a_19255_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X15138 vssd1 a_22843_9295# _0451_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X15139 vccd1 _0414_ a_3171_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15140 vssd1 a_12127_21959# _0709_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X15141 vssd1 _0447_ a_12950_16988# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X15142 a_17095_5639# _0445_ a_17329_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X15145 a_2139_12265# _0389_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15146 a_17727_17999# a_17029_18005# a_17470_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15147 vccd1 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ temp1.capload\[5\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15148 _0715_ a_9167_21601# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X15149 vccd1 _0261_ a_18979_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15150 a_5142_7775# a_4974_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15151 a_15469_26935# cal_lut\[91\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X15152 a_10229_23983# _0682_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X15153 a_27203_22173# a_26339_21807# a_26946_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15154 a_3575_15797# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.143 ps=1.33 w=0.42 l=0.15
X15155 vccd1 a_9447_8207# a_9615_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15156 a_8378_15823# a_7939_15829# a_8293_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15157 vssd1 a_2060_30199# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X15158 vccd1 _0517_ a_9423_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15159 a_24573_8751# a_24407_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15160 a_25235_22351# _0237_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X15161 _0557_ net16 a_12737_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X15162 a_3785_17999# _0422_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15163 a_24823_15444# _0244_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X15164 vssd1 a_2778_24527# clknet_0_temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15165 vssd1 _0420_ _0423_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X15166 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15167 _0655_ a_12162_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X15168 a_4068_31599# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X15169 vssd1 _0865_ a_15575_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15170 a_19609_4399# _0117_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X15171 vccd1 a_13146_23007# a_13073_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15172 cal_lut\[158\] a_22219_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15173 a_16911_29575# a_17007_29397# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X15174 vccd1 a_15725_15797# _0543_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X15175 _0083_ a_18979_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X15176 a_11884_21807# _0631_ a_11581_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X15177 a_20779_15253# _0850_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X15178 a_12518_1679# a_12079_1685# a_12433_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15179 a_3606_10660# a_3406_10505# a_3755_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X15180 a_20069_7663# _0110_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15181 vccd1 net35 a_20727_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15183 _0050_ a_14747_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15184 vccd1 a_6182_22895# clknet_1_1__leaf_io_in[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15185 a_1917_19881# _0418_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15186 a_23055_13469# a_22273_13103# a_22971_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15188 a_19465_17455# _0508_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X15189 a_18142_28068# a_17942_27913# a_18291_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X15192 a_6555_8207# a_6375_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15193 a_13990_26703# a_13551_26709# a_13905_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15194 a_20132_19394# dbg_result[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X15195 vssd1 a_25271_24349# a_25439_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15196 vccd1 io_in[0] a_6458_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15197 a_12269_18319# _0588_ a_11950_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X15198 clknet_0__0380_ a_7102_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15199 vssd1 a_6458_20175# clknet_0_io_in[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15200 vccd1 a_2071_11791# _0391_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X15201 a_10402_3677# a_10129_3311# a_10317_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15202 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15203 cal_lut\[150\] a_17895_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15204 vccd1 _0882_ a_9411_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15206 clknet_1_1__leaf_net67 a_3685_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15207 a_21166_2589# a_20727_2223# a_21081_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15209 vccd1 a_3848_27399# _0830_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X15212 vccd1 ctr\[2\] a_2695_14013# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.0588 ps=0.7 w=0.42 l=0.15
X15213 vccd1 a_1477_10901# clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15214 vssd1 _0657_ a_23361_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X15215 a_2153_11791# _0389_ a_2071_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X15216 a_16857_27023# cal_lut\[91\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X15217 vccd1 a_19827_25589# a_19743_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15218 a_2959_25071# _0803_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15219 vccd1 net49 temp1.capload\[0\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15220 a_9316_10927# _0451_ a_9126_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X15221 a_5911_22057# _0432_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15222 a_9071_14735# a_8289_14741# a_8987_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15223 vccd1 _0481_ a_9963_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X15224 vssd1 _0417_ a_2327_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15225 vssd1 _0364_ a_16955_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15226 a_6892_30083# ctr\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X15227 a_6823_17999# a_6375_18005# a_6729_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15228 _0345_ a_24771_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X15229 a_9253_21601# _0677_ a_9167_21601# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X15231 a_17930_25183# a_17762_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15233 a_24137_18543# cal_lut\[27\] a_24065_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15234 vccd1 _0160_ a_25941_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X15235 a_6516_20871# a_6646_21041# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X15237 a_9390_1501# a_8951_1135# a_9305_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15238 vssd1 a_12099_15547# a_12057_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15239 a_6817_3677# a_6283_3311# a_6722_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15240 vccd1 clknet_0_net67 a_3869_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15241 vccd1 a_7410_14709# dbg_result[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15242 a_22530_14709# a_22362_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15243 vccd1 cal_lut\[185\] a_16859_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15244 a_4032_25847# _0828_ a_4174_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X15245 vccd1 a_11214_5599# a_11141_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15247 a_4129_23439# _0790_ a_3695_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
X15248 vssd1 a_25842_17567# a_25800_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X15249 vccd1 _0784_ a_3933_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X15250 a_17677_1679# _0185_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15251 cal_lut\[103\] a_20287_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15252 vccd1 a_2778_24527# clknet_0_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15253 vccd1 _0476_ a_8675_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X15254 a_10779_28701# a_10331_28335# a_10685_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15255 a_17456_16617# _0246_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15256 vssd1 a_15725_15797# _0543_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X15257 vssd1 a_7718_14303# a_7676_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X15258 cal_lut\[100\] a_13847_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15259 a_12623_29967# net13 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X15260 a_10294_13215# a_10126_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15261 vccd1 net41 a_14931_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15262 cal_lut\[132\] a_14675_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15263 vssd1 _0443_ a_21029_6369# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X15264 vssd1 a_10294_11445# a_10252_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X15265 a_21675_2589# a_20893_2223# a_21591_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15266 vssd1 a_3869_11989# clknet_1_0__leaf_net67 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X15267 vssd1 a_18355_1653# a_18313_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15268 vssd1 _0456_ a_22740_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X15269 a_2014_12533# a_1846_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15270 a_24377_20553# a_23823_20393# a_24030_20452# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X15271 a_22322_4649# _0283_ a_22240_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15272 a_7691_2589# a_6909_2223# a_7607_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15273 vccd1 a_27583_9514# _0170_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15275 vccd1 _0476_ a_4531_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X15276 a_22362_14735# a_22089_14741# a_22277_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15277 cal_lut\[156\] a_18723_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15278 a_15795_28879# a_15097_28885# a_15538_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15279 a_20157_16917# a_19991_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15280 a_4605_12937# a_3615_12565# a_4479_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15281 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_1407_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X15282 a_17831_16189# a_17611_16201# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X15283 vccd1 a_1753_26133# clknet_1_1__leaf_temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15284 vccd1 a_2566_15797# a_2493_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15285 a_5996_21807# ctr\[9\] a_5693_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X15286 vssd1 _0475_ a_18140_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X15287 a_14153_20884# _0485_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X15288 vccd1 a_14158_26677# a_14085_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15289 vssd1 a_14103_17455# _0447_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15292 vssd1 a_13459_4399# _0283_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X15293 a_20004_27081# a_19605_26709# a_19878_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15294 vccd1 a_21759_4667# a_21675_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15295 vccd1 _0835_ a_6835_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15296 vssd1 cal_lut\[1\] a_6737_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15297 vccd1 a_22711_6549# _0343_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X15298 a_20676_9001# _0283_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15300 a_25823_23439# a_25125_23445# a_25566_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15301 a_22013_17027# _0684_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X15302 a_2605_21263# _0772_ a_2511_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X15303 vssd1 _0720_ a_10883_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0878 ps=0.92 w=0.65 l=0.15
X15306 a_24459_8181# cal_lut\[164\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X15307 a_6020_10927# a_5621_10927# a_5894_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15308 a_9678_24233# _0712_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X15309 _0260_ a_13367_10391# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X15310 vccd1 a_23903_18695# _0642_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X15311 dbg_result[3] a_7410_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X15312 a_15186_13647# a_14747_13653# a_15101_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15313 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd net11 a_9049_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X15314 a_6437_27247# a_5883_27221# a_6090_27221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X15315 vccd1 net35 a_18335_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15317 vssd1 a_12851_2589# a_13019_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15318 a_22247_9991# _0452_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X15319 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15320 _0787_ ctr\[6\] a_5630_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X15322 vccd1 _0450_ a_21831_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15323 io_out[0] a_2023_19319# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15324 a_9221_2223# a_8951_2589# a_9131_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X15325 vccd1 _0863_ a_11527_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X15326 vssd1 a_15519_27791# a_15687_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15327 vccd1 a_4789_11703# net75 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X15328 _0813_ a_5487_29217# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X15330 a_15427_21263# a_14563_21269# a_15170_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15332 clknet_0_temp1.i_precharge_n a_2778_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15333 _0254_ a_17456_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X15334 a_5825_15823# _0839_ _0192_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15335 vssd1 _0339_ a_17415_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15336 vccd1 _0330_ a_13459_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X15337 a_5341_17429# clknet_0_io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15338 a_22005_21629# _0531_ a_21923_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15339 _0866_ a_18192_15529# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X15340 a_16807_11293# a_15943_10927# a_16550_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X15341 vccd1 _0227_ a_19531_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15342 vccd1 ctr\[3\] a_2887_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15343 a_2921_17999# _0420_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X15344 a_12163_30287# net14 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X15346 vccd1 net11 a_9319_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X15348 a_19878_28879# a_19605_28885# a_19793_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15349 a_3066_27569# a_3017_27399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X15350 vccd1 a_11030_27383# a_10964_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X15351 a_5073_14735# _0205_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X15352 a_19694_15645# a_19421_15279# a_19609_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X15353 vccd1 _0498_ a_16220_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X15354 vccd1 _0341_ a_26339_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X15355 a_15097_21263# a_14563_21269# a_15002_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15356 vssd1 a_7607_2589# a_7775_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15357 _0403_ net73 a_7381_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15359 a_11847_3073# _0330_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X15360 _0848_ a_12995_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X15361 vccd1 a_17107_4073# a_17114_3977# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15362 a_6522_29535# a_6354_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15363 vssd1 clknet_1_1__leaf_io_in[0] a_10423_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15364 vssd1 a_8419_11195# a_8377_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15365 a_4040_11587# ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X15366 a_2010_24759# _0410_ a_2330_24887# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X15367 a_8390_23439# clknet_0__0380_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15368 a_21090_26159# a_20775_26311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X15369 a_16477_11293# a_15943_10927# a_16382_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15370 vssd1 a_3117_12533# _0203_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X15371 a_23754_26980# a_23547_26921# a_23930_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X15372 a_4997_23805# ctr\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15373 vccd1 _0425_ a_8397_20983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X15374 a_8532_31751# net11 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X15375 vssd1 a_6779_29789# a_6947_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15376 vccd1 _0410_ _0804_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15377 vccd1 a_2747_18517# net22 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X15378 _0641_ a_22659_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X15379 vssd1 a_13997_28023# _0271_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X15380 vssd1 _0421_ _0429_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15381 vssd1 a_10843_2197# _0373_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X15382 clknet_1_1__leaf__0380_ a_8390_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X15383 a_8853_21583# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15384 a_5460_17999# net72 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15385 a_3965_9839# a_3799_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15386 _0425_ a_7631_17171# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
R35 vssd1 net49 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X15388 vccd1 a_17286_9269# a_17213_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15389 a_25313_23439# _0062_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15390 a_2221_13255# _0411_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X15391 a_12644_2057# a_12245_1685# a_12518_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15392 vccd1 a_20839_22325# a_20755_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15393 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd _0419_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15394 _0434_ _0421_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15395 vccd1 net26 a_9963_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15396 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_3891_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X15397 a_25769_17821# a_25235_17455# a_25674_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15398 cal_lut\[118\] a_20287_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15399 vccd1 a_4811_30511# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X15400 net9 a_9687_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X15401 a_13040_6147# _0299_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15402 a_5573_29217# ctr\[9\] a_5487_29217# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X15403 a_15370_19407# a_15115_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.312 ps=2.12 w=1 l=0.15
X15404 vssd1 _0486_ a_15093_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X15406 a_21983_4943# cal_lut\[151\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X15408 vccd1 a_5841_19605# a_5871_19958# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15409 a_16187_23671# _0464_ a_16361_23777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X15410 vccd1 a_27491_17130# _0073_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15411 a_17489_1685# a_17323_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15412 _0489_ a_15391_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X15413 a_21292_2223# a_20893_2223# a_21166_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15414 a_23119_24349# _0216_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X15415 a_11141_5853# a_10607_5487# a_11046_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X15416 a_5675_9295# a_4977_9301# a_5418_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15417 a_13213_16911# _0438_ a_13129_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X15418 vccd1 a_18107_8439# _0607_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X15419 vccd1 cal_lut\[51\] a_16859_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15420 vssd1 ctr\[7\] a_5864_26819# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15421 a_15943_7232# cal_lut\[138\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X15422 vssd1 a_11857_18517# _0628_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X15423 a_7476_21583# _0437_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X15424 a_23273_27247# a_22726_27521# a_22926_27221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X15425 clknet_1_1__leaf_temp1.i_precharge_n a_1753_26133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15427 a_7011_31599# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X15428 vccd1 a_13111_1653# a_13027_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15429 a_17493_6575# _0112_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15430 a_2099_18695# _0420_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X15431 a_24761_7119# _0163_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15432 a_23757_10927# _0506_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X15433 a_7716_22325# _0755_ a_8108_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X15434 a_17661_4233# a_17114_3977# a_17314_4132# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X15435 vccd1 a_12672_30199# a_12623_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X15437 vssd1 _0771_ a_2797_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15438 _0433_ a_8544_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X15440 a_9516_1135# a_9117_1135# a_9390_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15441 a_5404_9001# _0838_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15442 a_19881_9301# a_19715_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15443 a_11877_26709# a_11711_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15444 a_26394_6687# a_26226_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15445 vccd1 a_6779_9117# a_6947_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15446 a_23792_10089# _0656_ a_23690_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X15447 a_21034_10499# _0283_ a_20952_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X15448 a_17075_22173# a_16293_21807# a_16991_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15449 vssd1 a_22695_1679# a_22863_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15450 a_15078_7093# a_14910_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X15451 a_8377_16367# a_7387_16367# a_8251_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15452 _0714_ _0711_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15453 vssd1 a_18751_23671# _0620_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X15454 vssd1 _0347_ a_26799_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15455 vssd1 a_5567_7931# a_5525_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15456 vccd1 a_8348_32375# a_8299_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X15457 vccd1 clknet_0_net67 a_3685_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15458 a_4747_10205# a_3965_9839# a_4663_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15459 a_15009_27791# _0091_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X15460 a_10964_27613# a_10423_27247# a_10871_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X15461 vssd1 _0864_ a_11987_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X15462 a_26394_6687# a_26226_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15463 a_23759_16733# a_23579_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15464 vccd1 a_3869_11989# clknet_1_0__leaf_net67 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15466 vssd1 _0438_ _0485_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15468 vccd1 net10 a_8123_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X15469 vssd1 a_17930_25183# a_17888_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X15471 _0859_ a_17088_12265# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X15475 vccd1 a_8143_14459# a_8059_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15476 vccd1 a_1937_6549# clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15477 a_12349_9661# a_12079_9295# a_12259_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X15478 a_24919_10901# a_25210_11201# a_25161_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X15479 vccd1 a_24835_13077# a_24842_13377# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X15480 vssd1 _0429_ a_4339_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X15482 a_20046_28853# a_19878_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X15483 vccd1 _0794_ a_5645_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15484 vssd1 _0721_ a_8268_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X15486 vssd1 _0767_ a_7665_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X15487 vssd1 a_9613_20693# a_9547_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X15488 _0443_ a_19915_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.331 ps=1.71 w=1 l=0.15
X15489 vccd1 a_17470_17973# a_17397_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X15490 vssd1 a_19367_13621# a_19325_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15491 a_4698_5853# a_4259_5487# a_4613_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15492 vssd1 a_5143_11445# a_4885_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X15493 vccd1 _0877_ a_25235_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X15494 _0193_ ctr\[3\] a_4733_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15495 vssd1 net26 a_14471_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 io_in[1] vssd1 1.17f
C1 dbg_delay vssd1 13.6f
C2 io_in[2] vssd1 1.1f
C3 io_in[3] vssd1 1.19f
C4 io_in[4] vssd1 1.33f
C5 io_in[5] vssd1 1.17f
C6 io_in[6] vssd1 1.1f
C7 io_in[7] vssd1 1.23f
C8 dbg_result[0] vssd1 17.1f
C9 dbg_result[1] vssd1 21f
C10 dbg_result[2] vssd1 16.9f
C11 io_out[0] vssd1 2.69f
C12 io_out[1] vssd1 1.41f
C13 io_in[0] vssd1 10.8f
C14 dbg_result[3] vssd1 19.6f
C15 io_out[2] vssd1 1.86f
C16 io_out[3] vssd1 2.22f
C17 io_out[4] vssd1 1.67f
C18 io_out[5] vssd1 2.78f
C19 dbg_result[4] vssd1 18f
C20 dbg_result[5] vssd1 19f
C21 io_out[6] vssd1 1.27f
C22 io_out[7] vssd1 1.32f
C23 vccd1 vssd1 3.42p
C24 a_14457_1135# vssd1 0.23f $ **FLOATING
C25 a_22059_1109# vssd1 0.604f $ **FLOATING
C26 a_21883_1109# vssd1 0.508f $ **FLOATING
C27 a_19439_1135# vssd1 0.524f $ **FLOATING
C28 a_17231_1135# vssd1 0.524f $ **FLOATING
C29 _0372_ vssd1 0.675f $ **FLOATING
C30 a_16859_1501# vssd1 0.508f $ **FLOATING
C31 a_16679_1501# vssd1 0.604f $ **FLOATING
C32 a_14967_1501# vssd1 0.609f $ **FLOATING
C33 a_15135_1403# vssd1 0.817f $ **FLOATING
C34 a_14542_1501# vssd1 0.626f $ **FLOATING
C35 a_14710_1247# vssd1 0.581f $ **FLOATING
C36 a_14269_1135# vssd1 1.43f $ **FLOATING
C37 a_14103_1135# vssd1 1.81f $ **FLOATING
C38 a_9305_1135# vssd1 0.23f $ **FLOATING
C39 a_11987_1135# vssd1 0.524f $ **FLOATING
C40 a_9815_1501# vssd1 0.609f $ **FLOATING
C41 a_9983_1403# vssd1 0.817f $ **FLOATING
C42 a_9390_1501# vssd1 0.626f $ **FLOATING
C43 a_9558_1247# vssd1 0.581f $ **FLOATING
C44 a_9117_1135# vssd1 1.43f $ **FLOATING
C45 a_8951_1135# vssd1 1.81f $ **FLOATING
C46 a_22185_1679# vssd1 0.23f $ **FLOATING
C47 a_20253_1679# vssd1 0.23f $ **FLOATING
C48 _0334_ vssd1 0.922f $ **FLOATING
C49 a_17677_1679# vssd1 0.23f $ **FLOATING
C50 a_15101_1679# vssd1 0.23f $ **FLOATING
C51 a_12433_1679# vssd1 0.23f $ **FLOATING
C52 _0370_ vssd1 0.837f $ **FLOATING
C53 a_10317_1679# vssd1 0.23f $ **FLOATING
C54 a_8293_1679# vssd1 0.23f $ **FLOATING
C55 a_22695_1679# vssd1 0.609f $ **FLOATING
C56 a_22863_1653# vssd1 0.817f $ **FLOATING
C57 a_22270_1679# vssd1 0.626f $ **FLOATING
C58 a_22438_1653# vssd1 0.581f $ **FLOATING
C59 a_21997_1685# vssd1 1.43f $ **FLOATING
C60 _0151_ vssd1 0.911f $ **FLOATING
C61 a_21831_1685# vssd1 1.81f $ **FLOATING
C62 a_21463_1679# vssd1 0.524f $ **FLOATING
C63 _0335_ vssd1 1f $ **FLOATING
C64 a_20763_1679# vssd1 0.609f $ **FLOATING
C65 a_20931_1653# vssd1 0.817f $ **FLOATING
C66 a_20338_1679# vssd1 0.626f $ **FLOATING
C67 a_20506_1653# vssd1 0.581f $ **FLOATING
C68 a_20065_1685# vssd1 1.43f $ **FLOATING
C69 _0150_ vssd1 1.19f $ **FLOATING
C70 a_19899_1685# vssd1 1.81f $ **FLOATING
C71 a_19439_1679# vssd1 0.524f $ **FLOATING
C72 a_18975_1679# vssd1 0.508f $ **FLOATING
C73 a_18795_1679# vssd1 0.604f $ **FLOATING
C74 a_18187_1679# vssd1 0.609f $ **FLOATING
C75 a_18355_1653# vssd1 0.817f $ **FLOATING
C76 a_17762_1679# vssd1 0.626f $ **FLOATING
C77 a_17930_1653# vssd1 0.581f $ **FLOATING
C78 a_17489_1685# vssd1 1.43f $ **FLOATING
C79 _0185_ vssd1 1.03f $ **FLOATING
C80 a_17323_1685# vssd1 1.81f $ **FLOATING
C81 a_16907_1985# vssd1 0.604f $ **FLOATING
C82 a_16731_1653# vssd1 0.508f $ **FLOATING
C83 a_16311_1679# vssd1 0.524f $ **FLOATING
C84 _0333_ vssd1 0.761f $ **FLOATING
C85 a_15611_1679# vssd1 0.609f $ **FLOATING
C86 a_15779_1653# vssd1 0.817f $ **FLOATING
C87 a_15186_1679# vssd1 0.626f $ **FLOATING
C88 a_15354_1653# vssd1 0.581f $ **FLOATING
C89 a_14913_1685# vssd1 1.43f $ **FLOATING
C90 _0184_ vssd1 0.911f $ **FLOATING
C91 a_14747_1685# vssd1 1.81f $ **FLOATING
C92 a_14379_1679# vssd1 0.524f $ **FLOATING
C93 _0371_ vssd1 0.725f $ **FLOATING
C94 a_13823_1679# vssd1 0.508f $ **FLOATING
C95 a_13643_1679# vssd1 0.604f $ **FLOATING
C96 a_12943_1679# vssd1 0.609f $ **FLOATING
C97 a_13111_1653# vssd1 0.817f $ **FLOATING
C98 a_12518_1679# vssd1 0.626f $ **FLOATING
C99 a_12686_1653# vssd1 0.581f $ **FLOATING
C100 a_12245_1685# vssd1 1.43f $ **FLOATING
C101 _0183_ vssd1 1.03f $ **FLOATING
C102 a_12079_1685# vssd1 1.81f $ **FLOATING
C103 a_11707_1679# vssd1 0.508f $ **FLOATING
C104 a_11527_1679# vssd1 0.604f $ **FLOATING
C105 a_10827_1679# vssd1 0.609f $ **FLOATING
C106 a_10995_1653# vssd1 0.817f $ **FLOATING
C107 a_10402_1679# vssd1 0.626f $ **FLOATING
C108 a_10570_1653# vssd1 0.581f $ **FLOATING
C109 a_10129_1685# vssd1 1.43f $ **FLOATING
C110 a_9963_1685# vssd1 1.81f $ **FLOATING
C111 a_9591_1679# vssd1 0.508f $ **FLOATING
C112 a_9411_1679# vssd1 0.604f $ **FLOATING
C113 a_8803_1679# vssd1 0.609f $ **FLOATING
C114 a_8971_1653# vssd1 0.817f $ **FLOATING
C115 a_8378_1679# vssd1 0.626f $ **FLOATING
C116 a_8546_1653# vssd1 0.581f $ **FLOATING
C117 a_8105_1685# vssd1 1.43f $ **FLOATING
C118 a_7939_1685# vssd1 1.81f $ **FLOATING
C119 a_7251_1898# vssd1 0.524f $ **FLOATING
C120 a_21081_2223# vssd1 0.23f $ **FLOATING
C121 a_22471_2589# vssd1 0.508f $ **FLOATING
C122 a_22291_2589# vssd1 0.604f $ **FLOATING
C123 a_21591_2589# vssd1 0.609f $ **FLOATING
C124 a_21759_2491# vssd1 0.817f $ **FLOATING
C125 a_21166_2589# vssd1 0.626f $ **FLOATING
C126 a_21334_2335# vssd1 0.581f $ **FLOATING
C127 a_20893_2223# vssd1 1.43f $ **FLOATING
C128 a_20727_2223# vssd1 1.81f $ **FLOATING
C129 a_20237_2223# vssd1 0.23f $ **FLOATING
C130 a_17217_2223# vssd1 0.23f $ **FLOATING
C131 _0154_ vssd1 1.23f $ **FLOATING
C132 a_19819_2223# vssd1 0.581f $ **FLOATING
C133 a_19890_2197# vssd1 0.626f $ **FLOATING
C134 a_19683_2197# vssd1 1.81f $ **FLOATING
C135 a_19690_2497# vssd1 1.43f $ **FLOATING
C136 a_19399_2197# vssd1 0.609f $ **FLOATING
C137 a_19303_2375# vssd1 0.817f $ **FLOATING
C138 a_17727_2589# vssd1 0.609f $ **FLOATING
C139 a_17895_2491# vssd1 0.817f $ **FLOATING
C140 a_17302_2589# vssd1 0.626f $ **FLOATING
C141 a_17470_2335# vssd1 0.581f $ **FLOATING
C142 a_17029_2223# vssd1 1.43f $ **FLOATING
C143 _0149_ vssd1 1.17f $ **FLOATING
C144 a_16863_2223# vssd1 1.81f $ **FLOATING
C145 _0148_ vssd1 1.23f $ **FLOATING
C146 a_12341_2223# vssd1 0.23f $ **FLOATING
C147 a_15439_2388# vssd1 0.524f $ **FLOATING
C148 a_14103_2223# vssd1 0.524f $ **FLOATING
C149 _0332_ vssd1 0.686f $ **FLOATING
C150 a_13639_2589# vssd1 0.508f $ **FLOATING
C151 a_13459_2589# vssd1 0.604f $ **FLOATING
C152 a_12851_2589# vssd1 0.609f $ **FLOATING
C153 a_13019_2491# vssd1 0.817f $ **FLOATING
C154 a_12426_2589# vssd1 0.626f $ **FLOATING
C155 a_12594_2335# vssd1 0.581f $ **FLOATING
C156 a_12153_2223# vssd1 1.43f $ **FLOATING
C157 a_11987_2223# vssd1 1.81f $ **FLOATING
C158 _0147_ vssd1 0.872f $ **FLOATING
C159 _0373_ vssd1 2.33f $ **FLOATING
C160 _0182_ vssd1 0.922f $ **FLOATING
C161 _0181_ vssd1 1.3f $ **FLOATING
C162 a_7097_2223# vssd1 0.23f $ **FLOATING
C163 a_11711_2223# vssd1 0.524f $ **FLOATING
C164 a_11019_2197# vssd1 0.604f $ **FLOATING
C165 a_10843_2197# vssd1 0.508f $ **FLOATING
C166 a_10055_2223# vssd1 0.524f $ **FLOATING
C167 _0369_ vssd1 0.895f $ **FLOATING
C168 _0368_ vssd1 0.725f $ **FLOATING
C169 a_9551_2388# vssd1 0.524f $ **FLOATING
C170 a_9131_2589# vssd1 0.508f $ **FLOATING
C171 a_8951_2589# vssd1 0.604f $ **FLOATING
C172 a_7607_2589# vssd1 0.609f $ **FLOATING
C173 a_7775_2491# vssd1 0.817f $ **FLOATING
C174 a_7182_2589# vssd1 0.626f $ **FLOATING
C175 a_7350_2335# vssd1 0.581f $ **FLOATING
C176 a_6909_2223# vssd1 1.43f $ **FLOATING
C177 _0186_ vssd1 0.994f $ **FLOATING
C178 a_6743_2223# vssd1 1.81f $ **FLOATING
C179 a_23457_3145# vssd1 0.23f $ **FLOATING
C180 _0153_ vssd1 1.03f $ **FLOATING
C181 _0338_ vssd1 1.08f $ **FLOATING
C182 a_15193_2767# vssd1 0.23f $ **FLOATING
C183 _0331_ vssd1 0.957f $ **FLOATING
C184 _0180_ vssd1 1.25f $ **FLOATING
C185 a_23039_3145# vssd1 0.581f $ **FLOATING
C186 a_23110_3044# vssd1 0.626f $ **FLOATING
C187 a_22910_2889# vssd1 1.43f $ **FLOATING
C188 a_22903_2985# vssd1 1.81f $ **FLOATING
C189 a_22619_2999# vssd1 0.609f $ **FLOATING
C190 a_22523_2999# vssd1 0.817f $ **FLOATING
C191 a_22151_3073# vssd1 0.604f $ **FLOATING
C192 a_21975_2741# vssd1 0.508f $ **FLOATING
C193 _0337_ vssd1 0.998f $ **FLOATING
C194 a_20867_2986# vssd1 0.524f $ **FLOATING
C195 a_19759_3073# vssd1 0.604f $ **FLOATING
C196 a_19583_2741# vssd1 0.508f $ **FLOATING
C197 a_17919_3073# vssd1 0.604f $ **FLOATING
C198 a_17743_2741# vssd1 0.508f $ **FLOATING
C199 a_15703_2767# vssd1 0.609f $ **FLOATING
C200 a_15871_2741# vssd1 0.817f $ **FLOATING
C201 a_15278_2767# vssd1 0.626f $ **FLOATING
C202 a_15446_2741# vssd1 0.581f $ **FLOATING
C203 a_15005_2773# vssd1 1.43f $ **FLOATING
C204 _0179_ vssd1 1.09f $ **FLOATING
C205 a_14839_2773# vssd1 1.81f $ **FLOATING
C206 a_12223_2741# vssd1 0.698f $ **FLOATING
C207 a_11847_3073# vssd1 0.604f $ **FLOATING
C208 a_11671_2741# vssd1 0.508f $ **FLOATING
C209 a_9963_2767# vssd1 0.524f $ **FLOATING
C210 a_9547_3073# vssd1 0.604f $ **FLOATING
C211 a_9371_2741# vssd1 0.508f $ **FLOATING
C212 _0367_ vssd1 0.881f $ **FLOATING
C213 a_8539_2986# vssd1 0.524f $ **FLOATING
C214 _0152_ vssd1 1.23f $ **FLOATING
C215 a_20437_3311# vssd1 0.23f $ **FLOATING
C216 a_23671_3311# vssd1 0.524f $ **FLOATING
C217 a_22659_3311# vssd1 0.524f $ **FLOATING
C218 _0336_ vssd1 1.07f $ **FLOATING
C219 a_20947_3677# vssd1 0.609f $ **FLOATING
C220 a_21115_3579# vssd1 0.817f $ **FLOATING
C221 a_20522_3677# vssd1 0.626f $ **FLOATING
C222 a_20690_3423# vssd1 0.581f $ **FLOATING
C223 a_20249_3311# vssd1 1.43f $ **FLOATING
C224 a_20083_3311# vssd1 1.81f $ **FLOATING
C225 _0156_ vssd1 0.872f $ **FLOATING
C226 a_18045_3311# vssd1 0.23f $ **FLOATING
C227 a_19807_3311# vssd1 0.524f $ **FLOATING
C228 _0340_ vssd1 0.647f $ **FLOATING
C229 a_19435_3677# vssd1 0.508f $ **FLOATING
C230 a_19255_3677# vssd1 0.604f $ **FLOATING
C231 _0330_ vssd1 11.6f $ **FLOATING
C232 a_18555_3677# vssd1 0.609f $ **FLOATING
C233 a_18723_3579# vssd1 0.817f $ **FLOATING
C234 a_18130_3677# vssd1 0.626f $ **FLOATING
C235 a_18298_3423# vssd1 0.581f $ **FLOATING
C236 a_17857_3311# vssd1 1.43f $ **FLOATING
C237 a_17691_3311# vssd1 1.81f $ **FLOATING
C238 _0155_ vssd1 0.872f $ **FLOATING
C239 _0366_ vssd1 1.17f $ **FLOATING
C240 a_11789_3311# vssd1 0.23f $ **FLOATING
C241 a_17415_3311# vssd1 0.524f $ **FLOATING
C242 _0339_ vssd1 0.934f $ **FLOATING
C243 a_16859_3677# vssd1 0.508f $ **FLOATING
C244 a_16679_3677# vssd1 0.604f $ **FLOATING
C245 a_16079_3285# vssd1 0.604f $ **FLOATING
C246 a_15903_3285# vssd1 0.508f $ **FLOATING
C247 a_15479_3677# vssd1 0.508f $ **FLOATING
C248 a_15299_3677# vssd1 0.604f $ **FLOATING
C249 a_14331_3285# vssd1 0.604f $ **FLOATING
C250 a_14155_3285# vssd1 0.508f $ **FLOATING
C251 a_12955_3476# vssd1 0.524f $ **FLOATING
C252 a_12299_3677# vssd1 0.609f $ **FLOATING
C253 a_12467_3579# vssd1 0.817f $ **FLOATING
C254 a_11874_3677# vssd1 0.626f $ **FLOATING
C255 a_12042_3423# vssd1 0.581f $ **FLOATING
C256 a_11601_3311# vssd1 1.43f $ **FLOATING
C257 a_11435_3311# vssd1 1.81f $ **FLOATING
C258 a_10317_3311# vssd1 0.23f $ **FLOATING
C259 a_10827_3677# vssd1 0.609f $ **FLOATING
C260 a_10995_3579# vssd1 0.817f $ **FLOATING
C261 a_10402_3677# vssd1 0.626f $ **FLOATING
C262 a_10570_3423# vssd1 0.581f $ **FLOATING
C263 a_10129_3311# vssd1 1.43f $ **FLOATING
C264 _0146_ vssd1 0.954f $ **FLOATING
C265 a_9963_3311# vssd1 1.81f $ **FLOATING
C266 a_6637_3311# vssd1 0.23f $ **FLOATING
C267 a_9595_3311# vssd1 0.698f $ **FLOATING
C268 a_8171_3476# vssd1 0.524f $ **FLOATING
C269 a_7147_3677# vssd1 0.609f $ **FLOATING
C270 a_7315_3579# vssd1 0.817f $ **FLOATING
C271 a_6722_3677# vssd1 0.626f $ **FLOATING
C272 a_6890_3423# vssd1 0.581f $ **FLOATING
C273 a_6449_3311# vssd1 1.43f $ **FLOATING
C274 a_6283_3311# vssd1 1.81f $ **FLOATING
C275 a_5451_3677# vssd1 0.508f $ **FLOATING
C276 a_5271_3677# vssd1 0.604f $ **FLOATING
C277 a_24653_4233# vssd1 0.23f $ **FLOATING
C278 a_22553_3855# vssd1 0.23f $ **FLOATING
C279 a_17661_4233# vssd1 0.23f $ **FLOATING
C280 a_15469_3855# vssd1 0.23f $ **FLOATING
C281 a_13997_3855# vssd1 0.23f $ **FLOATING
C282 a_12525_3855# vssd1 0.23f $ **FLOATING
C283 _0363_ vssd1 11.4f $ **FLOATING
C284 _0314_ vssd1 1.83f $ **FLOATING
C285 _0329_ vssd1 1.19f $ **FLOATING
C286 a_9358_3855# vssd1 0.333f $ **FLOATING
C287 a_8017_3855# vssd1 0.23f $ **FLOATING
C288 _0133_ vssd1 1.06f $ **FLOATING
C289 a_5165_3855# vssd1 0.23f $ **FLOATING
C290 _0116_ vssd1 1.36f $ **FLOATING
C291 a_24235_4233# vssd1 0.581f $ **FLOATING
C292 a_24306_4132# vssd1 0.626f $ **FLOATING
C293 a_24106_3977# vssd1 1.43f $ **FLOATING
C294 a_24099_4073# vssd1 1.81f $ **FLOATING
C295 a_23815_4087# vssd1 0.609f $ **FLOATING
C296 a_23719_4087# vssd1 0.817f $ **FLOATING
C297 a_23063_3855# vssd1 0.609f $ **FLOATING
C298 a_23231_3829# vssd1 0.817f $ **FLOATING
C299 a_22638_3855# vssd1 0.626f $ **FLOATING
C300 a_22806_3829# vssd1 0.581f $ **FLOATING
C301 a_22365_3861# vssd1 1.43f $ **FLOATING
C302 a_22199_3861# vssd1 1.81f $ **FLOATING
C303 a_20727_3855# vssd1 0.524f $ **FLOATING
C304 _0298_ vssd1 0.725f $ **FLOATING
C305 a_19763_4074# vssd1 0.524f $ **FLOATING
C306 a_19343_3855# vssd1 0.508f $ **FLOATING
C307 a_19163_3855# vssd1 0.604f $ **FLOATING
C308 a_17243_4233# vssd1 0.581f $ **FLOATING
C309 a_17314_4132# vssd1 0.626f $ **FLOATING
C310 a_17114_3977# vssd1 1.43f $ **FLOATING
C311 a_17107_4073# vssd1 1.81f $ **FLOATING
C312 a_16823_4087# vssd1 0.609f $ **FLOATING
C313 a_16727_4087# vssd1 0.817f $ **FLOATING
C314 a_15979_3855# vssd1 0.609f $ **FLOATING
C315 a_16147_3829# vssd1 0.817f $ **FLOATING
C316 a_15554_3855# vssd1 0.626f $ **FLOATING
C317 a_15722_3829# vssd1 0.581f $ **FLOATING
C318 a_15281_3861# vssd1 1.43f $ **FLOATING
C319 a_15115_3861# vssd1 1.81f $ **FLOATING
C320 a_14507_3855# vssd1 0.609f $ **FLOATING
C321 a_14675_3829# vssd1 0.817f $ **FLOATING
C322 a_14082_3855# vssd1 0.626f $ **FLOATING
C323 a_14250_3829# vssd1 0.581f $ **FLOATING
C324 a_13809_3861# vssd1 1.43f $ **FLOATING
C325 a_13643_3861# vssd1 1.81f $ **FLOATING
C326 a_13035_3855# vssd1 0.609f $ **FLOATING
C327 a_13203_3829# vssd1 0.817f $ **FLOATING
C328 a_12610_3855# vssd1 0.626f $ **FLOATING
C329 a_12778_3829# vssd1 0.581f $ **FLOATING
C330 a_12337_3861# vssd1 1.43f $ **FLOATING
C331 _0130_ vssd1 1.16f $ **FLOATING
C332 a_12171_3861# vssd1 1.81f $ **FLOATING
C333 net25 vssd1 10.3f $ **FLOATING
C334 a_11579_3829# vssd1 0.698f $ **FLOATING
C335 a_10835_4161# vssd1 0.604f $ **FLOATING
C336 a_10659_3829# vssd1 0.508f $ **FLOATING
C337 a_10051_3855# vssd1 0.508f $ **FLOATING
C338 a_9871_3855# vssd1 0.604f $ **FLOATING
C339 cal_lut\[181\] vssd1 2.41f $ **FLOATING
C340 a_9201_3829# vssd1 0.723f $ **FLOATING
C341 a_8527_3855# vssd1 0.609f $ **FLOATING
C342 a_8695_3829# vssd1 0.817f $ **FLOATING
C343 a_8102_3855# vssd1 0.626f $ **FLOATING
C344 a_8270_3829# vssd1 0.581f $ **FLOATING
C345 a_7829_3861# vssd1 1.43f $ **FLOATING
C346 _0132_ vssd1 1.05f $ **FLOATING
C347 a_7663_3861# vssd1 1.81f $ **FLOATING
C348 a_6791_4074# vssd1 0.524f $ **FLOATING
C349 a_5675_3855# vssd1 0.609f $ **FLOATING
C350 a_5843_3829# vssd1 0.817f $ **FLOATING
C351 a_5250_3855# vssd1 0.626f $ **FLOATING
C352 a_5418_3829# vssd1 0.581f $ **FLOATING
C353 a_4977_3861# vssd1 1.43f $ **FLOATING
C354 a_4811_3861# vssd1 1.81f $ **FLOATING
C355 _0115_ vssd1 1.49f $ **FLOATING
C356 _0297_ vssd1 1.11f $ **FLOATING
C357 cal_lut\[152\] vssd1 2.56f $ **FLOATING
C358 a_21081_4399# vssd1 0.23f $ **FLOATING
C359 _0296_ vssd1 1.31f $ **FLOATING
C360 a_23811_4564# vssd1 0.524f $ **FLOATING
C361 a_23344_4649# vssd1 0.502f $ **FLOATING
C362 a_22843_4399# vssd1 0.619f $ **FLOATING
C363 a_22240_4649# vssd1 0.502f $ **FLOATING
C364 a_21591_4765# vssd1 0.609f $ **FLOATING
C365 a_21759_4667# vssd1 0.817f $ **FLOATING
C366 a_21166_4765# vssd1 0.626f $ **FLOATING
C367 a_21334_4511# vssd1 0.581f $ **FLOATING
C368 a_20893_4399# vssd1 1.43f $ **FLOATING
C369 _0114_ vssd1 0.954f $ **FLOATING
C370 a_20727_4399# vssd1 1.81f $ **FLOATING
C371 a_19609_4399# vssd1 0.23f $ **FLOATING
C372 a_20119_4765# vssd1 0.609f $ **FLOATING
C373 a_20287_4667# vssd1 0.817f $ **FLOATING
C374 a_19694_4765# vssd1 0.626f $ **FLOATING
C375 a_19862_4511# vssd1 0.581f $ **FLOATING
C376 a_19421_4399# vssd1 1.43f $ **FLOATING
C377 _0117_ vssd1 0.994f $ **FLOATING
C378 a_19255_4399# vssd1 1.81f $ **FLOATING
C379 a_17875_4399# vssd1 0.648f $ **FLOATING
C380 _0177_ vssd1 1.31f $ **FLOATING
C381 a_16955_4399# vssd1 0.524f $ **FLOATING
C382 _0364_ vssd1 1.11f $ **FLOATING
C383 net31 vssd1 10.3f $ **FLOATING
C384 _0178_ vssd1 0.955f $ **FLOATING
C385 _0131_ vssd1 0.994f $ **FLOATING
C386 a_16640_4373# vssd1 0.648f $ **FLOATING
C387 _0365_ vssd1 1.07f $ **FLOATING
C388 a_15531_4564# vssd1 0.524f $ **FLOATING
C389 _0313_ vssd1 1.11f $ **FLOATING
C390 a_14151_4564# vssd1 0.524f $ **FLOATING
C391 a_13459_4399# vssd1 0.648f $ **FLOATING
C392 _0312_ vssd1 1.17f $ **FLOATING
C393 _0129_ vssd1 1.19f $ **FLOATING
C394 a_12535_4765# vssd1 0.508f $ **FLOATING
C395 a_12355_4765# vssd1 0.604f $ **FLOATING
C396 a_11759_4564# vssd1 0.524f $ **FLOATING
C397 a_10699_4399# vssd1 1.2f $ **FLOATING
C398 a_9542_4649# vssd1 0.333f $ **FLOATING
C399 cal_lut\[133\] vssd1 2.09f $ **FLOATING
C400 _0315_ vssd1 0.891f $ **FLOATING
C401 _0134_ vssd1 1.18f $ **FLOATING
C402 a_10108_4373# vssd1 0.648f $ **FLOATING
C403 cal_lut\[182\] vssd1 2.61f $ **FLOATING
C404 cal_lut\[134\] vssd1 3.34f $ **FLOATING
C405 a_9385_4373# vssd1 0.723f $ **FLOATING
C406 a_7439_4373# vssd1 0.698f $ **FLOATING
C407 a_7005_4551# vssd1 0.502f $ **FLOATING
C408 _0317_ vssd1 1.07f $ **FLOATING
C409 a_5687_4564# vssd1 0.524f $ **FLOATING
C410 a_5324_4373# vssd1 0.648f $ **FLOATING
C411 a_1407_4399# vssd1 0.698f $ **FLOATING
C412 a_25941_5321# vssd1 0.23f $ **FLOATING
C413 a_23117_4943# vssd1 0.203f $ **FLOATING
C414 a_21983_4943# vssd1 0.203f $ **FLOATING
C415 _0295_ vssd1 1.22f $ **FLOATING
C416 a_13629_4943# vssd1 0.23f $ **FLOATING
C417 _0311_ vssd1 0.947f $ **FLOATING
C418 a_8201_4943# vssd1 0.23f $ **FLOATING
C419 a_25523_5321# vssd1 0.581f $ **FLOATING
C420 a_25594_5220# vssd1 0.626f $ **FLOATING
C421 a_25394_5065# vssd1 1.43f $ **FLOATING
C422 a_25387_5161# vssd1 1.81f $ **FLOATING
C423 a_25103_5175# vssd1 0.609f $ **FLOATING
C424 a_25007_5175# vssd1 0.817f $ **FLOATING
C425 a_23763_4943# vssd1 1.2f $ **FLOATING
C426 _0478_ vssd1 0.854f $ **FLOATING
C427 cal_lut\[116\] vssd1 1.53f $ **FLOATING
C428 a_22988_4917# vssd1 0.655f $ **FLOATING
C429 cal_lut\[115\] vssd1 1.55f $ **FLOATING
C430 a_22523_5175# vssd1 0.619f $ **FLOATING
C431 a_21889_4943# vssd1 0.655f $ **FLOATING
C432 cal_lut\[151\] vssd1 3.08f $ **FLOATING
C433 _0687_ vssd1 0.801f $ **FLOATING
C434 a_20676_5059# vssd1 0.502f $ **FLOATING
C435 a_20175_5056# vssd1 0.619f $ **FLOATING
C436 cal_lut\[154\] vssd1 3.32f $ **FLOATING
C437 cal_lut\[156\] vssd1 2.13f $ **FLOATING
C438 a_18383_5175# vssd1 0.619f $ **FLOATING
C439 a_17927_4917# vssd1 0.698f $ **FLOATING
C440 a_17560_4917# vssd1 0.648f $ **FLOATING
C441 a_16127_5056# vssd1 0.619f $ **FLOATING
C442 cal_lut\[179\] vssd1 2.03f $ **FLOATING
C443 cal_lut\[178\] vssd1 2.26f $ **FLOATING
C444 a_15715_5175# vssd1 0.619f $ **FLOATING
C445 a_14795_5162# vssd1 0.524f $ **FLOATING
C446 a_14139_4943# vssd1 0.609f $ **FLOATING
C447 a_14307_4917# vssd1 0.817f $ **FLOATING
C448 a_13714_4943# vssd1 0.626f $ **FLOATING
C449 a_13882_4917# vssd1 0.581f $ **FLOATING
C450 a_13441_4949# vssd1 1.43f $ **FLOATING
C451 a_13275_4949# vssd1 1.81f $ **FLOATING
C452 a_12539_5056# vssd1 0.619f $ **FLOATING
C453 a_11660_5059# vssd1 0.502f $ **FLOATING
C454 a_10280_5059# vssd1 0.502f $ **FLOATING
C455 a_8711_4943# vssd1 0.609f $ **FLOATING
C456 a_8879_4917# vssd1 0.817f $ **FLOATING
C457 a_8286_4943# vssd1 0.626f $ **FLOATING
C458 a_8454_4917# vssd1 0.581f $ **FLOATING
C459 a_8013_4949# vssd1 1.43f $ **FLOATING
C460 _0145_ vssd1 0.872f $ **FLOATING
C461 a_7847_4949# vssd1 1.81f $ **FLOATING
C462 a_7571_4943# vssd1 0.524f $ **FLOATING
C463 _0318_ vssd1 0.945f $ **FLOATING
C464 a_7067_5162# vssd1 0.524f $ **FLOATING
C465 a_6637_5175# vssd1 0.502f $ **FLOATING
C466 a_5499_5249# vssd1 0.604f $ **FLOATING
C467 a_5323_4917# vssd1 0.508f $ **FLOATING
C468 a_4947_5249# vssd1 0.604f $ **FLOATING
C469 a_4771_4917# vssd1 0.508f $ **FLOATING
C470 _0160_ vssd1 0.922f $ **FLOATING
C471 a_25879_5487# vssd1 0.524f $ **FLOATING
C472 a_25389_5487# vssd1 0.23f $ **FLOATING
C473 a_19609_5487# vssd1 0.23f $ **FLOATING
C474 a_24971_5487# vssd1 0.581f $ **FLOATING
C475 a_25042_5461# vssd1 0.626f $ **FLOATING
C476 a_24835_5461# vssd1 1.81f $ **FLOATING
C477 a_24842_5761# vssd1 1.43f $ **FLOATING
C478 a_24551_5461# vssd1 0.609f $ **FLOATING
C479 a_24455_5639# vssd1 0.817f $ **FLOATING
C480 a_20775_5639# vssd1 0.619f $ **FLOATING
C481 a_20119_5853# vssd1 0.609f $ **FLOATING
C482 a_20287_5755# vssd1 0.817f $ **FLOATING
C483 a_19694_5853# vssd1 0.626f $ **FLOATING
C484 a_19862_5599# vssd1 0.581f $ **FLOATING
C485 a_19421_5487# vssd1 1.43f $ **FLOATING
C486 a_19255_5487# vssd1 1.81f $ **FLOATING
C487 cal_lut\[155\] vssd1 3.16f $ **FLOATING
C488 cal_lut\[131\] vssd1 4.13f $ **FLOATING
C489 a_16220_5737# vssd1 0.259f $ **FLOATING
C490 a_14733_5487# vssd1 0.23f $ **FLOATING
C491 a_18475_5639# vssd1 0.619f $ **FLOATING
C492 a_18015_5639# vssd1 0.619f $ **FLOATING
C493 a_17507_5487# vssd1 0.619f $ **FLOATING
C494 a_17095_5639# vssd1 0.619f $ **FLOATING
C495 a_16390_5487# vssd1 0.672f $ **FLOATING
C496 _0616_ vssd1 0.949f $ **FLOATING
C497 _0615_ vssd1 1.43f $ **FLOATING
C498 _0614_ vssd1 0.857f $ **FLOATING
C499 cal_lut\[149\] vssd1 3.37f $ **FLOATING
C500 a_15243_5853# vssd1 0.609f $ **FLOATING
C501 a_15411_5755# vssd1 0.817f $ **FLOATING
C502 a_14818_5853# vssd1 0.626f $ **FLOATING
C503 a_14986_5599# vssd1 0.581f $ **FLOATING
C504 a_14545_5487# vssd1 1.43f $ **FLOATING
C505 _0119_ vssd1 0.955f $ **FLOATING
C506 a_14379_5487# vssd1 1.81f $ **FLOATING
C507 _0118_ vssd1 1.15f $ **FLOATING
C508 a_13672_5737# vssd1 0.259f $ **FLOATING
C509 a_12079_5737# vssd1 0.333f $ **FLOATING
C510 a_10961_5487# vssd1 0.23f $ **FLOATING
C511 a_14151_5652# vssd1 0.524f $ **FLOATING
C512 cal_lut\[184\] vssd1 2.93f $ **FLOATING
C513 _0566_ vssd1 1.89f $ **FLOATING
C514 _0568_ vssd1 1.1f $ **FLOATING
C515 a_13241_5633# vssd1 0.672f $ **FLOATING
C516 a_12162_5737# vssd1 0.723f $ **FLOATING
C517 cal_lut\[129\] vssd1 1.49f $ **FLOATING
C518 cal_lut\[183\] vssd1 2.9f $ **FLOATING
C519 a_11471_5853# vssd1 0.609f $ **FLOATING
C520 a_11639_5755# vssd1 0.817f $ **FLOATING
C521 a_11046_5853# vssd1 0.626f $ **FLOATING
C522 a_11214_5599# vssd1 0.581f $ **FLOATING
C523 a_10773_5487# vssd1 1.43f $ **FLOATING
C524 a_10607_5487# vssd1 1.81f $ **FLOATING
C525 _0128_ vssd1 0.872f $ **FLOATING
C526 a_9595_5737# vssd1 0.333f $ **FLOATING
C527 _0328_ vssd1 0.863f $ **FLOATING
C528 cal_lut\[136\] vssd1 4.55f $ **FLOATING
C529 a_6453_5487# vssd1 0.23f $ **FLOATING
C530 a_10331_5487# vssd1 0.524f $ **FLOATING
C531 _0310_ vssd1 0.998f $ **FLOATING
C532 a_9678_5737# vssd1 0.723f $ **FLOATING
C533 cal_lut\[146\] vssd1 2.42f $ **FLOATING
C534 a_7891_5461# vssd1 0.604f $ **FLOATING
C535 a_7715_5461# vssd1 0.508f $ **FLOATING
C536 a_6963_5853# vssd1 0.609f $ **FLOATING
C537 a_7131_5755# vssd1 0.817f $ **FLOATING
C538 a_6538_5853# vssd1 0.626f $ **FLOATING
C539 a_6706_5599# vssd1 0.581f $ **FLOATING
C540 a_6265_5487# vssd1 1.43f $ **FLOATING
C541 _0135_ vssd1 1.19f $ **FLOATING
C542 a_6099_5487# vssd1 1.81f $ **FLOATING
C543 cal_lut\[137\] vssd1 7.21f $ **FLOATING
C544 a_4613_5487# vssd1 0.23f $ **FLOATING
C545 a_5123_5853# vssd1 0.609f $ **FLOATING
C546 a_5291_5755# vssd1 0.817f $ **FLOATING
C547 a_4698_5853# vssd1 0.626f $ **FLOATING
C548 a_4866_5599# vssd1 0.581f $ **FLOATING
C549 a_4425_5487# vssd1 1.43f $ **FLOATING
C550 a_4259_5487# vssd1 1.81f $ **FLOATING
C551 _0136_ vssd1 0.872f $ **FLOATING
C552 a_3983_5487# vssd1 0.524f $ **FLOATING
C553 _0319_ vssd1 1.43f $ **FLOATING
C554 _0345_ vssd1 1.2f $ **FLOATING
C555 _0159_ vssd1 1.41f $ **FLOATING
C556 a_22645_6031# vssd1 0.23f $ **FLOATING
C557 a_20572_6031# vssd1 0.259f $ **FLOATING
C558 _0113_ vssd1 1.16f $ **FLOATING
C559 _0301_ vssd1 1.27f $ **FLOATING
C560 _0300_ vssd1 1.31f $ **FLOATING
C561 cal_lut\[128\] vssd1 1.58f $ **FLOATING
C562 a_9397_6031# vssd1 0.23f $ **FLOATING
C563 a_7097_6031# vssd1 0.23f $ **FLOATING
C564 a_5073_6031# vssd1 0.23f $ **FLOATING
C565 _0346_ vssd1 0.725f $ **FLOATING
C566 a_26203_6250# vssd1 0.524f $ **FLOATING
C567 a_25783_6031# vssd1 0.508f $ **FLOATING
C568 cal_lut\[161\] vssd1 4.8f $ **FLOATING
C569 a_25603_6031# vssd1 0.604f $ **FLOATING
C570 a_25143_6031# vssd1 0.698f $ **FLOATING
C571 a_24771_6031# vssd1 0.508f $ **FLOATING
C572 a_24591_6031# vssd1 0.604f $ **FLOATING
C573 a_24315_6031# vssd1 0.524f $ **FLOATING
C574 _0344_ vssd1 0.647f $ **FLOATING
C575 a_23943_6031# vssd1 0.508f $ **FLOATING
C576 a_23763_6031# vssd1 0.604f $ **FLOATING
C577 a_23155_6031# vssd1 0.609f $ **FLOATING
C578 a_23323_6005# vssd1 0.817f $ **FLOATING
C579 a_22730_6031# vssd1 0.626f $ **FLOATING
C580 a_22898_6005# vssd1 0.581f $ **FLOATING
C581 a_22457_6037# vssd1 1.43f $ **FLOATING
C582 a_22291_6037# vssd1 1.81f $ **FLOATING
C583 a_21879_6250# vssd1 0.524f $ **FLOATING
C584 a_20943_6369# vssd1 0.56f $ **FLOATING
C585 cal_lut\[160\] vssd1 3.35f $ **FLOATING
C586 _0584_ vssd1 1.11f $ **FLOATING
C587 _0585_ vssd1 0.974f $ **FLOATING
C588 a_20141_6005# vssd1 0.672f $ **FLOATING
C589 a_18887_6031# vssd1 0.524f $ **FLOATING
C590 _0294_ vssd1 0.647f $ **FLOATING
C591 a_18515_6031# vssd1 0.508f $ **FLOATING
C592 a_18335_6031# vssd1 0.604f $ **FLOATING
C593 a_17599_6039# vssd1 0.648f $ **FLOATING
C594 a_16035_6144# vssd1 0.619f $ **FLOATING
C595 a_14651_6031# vssd1 0.508f $ **FLOATING
C596 cal_lut\[119\] vssd1 2.28f $ **FLOATING
C597 a_14471_6031# vssd1 0.604f $ **FLOATING
C598 a_13040_6147# vssd1 0.502f $ **FLOATING
C599 cal_lut\[118\] vssd1 5.21f $ **FLOATING
C600 a_12539_6144# vssd1 0.619f $ **FLOATING
C601 cal_lut\[130\] vssd1 2.19f $ **FLOATING
C602 a_9907_6031# vssd1 0.609f $ **FLOATING
C603 a_10075_6005# vssd1 0.817f $ **FLOATING
C604 a_9482_6031# vssd1 0.626f $ **FLOATING
C605 a_9650_6005# vssd1 0.581f $ **FLOATING
C606 a_9209_6037# vssd1 1.43f $ **FLOATING
C607 _0127_ vssd1 0.872f $ **FLOATING
C608 a_9043_6037# vssd1 1.81f $ **FLOATING
C609 a_8767_6031# vssd1 0.524f $ **FLOATING
C610 a_7607_6031# vssd1 0.609f $ **FLOATING
C611 a_7775_6005# vssd1 0.817f $ **FLOATING
C612 a_7182_6031# vssd1 0.626f $ **FLOATING
C613 a_7350_6005# vssd1 0.581f $ **FLOATING
C614 a_6909_6037# vssd1 1.43f $ **FLOATING
C615 a_6743_6037# vssd1 1.81f $ **FLOATING
C616 a_5583_6031# vssd1 0.609f $ **FLOATING
C617 a_5751_6005# vssd1 0.817f $ **FLOATING
C618 a_5158_6031# vssd1 0.626f $ **FLOATING
C619 a_5326_6005# vssd1 0.581f $ **FLOATING
C620 a_4885_6037# vssd1 1.43f $ **FLOATING
C621 _0137_ vssd1 0.872f $ **FLOATING
C622 a_4719_6037# vssd1 1.81f $ **FLOATING
C623 a_4443_6031# vssd1 0.524f $ **FLOATING
C624 _0320_ vssd1 1.26f $ **FLOATING
C625 temp1.capload\[1\].cap_56.HI vssd1 0.415f $ **FLOATING
C626 temp1.capload\[6\].cap.Y vssd1 0.281f $ **FLOATING
C627 a_1407_6031# vssd1 0.524f $ **FLOATING
C628 a_26141_6575# vssd1 0.23f $ **FLOATING
C629 a_26651_6941# vssd1 0.609f $ **FLOATING
C630 a_26819_6843# vssd1 0.817f $ **FLOATING
C631 a_26226_6941# vssd1 0.626f $ **FLOATING
C632 a_26394_6687# vssd1 0.581f $ **FLOATING
C633 a_25953_6575# vssd1 1.43f $ **FLOATING
C634 _0161_ vssd1 0.955f $ **FLOATING
C635 a_25787_6575# vssd1 1.81f $ **FLOATING
C636 a_24731_6740# vssd1 0.524f $ **FLOATING
C637 a_23211_6575# vssd1 0.648f $ **FLOATING
C638 a_21541_6575# vssd1 0.23f $ **FLOATING
C639 a_22887_6549# vssd1 0.604f $ **FLOATING
C640 a_22711_6549# vssd1 0.508f $ **FLOATING
C641 a_22051_6941# vssd1 0.609f $ **FLOATING
C642 a_22219_6843# vssd1 0.817f $ **FLOATING
C643 a_21626_6941# vssd1 0.626f $ **FLOATING
C644 a_21794_6687# vssd1 0.581f $ **FLOATING
C645 a_21353_6575# vssd1 1.43f $ **FLOATING
C646 _0157_ vssd1 1.08f $ **FLOATING
C647 a_21187_6575# vssd1 1.81f $ **FLOATING
C648 _0342_ vssd1 1.22f $ **FLOATING
C649 a_17493_6575# vssd1 0.23f $ **FLOATING
C650 a_20815_6941# vssd1 0.508f $ **FLOATING
C651 a_20635_6941# vssd1 0.604f $ **FLOATING
C652 a_18003_6941# vssd1 0.609f $ **FLOATING
C653 a_18171_6843# vssd1 0.817f $ **FLOATING
C654 a_17578_6941# vssd1 0.626f $ **FLOATING
C655 a_17746_6687# vssd1 0.581f $ **FLOATING
C656 a_17305_6575# vssd1 1.43f $ **FLOATING
C657 a_17139_6575# vssd1 1.81f $ **FLOATING
C658 _0309_ vssd1 1.28f $ **FLOATING
C659 a_8951_6825# vssd1 0.333f $ **FLOATING
C660 a_7741_6575# vssd1 0.23f $ **FLOATING
C661 a_14699_6549# vssd1 0.604f $ **FLOATING
C662 a_14523_6549# vssd1 0.508f $ **FLOATING
C663 a_13183_6575# vssd1 0.524f $ **FLOATING
C664 a_11247_6941# vssd1 0.508f $ **FLOATING
C665 a_11067_6941# vssd1 0.604f $ **FLOATING
C666 a_10379_6740# vssd1 0.524f $ **FLOATING
C667 a_9765_6727# vssd1 0.502f $ **FLOATING
C668 a_9034_6825# vssd1 0.723f $ **FLOATING
C669 cal_lut\[127\] vssd1 1.34f $ **FLOATING
C670 cal_lut\[145\] vssd1 2.16f $ **FLOATING
C671 a_8251_6941# vssd1 0.609f $ **FLOATING
C672 a_8419_6843# vssd1 0.817f $ **FLOATING
C673 a_7826_6941# vssd1 0.626f $ **FLOATING
C674 a_7994_6687# vssd1 0.581f $ **FLOATING
C675 a_7553_6575# vssd1 1.43f $ **FLOATING
C676 a_7387_6575# vssd1 1.81f $ **FLOATING
C677 _0144_ vssd1 1.1f $ **FLOATING
C678 temp1.capload\[1\].cap.Y vssd1 0.281f $ **FLOATING
C679 a_6879_6549# vssd1 0.604f $ **FLOATING
C680 a_6703_6549# vssd1 0.508f $ **FLOATING
C681 a_6375_6575# vssd1 0.524f $ **FLOATING
C682 _0327_ vssd1 0.725f $ **FLOATING
C683 a_1937_6549# vssd1 4.03f $ **FLOATING
C684 net56 vssd1 1.29f $ **FLOATING
C685 a_27337_7119# vssd1 0.23f $ **FLOATING
C686 a_24761_7119# vssd1 0.23f $ **FLOATING
C687 _0348_ vssd1 1.21f $ **FLOATING
C688 _0158_ vssd1 1.19f $ **FLOATING
C689 _0112_ vssd1 1.4f $ **FLOATING
C690 a_14825_7119# vssd1 0.23f $ **FLOATING
C691 _0306_ vssd1 1.22f $ **FLOATING
C692 a_11881_7119# vssd1 0.23f $ **FLOATING
C693 a_10317_7119# vssd1 0.23f $ **FLOATING
C694 _0126_ vssd1 1.28f $ **FLOATING
C695 a_6729_7119# vssd1 0.23f $ **FLOATING
C696 a_4413_7497# vssd1 0.23f $ **FLOATING
C697 a_27847_7119# vssd1 0.609f $ **FLOATING
C698 a_28015_7093# vssd1 0.817f $ **FLOATING
C699 a_27422_7119# vssd1 0.626f $ **FLOATING
C700 a_27590_7093# vssd1 0.581f $ **FLOATING
C701 a_27149_7125# vssd1 1.43f $ **FLOATING
C702 a_26983_7125# vssd1 1.81f $ **FLOATING
C703 a_26519_7119# vssd1 0.508f $ **FLOATING
C704 a_26339_7119# vssd1 0.604f $ **FLOATING
C705 a_25271_7119# vssd1 0.609f $ **FLOATING
C706 a_25439_7093# vssd1 0.817f $ **FLOATING
C707 a_24846_7119# vssd1 0.626f $ **FLOATING
C708 a_25014_7093# vssd1 0.581f $ **FLOATING
C709 a_24573_7125# vssd1 1.43f $ **FLOATING
C710 _0163_ vssd1 1.22f $ **FLOATING
C711 a_24407_7125# vssd1 1.81f $ **FLOATING
C712 a_24035_7119# vssd1 0.508f $ **FLOATING
C713 a_23855_7119# vssd1 0.604f $ **FLOATING
C714 a_23351_7338# vssd1 0.524f $ **FLOATING
C715 _0343_ vssd1 0.883f $ **FLOATING
C716 a_22431_7338# vssd1 0.524f $ **FLOATING
C717 a_19619_7119# vssd1 0.508f $ **FLOATING
C718 a_19439_7119# vssd1 0.604f $ **FLOATING
C719 a_18519_7119# vssd1 0.524f $ **FLOATING
C720 _0293_ vssd1 1.06f $ **FLOATING
C721 a_18107_7338# vssd1 0.524f $ **FLOATING
C722 a_17783_7119# vssd1 0.524f $ **FLOATING
C723 a_17415_7119# vssd1 0.698f $ **FLOATING
C724 a_16996_7235# vssd1 0.502f $ **FLOATING
C725 a_15943_7232# vssd1 0.619f $ **FLOATING
C726 a_15335_7119# vssd1 0.609f $ **FLOATING
C727 a_15503_7093# vssd1 0.817f $ **FLOATING
C728 a_14910_7119# vssd1 0.626f $ **FLOATING
C729 a_15078_7093# vssd1 0.581f $ **FLOATING
C730 a_14637_7125# vssd1 1.43f $ **FLOATING
C731 _0125_ vssd1 0.872f $ **FLOATING
C732 a_14471_7125# vssd1 1.81f $ **FLOATING
C733 a_14195_7119# vssd1 0.524f $ **FLOATING
C734 _0307_ vssd1 0.961f $ **FLOATING
C735 a_13592_7235# vssd1 0.502f $ **FLOATING
C736 cal_lut\[148\] vssd1 3.17f $ **FLOATING
C737 a_13139_7351# vssd1 0.619f $ **FLOATING
C738 a_12391_7119# vssd1 0.609f $ **FLOATING
C739 a_12559_7093# vssd1 0.817f $ **FLOATING
C740 a_11966_7119# vssd1 0.626f $ **FLOATING
C741 a_12134_7093# vssd1 0.581f $ **FLOATING
C742 a_11693_7125# vssd1 1.43f $ **FLOATING
C743 a_11527_7125# vssd1 1.81f $ **FLOATING
C744 a_10827_7119# vssd1 0.609f $ **FLOATING
C745 a_10995_7093# vssd1 0.817f $ **FLOATING
C746 a_10402_7119# vssd1 0.626f $ **FLOATING
C747 a_10570_7093# vssd1 0.581f $ **FLOATING
C748 a_10129_7125# vssd1 1.43f $ **FLOATING
C749 _0122_ vssd1 1.01f $ **FLOATING
C750 a_9963_7125# vssd1 1.81f $ **FLOATING
C751 _0308_ vssd1 0.758f $ **FLOATING
C752 a_8447_7338# vssd1 0.524f $ **FLOATING
C753 a_7980_7235# vssd1 0.502f $ **FLOATING
C754 a_7239_7119# vssd1 0.609f $ **FLOATING
C755 a_7407_7093# vssd1 0.817f $ **FLOATING
C756 a_6814_7119# vssd1 0.626f $ **FLOATING
C757 a_6982_7093# vssd1 0.581f $ **FLOATING
C758 a_6541_7125# vssd1 1.43f $ **FLOATING
C759 a_6375_7125# vssd1 1.81f $ **FLOATING
C760 a_4951_7338# vssd1 0.524f $ **FLOATING
C761 a_3995_7497# vssd1 0.581f $ **FLOATING
C762 a_4066_7396# vssd1 0.626f $ **FLOATING
C763 a_3866_7241# vssd1 1.43f $ **FLOATING
C764 a_3859_7337# vssd1 1.81f $ **FLOATING
C765 a_3575_7351# vssd1 0.609f $ **FLOATING
C766 a_3479_7351# vssd1 0.817f $ **FLOATING
C767 temp1.capload\[0\].cap_49.HI vssd1 0.415f $ **FLOATING
C768 temp1.capload\[5\].cap_60.HI vssd1 0.415f $ **FLOATING
C769 temp1.capload\[4\].cap_59.HI vssd1 0.415f $ **FLOATING
C770 temp1.capload\[8\].cap_63.HI vssd1 0.415f $ **FLOATING
C771 temp1.capload\[4\].cap.Y vssd1 0.281f $ **FLOATING
C772 net59 vssd1 0.97f $ **FLOATING
C773 temp1.capload\[14\].cap_54.HI vssd1 0.415f $ **FLOATING
C774 _0162_ vssd1 1.02f $ **FLOATING
C775 a_23197_7663# vssd1 0.23f $ **FLOATING
C776 a_26799_7663# vssd1 0.524f $ **FLOATING
C777 _0347_ vssd1 0.81f $ **FLOATING
C778 a_23707_8029# vssd1 0.609f $ **FLOATING
C779 a_23875_7931# vssd1 0.817f $ **FLOATING
C780 a_23282_8029# vssd1 0.626f $ **FLOATING
C781 a_23450_7775# vssd1 0.581f $ **FLOATING
C782 a_23009_7663# vssd1 1.43f $ **FLOATING
C783 _0109_ vssd1 0.994f $ **FLOATING
C784 a_22843_7663# vssd1 1.81f $ **FLOATING
C785 cal_lut\[159\] vssd1 2.65f $ **FLOATING
C786 _0292_ vssd1 2.02f $ **FLOATING
C787 a_20069_7663# vssd1 0.23f $ **FLOATING
C788 a_22291_7663# vssd1 0.619f $ **FLOATING
C789 a_21265_7815# vssd1 0.502f $ **FLOATING
C790 a_20579_8029# vssd1 0.609f $ **FLOATING
C791 a_20747_7931# vssd1 0.817f $ **FLOATING
C792 a_20154_8029# vssd1 0.626f $ **FLOATING
C793 a_20322_7775# vssd1 0.581f $ **FLOATING
C794 a_19881_7663# vssd1 1.43f $ **FLOATING
C795 a_19715_7663# vssd1 1.81f $ **FLOATING
C796 cal_lut\[144\] vssd1 7.26f $ **FLOATING
C797 a_19255_7663# vssd1 0.619f $ **FLOATING
C798 net32 vssd1 6.04f $ **FLOATING
C799 a_18673_7663# vssd1 0.23f $ **FLOATING
C800 _0111_ vssd1 0.955f $ **FLOATING
C801 a_18255_7663# vssd1 0.581f $ **FLOATING
C802 a_18326_7637# vssd1 0.626f $ **FLOATING
C803 a_18119_7637# vssd1 1.81f $ **FLOATING
C804 a_18126_7937# vssd1 1.43f $ **FLOATING
C805 a_17835_7637# vssd1 0.609f $ **FLOATING
C806 a_17739_7815# vssd1 0.817f $ **FLOATING
C807 a_17323_7663# vssd1 0.648f $ **FLOATING
C808 a_16340_7913# vssd1 0.259f $ **FLOATING
C809 a_14457_7663# vssd1 0.23f $ **FLOATING
C810 a_16757_7637# vssd1 0.713f $ **FLOATING
C811 cal_lut\[150\] vssd1 5.33f $ **FLOATING
C812 _0544_ vssd1 0.9f $ **FLOATING
C813 a_15909_7809# vssd1 0.672f $ **FLOATING
C814 a_14967_8029# vssd1 0.609f $ **FLOATING
C815 a_15135_7931# vssd1 0.817f $ **FLOATING
C816 a_14542_8029# vssd1 0.626f $ **FLOATING
C817 a_14710_7775# vssd1 0.581f $ **FLOATING
C818 a_14269_7663# vssd1 1.43f $ **FLOATING
C819 _0124_ vssd1 1.68f $ **FLOATING
C820 a_14103_7663# vssd1 1.81f $ **FLOATING
C821 a_13028_7913# vssd1 0.259f $ **FLOATING
C822 _0123_ vssd1 1.04f $ **FLOATING
C823 net26 vssd1 12.5f $ **FLOATING
C824 _0304_ vssd1 1.05f $ **FLOATING
C825 _0143_ vssd1 0.96f $ **FLOATING
C826 a_4889_7663# vssd1 0.23f $ **FLOATING
C827 cal_lut\[124\] vssd1 1.75f $ **FLOATING
C828 _0570_ vssd1 0.903f $ **FLOATING
C829 _0571_ vssd1 1.41f $ **FLOATING
C830 _0572_ vssd1 0.786f $ **FLOATING
C831 a_12597_7809# vssd1 0.672f $ **FLOATING
C832 a_12079_7663# vssd1 0.619f $ **FLOATING
C833 a_11527_7663# vssd1 0.524f $ **FLOATING
C834 _0305_ vssd1 1.27f $ **FLOATING
C835 a_10659_7637# vssd1 0.698f $ **FLOATING
C836 a_10235_8029# vssd1 0.508f $ **FLOATING
C837 a_10055_8029# vssd1 0.604f $ **FLOATING
C838 _0290_ vssd1 14.1f $ **FLOATING
C839 a_8999_7828# vssd1 0.524f $ **FLOATING
C840 a_6559_7663# vssd1 0.524f $ **FLOATING
C841 _0326_ vssd1 0.647f $ **FLOATING
C842 a_6187_8029# vssd1 0.508f $ **FLOATING
C843 a_6007_8029# vssd1 0.604f $ **FLOATING
C844 a_5399_8029# vssd1 0.609f $ **FLOATING
C845 a_5567_7931# vssd1 0.817f $ **FLOATING
C846 a_4974_8029# vssd1 0.626f $ **FLOATING
C847 a_5142_7775# vssd1 0.581f $ **FLOATING
C848 a_4701_7663# vssd1 1.43f $ **FLOATING
C849 _0142_ vssd1 0.955f $ **FLOATING
C850 a_4535_7663# vssd1 1.81f $ **FLOATING
C851 _0325_ vssd1 1.1f $ **FLOATING
C852 temp1.capload\[6\].cap_61.HI vssd1 0.415f $ **FLOATING
C853 temp1.capload\[5\].cap.Y vssd1 0.281f $ **FLOATING
C854 temp1.capload\[0\].cap.Y vssd1 0.281f $ **FLOATING
C855 temp1.capload\[8\].cap.Y vssd1 0.281f $ **FLOATING
C856 a_4163_8029# vssd1 0.508f $ **FLOATING
C857 cal_lut\[142\] vssd1 5.29f $ **FLOATING
C858 a_3983_8029# vssd1 0.604f $ **FLOATING
C859 a_3155_7663# vssd1 0.698f $ **FLOATING
C860 net60 vssd1 1.09f $ **FLOATING
C861 net49 vssd1 1.19f $ **FLOATING
C862 net63 vssd1 1.09f $ **FLOATING
C863 net61 vssd1 1.51f $ **FLOATING
C864 temp1.capload\[14\].cap.Y vssd1 0.281f $ **FLOATING
C865 net54 vssd1 1.1f $ **FLOATING
C866 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_ vssd1 7.15f $ **FLOATING
C867 a_25773_8207# vssd1 0.23f $ **FLOATING
C868 _0289_ vssd1 1.37f $ **FLOATING
C869 a_22185_8207# vssd1 0.23f $ **FLOATING
C870 _0583_ vssd1 1.64f $ **FLOATING
C871 _0110_ vssd1 0.975f $ **FLOATING
C872 _0545_ vssd1 0.857f $ **FLOATING
C873 a_11693_8207# vssd1 0.214f $ **FLOATING
C874 a_11609_8207# vssd1 0.167f $ **FLOATING
C875 a_8937_8207# vssd1 0.23f $ **FLOATING
C876 _0303_ vssd1 1.23f $ **FLOATING
C877 _0141_ vssd1 1.71f $ **FLOATING
C878 a_4259_8207# vssd1 0.227f $ **FLOATING
C879 a_27211_8513# vssd1 0.604f $ **FLOATING
C880 a_27035_8181# vssd1 0.508f $ **FLOATING
C881 a_26283_8207# vssd1 0.609f $ **FLOATING
C882 a_26451_8181# vssd1 0.817f $ **FLOATING
C883 a_25858_8207# vssd1 0.626f $ **FLOATING
C884 a_26026_8181# vssd1 0.581f $ **FLOATING
C885 a_25585_8213# vssd1 1.43f $ **FLOATING
C886 _0165_ vssd1 0.872f $ **FLOATING
C887 a_25419_8213# vssd1 1.81f $ **FLOATING
C888 net34 vssd1 9.98f $ **FLOATING
C889 a_25143_8207# vssd1 0.524f $ **FLOATING
C890 a_24635_8513# vssd1 0.604f $ **FLOATING
C891 a_24459_8181# vssd1 0.508f $ **FLOATING
C892 a_23804_8323# vssd1 0.502f $ **FLOATING
C893 cal_lut\[117\] vssd1 5.13f $ **FLOATING
C894 a_23351_8439# vssd1 0.619f $ **FLOATING
C895 a_22695_8207# vssd1 0.609f $ **FLOATING
C896 a_22863_8181# vssd1 0.817f $ **FLOATING
C897 a_22270_8207# vssd1 0.626f $ **FLOATING
C898 a_22438_8181# vssd1 0.581f $ **FLOATING
C899 a_21997_8213# vssd1 1.43f $ **FLOATING
C900 a_21831_8213# vssd1 1.81f $ **FLOATING
C901 net33 vssd1 12.7f $ **FLOATING
C902 a_21003_8320# vssd1 0.619f $ **FLOATING
C903 cal_lut\[111\] vssd1 1.31f $ **FLOATING
C904 cal_lut\[166\] vssd1 3.94f $ **FLOATING
C905 a_20499_8439# vssd1 0.619f $ **FLOATING
C906 a_19807_8207# vssd1 0.524f $ **FLOATING
C907 _0291_ vssd1 1.09f $ **FLOATING
C908 cal_lut\[113\] vssd1 2.32f $ **FLOATING
C909 a_18107_8439# vssd1 0.619f $ **FLOATING
C910 a_17651_8181# vssd1 0.698f $ **FLOATING
C911 a_16771_8320# vssd1 0.619f $ **FLOATING
C912 cal_lut\[143\] vssd1 6.92f $ **FLOATING
C913 a_15851_8320# vssd1 0.619f $ **FLOATING
C914 cal_lut\[180\] vssd1 6.15f $ **FLOATING
C915 a_14287_8320# vssd1 0.619f $ **FLOATING
C916 cal_lut\[112\] vssd1 2.86f $ **FLOATING
C917 _0441_ vssd1 14.4f $ **FLOATING
C918 a_11527_8207# vssd1 0.972f $ **FLOATING
C919 cal_lut\[123\] vssd1 2.03f $ **FLOATING
C920 a_10699_8320# vssd1 0.619f $ **FLOATING
C921 cal_lut\[135\] vssd1 4.74f $ **FLOATING
C922 a_9447_8207# vssd1 0.609f $ **FLOATING
C923 a_9615_8181# vssd1 0.817f $ **FLOATING
C924 a_9022_8207# vssd1 0.626f $ **FLOATING
C925 a_9190_8181# vssd1 0.581f $ **FLOATING
C926 a_8749_8213# vssd1 1.43f $ **FLOATING
C927 _0121_ vssd1 1.03f $ **FLOATING
C928 a_8583_8213# vssd1 1.81f $ **FLOATING
C929 net23 vssd1 12f $ **FLOATING
C930 a_8164_8323# vssd1 0.502f $ **FLOATING
C931 a_7704_8323# vssd1 0.502f $ **FLOATING
C932 _0299_ vssd1 11.1f $ **FLOATING
C933 a_6555_8207# vssd1 0.508f $ **FLOATING
C934 a_6375_8207# vssd1 0.604f $ **FLOATING
C935 _0324_ vssd1 0.725f $ **FLOATING
C936 a_5779_8426# vssd1 0.524f $ **FLOATING
C937 a_5359_8207# vssd1 0.508f $ **FLOATING
C938 a_5179_8207# vssd1 0.604f $ **FLOATING
C939 _0316_ vssd1 11.7f $ **FLOATING
C940 a_4912_8439# vssd1 0.535f $ **FLOATING
C941 net24 vssd1 7.62f $ **FLOATING
C942 a_4593_8439# vssd1 0.5f $ **FLOATING
C943 a_4406_8181# vssd1 0.578f $ **FLOATING
C944 a_4310_8439# vssd1 0.498f $ **FLOATING
C945 a_2489_8181# vssd1 4.03f $ **FLOATING
C946 temp1.capload\[12\].cap_52.HI vssd1 0.415f $ **FLOATING
C947 temp1.capload\[12\].cap.Y vssd1 0.281f $ **FLOATING
C948 net52 vssd1 0.821f $ **FLOATING
C949 a_1407_8207# vssd1 0.524f $ **FLOATING
C950 a_27245_8751# vssd1 0.23f $ **FLOATING
C951 a_27755_9117# vssd1 0.609f $ **FLOATING
C952 a_27923_9019# vssd1 0.817f $ **FLOATING
C953 a_27330_9117# vssd1 0.626f $ **FLOATING
C954 a_27498_8863# vssd1 0.581f $ **FLOATING
C955 a_27057_8751# vssd1 1.43f $ **FLOATING
C956 a_26891_8751# vssd1 1.81f $ **FLOATING
C957 _0166_ vssd1 0.872f $ **FLOATING
C958 _0350_ vssd1 1.14f $ **FLOATING
C959 a_24761_8751# vssd1 0.23f $ **FLOATING
C960 a_26615_8751# vssd1 0.524f $ **FLOATING
C961 _0351_ vssd1 0.973f $ **FLOATING
C962 _0341_ vssd1 10.5f $ **FLOATING
C963 a_26107_8725# vssd1 0.604f $ **FLOATING
C964 a_25931_8725# vssd1 0.508f $ **FLOATING
C965 a_25271_9117# vssd1 0.609f $ **FLOATING
C966 a_25439_9019# vssd1 0.817f $ **FLOATING
C967 a_24846_9117# vssd1 0.626f $ **FLOATING
C968 a_25014_8863# vssd1 0.581f $ **FLOATING
C969 a_24573_8751# vssd1 1.43f $ **FLOATING
C970 a_24407_8751# vssd1 1.81f $ **FLOATING
C971 _0164_ vssd1 0.911f $ **FLOATING
C972 cal_lut\[165\] vssd1 2.17f $ **FLOATING
C973 cal_lut\[153\] vssd1 3.93f $ **FLOATING
C974 _0108_ vssd1 1.29f $ **FLOATING
C975 cal_lut\[125\] vssd1 3.19f $ **FLOATING
C976 cal_lut\[120\] vssd1 6.17f $ **FLOATING
C977 cal_lut\[126\] vssd1 5.68f $ **FLOATING
C978 cal_lut\[132\] vssd1 6.05f $ **FLOATING
C979 _0569_ vssd1 1.93f $ **FLOATING
C980 _0573_ vssd1 1.25f $ **FLOATING
C981 a_24039_8751# vssd1 0.524f $ **FLOATING
C982 _0349_ vssd1 0.973f $ **FLOATING
C983 a_23395_8751# vssd1 0.619f $ **FLOATING
C984 a_22659_8751# vssd1 0.619f $ **FLOATING
C985 a_21371_8751# vssd1 0.524f $ **FLOATING
C986 _0288_ vssd1 0.797f $ **FLOATING
C987 a_20676_9001# vssd1 0.502f $ **FLOATING
C988 a_18795_8751# vssd1 0.524f $ **FLOATING
C989 a_18519_8751# vssd1 0.524f $ **FLOATING
C990 _0287_ vssd1 0.764f $ **FLOATING
C991 a_17871_9117# vssd1 0.508f $ **FLOATING
C992 a_17691_9117# vssd1 0.604f $ **FLOATING
C993 a_16771_8751# vssd1 0.619f $ **FLOATING
C994 a_15991_8903# vssd1 0.619f $ **FLOATING
C995 a_15483_8751# vssd1 0.619f $ **FLOATING
C996 a_15023_8751# vssd1 0.619f $ **FLOATING
C997 a_14163_8903# vssd1 0.56f $ **FLOATING
C998 a_13091_9001# vssd1 0.702f $ **FLOATING
C999 a_12723_8751# vssd1 0.524f $ **FLOATING
C1000 a_12141_8751# vssd1 0.23f $ **FLOATING
C1001 _0649_ vssd1 0.959f $ **FLOATING
C1002 a_9963_9001# vssd1 0.333f $ **FLOATING
C1003 a_7741_8751# vssd1 0.23f $ **FLOATING
C1004 a_11723_8751# vssd1 0.581f $ **FLOATING
C1005 a_11794_8725# vssd1 0.626f $ **FLOATING
C1006 a_11587_8725# vssd1 1.81f $ **FLOATING
C1007 a_11594_9025# vssd1 1.43f $ **FLOATING
C1008 a_11303_8725# vssd1 0.609f $ **FLOATING
C1009 a_11207_8903# vssd1 0.817f $ **FLOATING
C1010 a_10699_8751# vssd1 0.619f $ **FLOATING
C1011 a_10046_9001# vssd1 0.723f $ **FLOATING
C1012 cal_lut\[122\] vssd1 1.7f $ **FLOATING
C1013 a_9411_8751# vssd1 0.619f $ **FLOATING
C1014 a_8251_9117# vssd1 0.609f $ **FLOATING
C1015 a_8419_9019# vssd1 0.817f $ **FLOATING
C1016 a_7826_9117# vssd1 0.626f $ **FLOATING
C1017 a_7994_8863# vssd1 0.581f $ **FLOATING
C1018 a_7553_8751# vssd1 1.43f $ **FLOATING
C1019 a_7387_8751# vssd1 1.81f $ **FLOATING
C1020 a_6269_8751# vssd1 0.23f $ **FLOATING
C1021 a_6779_9117# vssd1 0.609f $ **FLOATING
C1022 a_6947_9019# vssd1 0.817f $ **FLOATING
C1023 a_6354_9117# vssd1 0.626f $ **FLOATING
C1024 a_6522_8863# vssd1 0.581f $ **FLOATING
C1025 a_6081_8751# vssd1 1.43f $ **FLOATING
C1026 a_5915_8751# vssd1 1.81f $ **FLOATING
C1027 cal_lut\[138\] vssd1 6.75f $ **FLOATING
C1028 cal_lut\[141\] vssd1 4.04f $ **FLOATING
C1029 temp1.capload\[2\].cap_57.HI vssd1 0.415f $ **FLOATING
C1030 a_4153_8751# vssd1 0.23f $ **FLOATING
C1031 cal_lut\[140\] vssd1 4.52f $ **FLOATING
C1032 a_5404_9001# vssd1 0.502f $ **FLOATING
C1033 a_4663_9117# vssd1 0.609f $ **FLOATING
C1034 a_4831_9019# vssd1 0.817f $ **FLOATING
C1035 a_4238_9117# vssd1 0.626f $ **FLOATING
C1036 a_4406_8863# vssd1 0.581f $ **FLOATING
C1037 a_3965_8751# vssd1 1.43f $ **FLOATING
C1038 a_3799_8751# vssd1 1.81f $ **FLOATING
C1039 _0140_ vssd1 1.1f $ **FLOATING
C1040 a_3325_8903# vssd1 0.502f $ **FLOATING
C1041 a_2971_8751# vssd1 0.524f $ **FLOATING
C1042 _0323_ vssd1 0.758f $ **FLOATING
C1043 temp1.capload\[2\].cap.Y vssd1 0.281f $ **FLOATING
C1044 temp1.capload\[15\].cap.Y vssd1 0.281f $ **FLOATING
C1045 temp1.capload\[13\].cap.Y vssd1 0.281f $ **FLOATING
C1046 temp1.capload\[9\].cap.Y vssd1 0.281f $ **FLOATING
C1047 net57 vssd1 0.821f $ **FLOATING
C1048 a_20069_9295# vssd1 0.23f $ **FLOATING
C1049 a_19225_9673# vssd1 0.23f $ **FLOATING
C1050 a_17033_9295# vssd1 0.23f $ **FLOATING
C1051 a_14776_9295# vssd1 0.259f $ **FLOATING
C1052 _0565_ vssd1 1.3f $ **FLOATING
C1053 a_13169_9295# vssd1 0.23f $ **FLOATING
C1054 _0278_ vssd1 0.931f $ **FLOATING
C1055 a_10129_9295# vssd1 0.214f $ **FLOATING
C1056 a_10045_9295# vssd1 0.167f $ **FLOATING
C1057 _0120_ vssd1 1.09f $ **FLOATING
C1058 _0139_ vssd1 1.13f $ **FLOATING
C1059 cal_lut\[139\] vssd1 3.27f $ **FLOATING
C1060 a_5165_9295# vssd1 0.23f $ **FLOATING
C1061 _0356_ vssd1 0.725f $ **FLOATING
C1062 a_27583_9514# vssd1 0.524f $ **FLOATING
C1063 a_27163_9295# vssd1 0.508f $ **FLOATING
C1064 a_26983_9295# vssd1 0.604f $ **FLOATING
C1065 a_24499_9295# vssd1 0.698f $ **FLOATING
C1066 a_22843_9295# vssd1 1.2f $ **FLOATING
C1067 a_21831_9408# vssd1 0.619f $ **FLOATING
C1068 a_21235_9514# vssd1 0.524f $ **FLOATING
C1069 a_20579_9295# vssd1 0.609f $ **FLOATING
C1070 a_20747_9269# vssd1 0.817f $ **FLOATING
C1071 a_20154_9295# vssd1 0.626f $ **FLOATING
C1072 a_20322_9269# vssd1 0.581f $ **FLOATING
C1073 a_19881_9301# vssd1 1.43f $ **FLOATING
C1074 _0107_ vssd1 1.54f $ **FLOATING
C1075 a_19715_9301# vssd1 1.81f $ **FLOATING
C1076 _0105_ vssd1 1.13f $ **FLOATING
C1077 a_18807_9673# vssd1 0.581f $ **FLOATING
C1078 a_18878_9572# vssd1 0.626f $ **FLOATING
C1079 a_18678_9417# vssd1 1.43f $ **FLOATING
C1080 a_18671_9513# vssd1 1.81f $ **FLOATING
C1081 a_18387_9527# vssd1 0.609f $ **FLOATING
C1082 a_18291_9527# vssd1 0.817f $ **FLOATING
C1083 a_17543_9295# vssd1 0.609f $ **FLOATING
C1084 a_17711_9269# vssd1 0.817f $ **FLOATING
C1085 a_17118_9295# vssd1 0.626f $ **FLOATING
C1086 a_17286_9269# vssd1 0.581f $ **FLOATING
C1087 a_16845_9301# vssd1 1.43f $ **FLOATING
C1088 a_16679_9301# vssd1 1.81f $ **FLOATING
C1089 a_16168_9411# vssd1 0.502f $ **FLOATING
C1090 a_15812_9269# vssd1 0.648f $ **FLOATING
C1091 cal_lut\[106\] vssd1 2.32f $ **FLOATING
C1092 a_15163_9527# vssd1 0.619f $ **FLOATING
C1093 _0562_ vssd1 0.779f $ **FLOATING
C1094 _0564_ vssd1 1.12f $ **FLOATING
C1095 a_14345_9269# vssd1 0.672f $ **FLOATING
C1096 a_13679_9295# vssd1 0.609f $ **FLOATING
C1097 a_13847_9269# vssd1 0.817f $ **FLOATING
C1098 a_13254_9295# vssd1 0.626f $ **FLOATING
C1099 a_13422_9269# vssd1 0.581f $ **FLOATING
C1100 a_12981_9301# vssd1 1.43f $ **FLOATING
C1101 _0099_ vssd1 1.03f $ **FLOATING
C1102 a_12815_9301# vssd1 1.81f $ **FLOATING
C1103 a_12259_9295# vssd1 0.508f $ **FLOATING
C1104 cal_lut\[99\] vssd1 2.13f $ **FLOATING
C1105 a_12079_9295# vssd1 0.604f $ **FLOATING
C1106 a_11527_9303# vssd1 0.648f $ **FLOATING
C1107 a_9963_9295# vssd1 0.972f $ **FLOATING
C1108 _0493_ vssd1 5.31f $ **FLOATING
C1109 cal_lut\[121\] vssd1 2.18f $ **FLOATING
C1110 _0693_ vssd1 0.876f $ **FLOATING
C1111 _0302_ vssd1 1.4f $ **FLOATING
C1112 a_7987_9514# vssd1 0.524f $ **FLOATING
C1113 _0322_ vssd1 1.09f $ **FLOATING
C1114 a_6607_9514# vssd1 0.524f $ **FLOATING
C1115 a_5675_9295# vssd1 0.609f $ **FLOATING
C1116 a_5843_9269# vssd1 0.817f $ **FLOATING
C1117 a_5250_9295# vssd1 0.626f $ **FLOATING
C1118 a_5418_9269# vssd1 0.581f $ **FLOATING
C1119 a_4977_9301# vssd1 1.43f $ **FLOATING
C1120 a_4811_9301# vssd1 1.81f $ **FLOATING
C1121 a_3707_9303# vssd1 0.648f $ **FLOATING
C1122 a_3339_9295# vssd1 0.698f $ **FLOATING
C1123 temp1.capload\[13\].cap_53.HI vssd1 0.415f $ **FLOATING
C1124 net53 vssd1 1.64f $ **FLOATING
C1125 temp1.capload\[15\].cap_55.HI vssd1 0.415f $ **FLOATING
C1126 net55 vssd1 1.22f $ **FLOATING
C1127 a_2235_9303# vssd1 0.648f $ **FLOATING
C1128 temp1.capload\[9\].cap_64.HI vssd1 0.415f $ **FLOATING
C1129 net64 vssd1 1.18f $ **FLOATING
C1130 temp1.capload\[3\].cap.Y vssd1 0.281f $ **FLOATING
C1131 temp1.capload\[7\].cap.Y vssd1 0.281f $ **FLOATING
C1132 a_27521_9839# vssd1 0.23f $ **FLOATING
C1133 a_28031_10205# vssd1 0.609f $ **FLOATING
C1134 a_28199_10107# vssd1 0.817f $ **FLOATING
C1135 a_27606_10205# vssd1 0.626f $ **FLOATING
C1136 a_27774_9951# vssd1 0.581f $ **FLOATING
C1137 a_27333_9839# vssd1 1.43f $ **FLOATING
C1138 _0170_ vssd1 0.955f $ **FLOATING
C1139 a_27167_9839# vssd1 1.81f $ **FLOATING
C1140 a_25957_9839# vssd1 0.23f $ **FLOATING
C1141 a_26467_10205# vssd1 0.609f $ **FLOATING
C1142 a_26635_10107# vssd1 0.817f $ **FLOATING
C1143 a_26042_10205# vssd1 0.626f $ **FLOATING
C1144 a_26210_9951# vssd1 0.581f $ **FLOATING
C1145 a_25769_9839# vssd1 1.43f $ **FLOATING
C1146 a_25603_9839# vssd1 1.81f $ **FLOATING
C1147 a_24630_10089# vssd1 0.333f $ **FLOATING
C1148 a_23792_10089# vssd1 0.259f $ **FLOATING
C1149 a_21081_9839# vssd1 0.23f $ **FLOATING
C1150 cal_lut\[170\] vssd1 2.27f $ **FLOATING
C1151 cal_lut\[164\] vssd1 2.76f $ **FLOATING
C1152 a_24473_9813# vssd1 0.723f $ **FLOATING
C1153 _0657_ vssd1 2.38f $ **FLOATING
C1154 _0658_ vssd1 1.21f $ **FLOATING
C1155 a_23361_9985# vssd1 0.672f $ **FLOATING
C1156 a_22875_9867# vssd1 0.56f $ **FLOATING
C1157 a_22247_9991# vssd1 0.619f $ **FLOATING
C1158 a_21591_10205# vssd1 0.609f $ **FLOATING
C1159 a_21759_10107# vssd1 0.817f $ **FLOATING
C1160 a_21166_10205# vssd1 0.626f $ **FLOATING
C1161 a_21334_9951# vssd1 0.581f $ **FLOATING
C1162 a_20893_9839# vssd1 1.43f $ **FLOATING
C1163 _0104_ vssd1 0.994f $ **FLOATING
C1164 a_20727_9839# vssd1 1.81f $ **FLOATING
C1165 cal_lut\[108\] vssd1 2.04f $ **FLOATING
C1166 cal_lut\[105\] vssd1 2.62f $ **FLOATING
C1167 _0285_ vssd1 1.32f $ **FLOATING
C1168 _0106_ vssd1 0.955f $ **FLOATING
C1169 a_15972_10089# vssd1 0.259f $ **FLOATING
C1170 _0098_ vssd1 1.25f $ **FLOATING
C1171 _0450_ vssd1 12.8f $ **FLOATING
C1172 _0699_ vssd1 2.12f $ **FLOATING
C1173 _0700_ vssd1 3.01f $ **FLOATING
C1174 _0138_ vssd1 1.33f $ **FLOATING
C1175 a_4153_9839# vssd1 0.23f $ **FLOATING
C1176 a_20267_9839# vssd1 0.619f $ **FLOATING
C1177 a_19333_9991# vssd1 0.502f $ **FLOATING
C1178 _0286_ vssd1 1.22f $ **FLOATING
C1179 a_17095_10004# vssd1 0.524f $ **FLOATING
C1180 net39 vssd1 12.8f $ **FLOATING
C1181 a_16731_9813# vssd1 0.698f $ **FLOATING
C1182 _0547_ vssd1 1.11f $ **FLOATING
C1183 _0548_ vssd1 1.24f $ **FLOATING
C1184 a_15541_9985# vssd1 0.672f $ **FLOATING
C1185 a_14375_10205# vssd1 0.508f $ **FLOATING
C1186 cal_lut\[100\] vssd1 1.67f $ **FLOATING
C1187 a_14195_10205# vssd1 0.604f $ **FLOATING
C1188 a_12263_9839# vssd1 0.524f $ **FLOATING
C1189 _0277_ vssd1 0.647f $ **FLOATING
C1190 a_11891_10205# vssd1 0.508f $ **FLOATING
C1191 a_11711_10205# vssd1 0.604f $ **FLOATING
C1192 a_10607_9839# vssd1 0.619f $ **FLOATING
C1193 a_9043_10089# vssd1 0.702f $ **FLOATING
C1194 a_7291_10205# vssd1 0.508f $ **FLOATING
C1195 a_7111_10205# vssd1 0.604f $ **FLOATING
C1196 _0321_ vssd1 1.21f $ **FLOATING
C1197 a_5871_10004# vssd1 0.524f $ **FLOATING
C1198 a_5451_10205# vssd1 0.508f $ **FLOATING
C1199 a_5271_10205# vssd1 0.604f $ **FLOATING
C1200 a_4663_10205# vssd1 0.609f $ **FLOATING
C1201 a_4831_10107# vssd1 0.817f $ **FLOATING
C1202 a_4238_10205# vssd1 0.626f $ **FLOATING
C1203 a_4406_9951# vssd1 0.581f $ **FLOATING
C1204 a_3965_9839# vssd1 1.43f $ **FLOATING
C1205 a_3799_9839# vssd1 1.81f $ **FLOATING
C1206 net3 vssd1 1.75f $ **FLOATING
C1207 a_3155_9839# vssd1 0.648f $ **FLOATING
C1208 temp1.capload\[11\].cap.Y vssd1 0.281f $ **FLOATING
C1209 a_2773_9991# vssd1 0.502f $ **FLOATING
C1210 net51 vssd1 0.96f $ **FLOATING
C1211 temp1.capload\[11\].cap_51.HI vssd1 0.415f $ **FLOATING
C1212 temp1.capload\[7\].cap_62.HI vssd1 0.415f $ **FLOATING
C1213 _0000_ vssd1 1.57f $ **FLOATING
C1214 a_1867_9839# vssd1 0.524f $ **FLOATING
C1215 _0837_ vssd1 1.02f $ **FLOATING
C1216 net62 vssd1 1.07f $ **FLOATING
C1217 _0169_ vssd1 0.975f $ **FLOATING
C1218 a_24262_10383# vssd1 0.333f $ **FLOATING
C1219 a_23683_10383# vssd1 0.167f $ **FLOATING
C1220 a_23481_10383# vssd1 0.214f $ **FLOATING
C1221 a_22596_10383# vssd1 0.259f $ **FLOATING
C1222 _0284_ vssd1 1.14f $ **FLOATING
C1223 a_17536_10383# vssd1 0.259f $ **FLOATING
C1224 a_11693_10383# vssd1 0.214f $ **FLOATING
C1225 a_11609_10383# vssd1 0.167f $ **FLOATING
C1226 a_10360_10383# vssd1 0.259f $ **FLOATING
C1227 a_8675_10383# vssd1 0.333f $ **FLOATING
C1228 a_14917_10383# vssd1 0.23f $ **FLOATING
C1229 a_27163_10383# vssd1 0.508f $ **FLOATING
C1230 cal_lut\[171\] vssd1 3.78f $ **FLOATING
C1231 a_26983_10383# vssd1 0.604f $ **FLOATING
C1232 _0355_ vssd1 0.725f $ **FLOATING
C1233 a_25927_10602# vssd1 0.524f $ **FLOATING
C1234 a_25507_10383# vssd1 0.508f $ **FLOATING
C1235 a_25327_10383# vssd1 0.604f $ **FLOATING
C1236 _0510_ vssd1 2.29f $ **FLOATING
C1237 cal_lut\[163\] vssd1 4.44f $ **FLOATING
C1238 a_24105_10357# vssd1 0.723f $ **FLOATING
C1239 _0695_ vssd1 0.564f $ **FLOATING
C1240 cal_lut\[109\] vssd1 2.27f $ **FLOATING
C1241 a_23355_10615# vssd1 0.972f $ **FLOATING
C1242 _0632_ vssd1 1.7f $ **FLOATING
C1243 _0633_ vssd1 1.14f $ **FLOATING
C1244 _0634_ vssd1 0.896f $ **FLOATING
C1245 a_22165_10357# vssd1 0.672f $ **FLOATING
C1246 a_20952_10499# vssd1 0.502f $ **FLOATING
C1247 _0283_ vssd1 17.4f $ **FLOATING
C1248 a_20032_10499# vssd1 0.502f $ **FLOATING
C1249 a_18659_10615# vssd1 0.619f $ **FLOATING
C1250 a_18055_10383# vssd1 0.508f $ **FLOATING
C1251 a_17875_10383# vssd1 0.604f $ **FLOATING
C1252 cal_lut\[107\] vssd1 2.05f $ **FLOATING
C1253 _0622_ vssd1 1.56f $ **FLOATING
C1254 _0623_ vssd1 1.2f $ **FLOATING
C1255 a_17105_10357# vssd1 0.672f $ **FLOATING
C1256 a_16035_10383# vssd1 0.524f $ **FLOATING
C1257 a_15427_10383# vssd1 0.609f $ **FLOATING
C1258 a_15595_10357# vssd1 0.817f $ **FLOATING
C1259 a_15002_10383# vssd1 0.626f $ **FLOATING
C1260 a_15170_10357# vssd1 0.581f $ **FLOATING
C1261 a_14729_10389# vssd1 1.43f $ **FLOATING
C1262 _0100_ vssd1 0.872f $ **FLOATING
C1263 a_14563_10389# vssd1 1.81f $ **FLOATING
C1264 a_14287_10383# vssd1 0.524f $ **FLOATING
C1265 _0279_ vssd1 1f $ **FLOATING
C1266 a_13367_10391# vssd1 0.648f $ **FLOATING
C1267 net1 vssd1 12.9f $ **FLOATING
C1268 a_12985_10615# vssd1 0.502f $ **FLOATING
C1269 _0659_ vssd1 5.55f $ **FLOATING
C1270 _0655_ vssd1 2.58f $ **FLOATING
C1271 _0654_ vssd1 0.865f $ **FLOATING
C1272 a_12310_10615# vssd1 0.702f $ **FLOATING
C1273 a_11527_10383# vssd1 0.972f $ **FLOATING
C1274 _0498_ vssd1 9.05f $ **FLOATING
C1275 cal_lut\[147\] vssd1 4.75f $ **FLOATING
C1276 _0653_ vssd1 1.03f $ **FLOATING
C1277 _0701_ vssd1 1.57f $ **FLOATING
C1278 _0696_ vssd1 6.09f $ **FLOATING
C1279 _0694_ vssd1 1.23f $ **FLOATING
C1280 _0697_ vssd1 0.826f $ **FLOATING
C1281 a_7097_10383# vssd1 0.23f $ **FLOATING
C1282 a_5517_10761# vssd1 0.23f $ **FLOATING
C1283 a_3953_10761# vssd1 0.23f $ **FLOATING
C1284 temp1.capload\[10\].cap.Y vssd1 0.281f $ **FLOATING
C1285 a_10746_10615# vssd1 0.702f $ **FLOATING
C1286 _0494_ vssd1 1.35f $ **FLOATING
C1287 a_9929_10357# vssd1 0.672f $ **FLOATING
C1288 a_8758_10383# vssd1 0.723f $ **FLOATING
C1289 cal_lut\[187\] vssd1 5.14f $ **FLOATING
C1290 a_7607_10383# vssd1 0.609f $ **FLOATING
C1291 a_7775_10357# vssd1 0.817f $ **FLOATING
C1292 a_7182_10383# vssd1 0.626f $ **FLOATING
C1293 a_7350_10357# vssd1 0.581f $ **FLOATING
C1294 a_6909_10389# vssd1 1.43f $ **FLOATING
C1295 a_6743_10389# vssd1 1.81f $ **FLOATING
C1296 _0375_ vssd1 1.04f $ **FLOATING
C1297 a_6055_10602# vssd1 0.524f $ **FLOATING
C1298 _0188_ vssd1 0.872f $ **FLOATING
C1299 a_5099_10761# vssd1 0.581f $ **FLOATING
C1300 a_5170_10660# vssd1 0.626f $ **FLOATING
C1301 a_4970_10505# vssd1 1.43f $ **FLOATING
C1302 a_4963_10601# vssd1 1.81f $ **FLOATING
C1303 a_4679_10615# vssd1 0.609f $ **FLOATING
C1304 a_4583_10615# vssd1 0.817f $ **FLOATING
C1305 a_3535_10761# vssd1 0.581f $ **FLOATING
C1306 a_3606_10660# vssd1 0.626f $ **FLOATING
C1307 a_3406_10505# vssd1 1.43f $ **FLOATING
C1308 a_3399_10601# vssd1 1.81f $ **FLOATING
C1309 a_3115_10615# vssd1 0.609f $ **FLOATING
C1310 a_2947_10615# vssd1 0.97f $ **FLOATING
C1311 a_1407_10383# vssd1 0.698f $ **FLOATING
C1312 _0357_ vssd1 0.895f $ **FLOATING
C1313 a_27491_11092# vssd1 0.524f $ **FLOATING
C1314 a_27071_11293# vssd1 0.508f $ **FLOATING
C1315 a_26891_11293# vssd1 0.604f $ **FLOATING
C1316 a_25757_10927# vssd1 0.23f $ **FLOATING
C1317 cal_lut\[177\] vssd1 8.15f $ **FLOATING
C1318 a_23959_11177# vssd1 0.167f $ **FLOATING
C1319 a_23757_11177# vssd1 0.214f $ **FLOATING
C1320 a_21081_10927# vssd1 0.23f $ **FLOATING
C1321 a_25339_10927# vssd1 0.581f $ **FLOATING
C1322 a_25410_10901# vssd1 0.626f $ **FLOATING
C1323 a_25203_10901# vssd1 1.81f $ **FLOATING
C1324 a_25210_11201# vssd1 1.43f $ **FLOATING
C1325 a_24919_10901# vssd1 0.609f $ **FLOATING
C1326 a_24823_11079# vssd1 0.817f $ **FLOATING
C1327 _0511_ vssd1 1.06f $ **FLOATING
C1328 _0509_ vssd1 1.49f $ **FLOATING
C1329 cal_lut\[110\] vssd1 5.06f $ **FLOATING
C1330 a_23631_11079# vssd1 0.972f $ **FLOATING
C1331 a_23151_10955# vssd1 0.56f $ **FLOATING
C1332 a_21591_11293# vssd1 0.609f $ **FLOATING
C1333 a_21759_11195# vssd1 0.817f $ **FLOATING
C1334 a_21166_11293# vssd1 0.626f $ **FLOATING
C1335 a_21334_11039# vssd1 0.581f $ **FLOATING
C1336 a_20893_10927# vssd1 1.43f $ **FLOATING
C1337 a_20727_10927# vssd1 1.81f $ **FLOATING
C1338 a_19609_10927# vssd1 0.23f $ **FLOATING
C1339 a_20119_11293# vssd1 0.609f $ **FLOATING
C1340 a_20287_11195# vssd1 0.817f $ **FLOATING
C1341 a_19694_11293# vssd1 0.626f $ **FLOATING
C1342 a_19862_11039# vssd1 0.581f $ **FLOATING
C1343 a_19421_10927# vssd1 1.43f $ **FLOATING
C1344 a_19255_10927# vssd1 1.81f $ **FLOATING
C1345 _0102_ vssd1 1.18f $ **FLOATING
C1346 cal_lut\[102\] vssd1 2.76f $ **FLOATING
C1347 a_16297_10927# vssd1 0.23f $ **FLOATING
C1348 a_18335_10927# vssd1 0.524f $ **FLOATING
C1349 _0281_ vssd1 0.81f $ **FLOATING
C1350 a_17907_10955# vssd1 0.56f $ **FLOATING
C1351 a_16807_11293# vssd1 0.609f $ **FLOATING
C1352 a_16975_11195# vssd1 0.817f $ **FLOATING
C1353 a_16382_11293# vssd1 0.626f $ **FLOATING
C1354 a_16550_11039# vssd1 0.581f $ **FLOATING
C1355 a_16109_10927# vssd1 1.43f $ **FLOATING
C1356 _0101_ vssd1 0.908f $ **FLOATING
C1357 a_15943_10927# vssd1 1.81f $ **FLOATING
C1358 _0280_ vssd1 0.959f $ **FLOATING
C1359 _0563_ vssd1 1.4f $ **FLOATING
C1360 _0567_ vssd1 3.06f $ **FLOATING
C1361 a_15524_11177# vssd1 0.502f $ **FLOATING
C1362 a_14611_11079# vssd1 0.619f $ **FLOATING
C1363 a_14151_11079# vssd1 0.619f $ **FLOATING
C1364 a_13245_10927# vssd1 0.23f $ **FLOATING
C1365 cal_lut\[98\] vssd1 2.42f $ **FLOATING
C1366 _0513_ vssd1 0.841f $ **FLOATING
C1367 _0512_ vssd1 7.18f $ **FLOATING
C1368 _0499_ vssd1 3.06f $ **FLOATING
C1369 _0497_ vssd1 0.703f $ **FLOATING
C1370 a_9043_11177# vssd1 0.333f $ **FLOATING
C1371 a_7741_10927# vssd1 0.23f $ **FLOATING
C1372 a_12827_10927# vssd1 0.581f $ **FLOATING
C1373 a_12898_10901# vssd1 0.626f $ **FLOATING
C1374 a_12691_10901# vssd1 1.81f $ **FLOATING
C1375 a_12698_11201# vssd1 1.43f $ **FLOATING
C1376 a_12407_10901# vssd1 0.609f $ **FLOATING
C1377 a_12311_11079# vssd1 0.817f $ **FLOATING
C1378 a_10851_11079# vssd1 0.56f $ **FLOATING
C1379 a_9779_11177# vssd1 0.702f $ **FLOATING
C1380 a_9126_11177# vssd1 0.723f $ **FLOATING
C1381 cal_lut\[188\] vssd1 3.24f $ **FLOATING
C1382 _0496_ vssd1 3.38f $ **FLOATING
C1383 a_8251_11293# vssd1 0.609f $ **FLOATING
C1384 a_8419_11195# vssd1 0.817f $ **FLOATING
C1385 a_7826_11293# vssd1 0.626f $ **FLOATING
C1386 a_7994_11039# vssd1 0.581f $ **FLOATING
C1387 a_7553_10927# vssd1 1.43f $ **FLOATING
C1388 a_7387_10927# vssd1 1.81f $ **FLOATING
C1389 _0187_ vssd1 0.955f $ **FLOATING
C1390 a_5809_10927# vssd1 0.23f $ **FLOATING
C1391 _0374_ vssd1 1.15f $ **FLOATING
C1392 a_7159_11092# vssd1 0.524f $ **FLOATING
C1393 a_6319_11293# vssd1 0.609f $ **FLOATING
C1394 a_6487_11195# vssd1 0.817f $ **FLOATING
C1395 a_5894_11293# vssd1 0.626f $ **FLOATING
C1396 a_6062_11039# vssd1 0.581f $ **FLOATING
C1397 a_5621_10927# vssd1 1.43f $ **FLOATING
C1398 a_5455_10927# vssd1 1.81f $ **FLOATING
C1399 _0201_ vssd1 0.955f $ **FLOATING
C1400 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_ vssd1 7.59f $ **FLOATING
C1401 a_5083_11293# vssd1 0.508f $ **FLOATING
C1402 cal_lut\[189\] vssd1 4.5f $ **FLOATING
C1403 a_4903_11293# vssd1 0.604f $ **FLOATING
C1404 a_3799_10927# vssd1 0.524f $ **FLOATING
C1405 _0392_ vssd1 0.719f $ **FLOATING
C1406 a_3288_11177# vssd1 0.502f $ **FLOATING
C1407 clknet_0_temp1.dcdel_capnode_notouch_ vssd1 5.97f $ **FLOATING
C1408 a_1477_10901# vssd1 4.03f $ **FLOATING
C1409 cal_lut\[172\] vssd1 7.62f $ **FLOATING
C1410 a_27521_11471# vssd1 0.23f $ **FLOATING
C1411 _0176_ vssd1 1.09f $ **FLOATING
C1412 a_22790_11471# vssd1 0.333f $ **FLOATING
C1413 a_21997_11471# vssd1 0.214f $ **FLOATING
C1414 a_21913_11471# vssd1 0.167f $ **FLOATING
C1415 a_21169_11471# vssd1 0.214f $ **FLOATING
C1416 a_21085_11471# vssd1 0.167f $ **FLOATING
C1417 _0103_ vssd1 1.24f $ **FLOATING
C1418 _0097_ vssd1 1.13f $ **FLOATING
C1419 a_10041_11471# vssd1 0.23f $ **FLOATING
C1420 _0037_ vssd1 1.06f $ **FLOATING
C1421 _0189_ vssd1 1.02f $ **FLOATING
C1422 a_28031_11471# vssd1 0.609f $ **FLOATING
C1423 a_28199_11445# vssd1 0.817f $ **FLOATING
C1424 a_27606_11471# vssd1 0.626f $ **FLOATING
C1425 a_27774_11445# vssd1 0.581f $ **FLOATING
C1426 a_27333_11477# vssd1 1.43f $ **FLOATING
C1427 _0171_ vssd1 0.961f $ **FLOATING
C1428 a_27167_11477# vssd1 1.81f $ **FLOATING
C1429 a_25419_11471# vssd1 0.524f $ **FLOATING
C1430 _0362_ vssd1 0.647f $ **FLOATING
C1431 a_25047_11471# vssd1 0.508f $ **FLOATING
C1432 a_24867_11471# vssd1 0.604f $ **FLOATING
C1433 _0451_ vssd1 19.6f $ **FLOATING
C1434 a_22633_11445# vssd1 0.723f $ **FLOATING
C1435 a_21831_11471# vssd1 0.972f $ **FLOATING
C1436 cal_lut\[157\] vssd1 5.09f $ **FLOATING
C1437 cal_lut\[103\] vssd1 2.21f $ **FLOATING
C1438 a_21003_11471# vssd1 0.972f $ **FLOATING
C1439 cal_lut\[158\] vssd1 4.44f $ **FLOATING
C1440 _0449_ vssd1 4f $ **FLOATING
C1441 cal_lut\[104\] vssd1 1.8f $ **FLOATING
C1442 _0457_ vssd1 1.98f $ **FLOATING
C1443 a_20175_11471# vssd1 0.524f $ **FLOATING
C1444 _0282_ vssd1 1.2f $ **FLOATING
C1445 a_19071_11584# vssd1 0.619f $ **FLOATING
C1446 cal_lut\[186\] vssd1 8.53f $ **FLOATING
C1447 a_12815_11471# vssd1 0.524f $ **FLOATING
C1448 _0276_ vssd1 1.16f $ **FLOATING
C1449 a_11891_11471# vssd1 0.508f $ **FLOATING
C1450 cal_lut\[39\] vssd1 1.84f $ **FLOATING
C1451 a_11711_11471# vssd1 0.604f $ **FLOATING
C1452 a_10551_11471# vssd1 0.609f $ **FLOATING
C1453 a_10719_11445# vssd1 0.817f $ **FLOATING
C1454 a_10126_11471# vssd1 0.626f $ **FLOATING
C1455 a_10294_11445# vssd1 0.581f $ **FLOATING
C1456 a_9853_11477# vssd1 1.43f $ **FLOATING
C1457 _0038_ vssd1 0.872f $ **FLOATING
C1458 a_9687_11477# vssd1 1.81f $ **FLOATING
C1459 a_9411_11471# vssd1 0.524f $ **FLOATING
C1460 _0882_ vssd1 0.686f $ **FLOATING
C1461 a_8947_11471# vssd1 0.508f $ **FLOATING
C1462 cal_lut\[38\] vssd1 1.39f $ **FLOATING
C1463 a_8767_11471# vssd1 0.604f $ **FLOATING
C1464 a_8351_11777# vssd1 0.604f $ **FLOATING
C1465 a_8175_11445# vssd1 0.508f $ **FLOATING
C1466 _0881_ vssd1 0.647f $ **FLOATING
C1467 a_7895_11690# vssd1 0.524f $ **FLOATING
C1468 a_6603_11777# vssd1 0.604f $ **FLOATING
C1469 cal_lut\[190\] vssd1 5.08f $ **FLOATING
C1470 a_6427_11445# vssd1 0.508f $ **FLOATING
C1471 a_5639_11471# vssd1 0.524f $ **FLOATING
C1472 _0376_ vssd1 0.961f $ **FLOATING
C1473 a_5143_11445# vssd1 0.788f $ **FLOATING
C1474 a_4885_11445# vssd1 0.794f $ **FLOATING
C1475 a_4789_11703# vssd1 0.553f $ **FLOATING
C1476 net75 vssd1 0.669f $ **FLOATING
C1477 a_3877_11703# vssd1 0.502f $ **FLOATING
C1478 temp1.capload\[3\].cap_58.HI vssd1 0.415f $ **FLOATING
C1479 net58 vssd1 2.04f $ **FLOATING
C1480 net50 vssd1 1.52f $ **FLOATING
C1481 _0391_ vssd1 1.22f $ **FLOATING
C1482 a_2309_11791# vssd1 0.211f $ **FLOATING
C1483 a_2071_11791# vssd1 0.706f $ **FLOATING
C1484 temp1.capload\[10\].cap_50.HI vssd1 0.415f $ **FLOATING
C1485 a_27351_12015# vssd1 0.524f $ **FLOATING
C1486 _0358_ vssd1 1.02f $ **FLOATING
C1487 a_26309_12015# vssd1 0.23f $ **FLOATING
C1488 cal_lut\[176\] vssd1 2.47f $ **FLOATING
C1489 a_20112_12265# vssd1 0.259f $ **FLOATING
C1490 a_18272_12265# vssd1 0.259f $ **FLOATING
C1491 a_14855_12265# vssd1 0.388f $ **FLOATING
C1492 _0175_ vssd1 1.24f $ **FLOATING
C1493 a_25891_12015# vssd1 0.581f $ **FLOATING
C1494 a_25962_11989# vssd1 0.626f $ **FLOATING
C1495 a_25755_11989# vssd1 1.81f $ **FLOATING
C1496 a_25762_12289# vssd1 1.43f $ **FLOATING
C1497 a_25471_11989# vssd1 0.609f $ **FLOATING
C1498 a_25375_12167# vssd1 0.817f $ **FLOATING
C1499 a_25051_12015# vssd1 0.524f $ **FLOATING
C1500 a_23671_12015# vssd1 0.524f $ **FLOATING
C1501 a_20943_12043# vssd1 0.56f $ **FLOATING
C1502 _0444_ vssd1 5.61f $ **FLOATING
C1503 cal_lut\[162\] vssd1 6.29f $ **FLOATING
C1504 _0524_ vssd1 1.07f $ **FLOATING
C1505 a_19681_12161# vssd1 0.672f $ **FLOATING
C1506 a_18645_12043# vssd1 0.713f $ **FLOATING
C1507 _0502_ vssd1 9.38f $ **FLOATING
C1508 cal_lut\[185\] vssd1 7.36f $ **FLOATING
C1509 _0607_ vssd1 2.14f $ **FLOATING
C1510 a_17841_12161# vssd1 0.672f $ **FLOATING
C1511 a_17088_12265# vssd1 0.502f $ **FLOATING
C1512 a_15943_12015# vssd1 0.619f $ **FLOATING
C1513 a_15299_12015# vssd1 0.619f $ **FLOATING
C1514 _0514_ vssd1 11.8f $ **FLOATING
C1515 _0440_ vssd1 12.6f $ **FLOATING
C1516 a_6729_12015# vssd1 0.23f $ **FLOATING
C1517 a_14156_11989# vssd1 0.648f $ **FLOATING
C1518 a_12815_12015# vssd1 0.524f $ **FLOATING
C1519 _0378_ vssd1 0.686f $ **FLOATING
C1520 a_12351_12381# vssd1 0.508f $ **FLOATING
C1521 cal_lut\[191\] vssd1 4.64f $ **FLOATING
C1522 a_12171_12381# vssd1 0.604f $ **FLOATING
C1523 a_7239_12381# vssd1 0.609f $ **FLOATING
C1524 a_7407_12283# vssd1 0.817f $ **FLOATING
C1525 a_6814_12381# vssd1 0.626f $ **FLOATING
C1526 a_6982_12127# vssd1 0.581f $ **FLOATING
C1527 a_6541_12015# vssd1 1.43f $ **FLOATING
C1528 a_6375_12015# vssd1 1.81f $ **FLOATING
C1529 _0190_ vssd1 0.872f $ **FLOATING
C1530 a_2139_12265# vssd1 0.253f $ **FLOATING
C1531 a_6099_12015# vssd1 0.524f $ **FLOATING
C1532 _0377_ vssd1 0.934f $ **FLOATING
C1533 a_3869_11989# vssd1 4.03f $ **FLOATING
C1534 a_2419_12015# vssd1 1.2f $ **FLOATING
C1535 a_1921_11989# vssd1 0.55f $ **FLOATING
C1536 a_1407_12015# vssd1 0.524f $ **FLOATING
C1537 a_27521_12559# vssd1 0.23f $ **FLOATING
C1538 _0361_ vssd1 0.911f $ **FLOATING
C1539 a_24653_12937# vssd1 0.23f $ **FLOATING
C1540 _0856_ vssd1 0.975f $ **FLOATING
C1541 a_22054_12559# vssd1 0.333f $ **FLOATING
C1542 a_20756_12559# vssd1 0.259f $ **FLOATING
C1543 _0683_ vssd1 1.14f $ **FLOATING
C1544 net19 vssd1 7.11f $ **FLOATING
C1545 a_17168_12559# vssd1 0.259f $ **FLOATING
C1546 a_18229_12559# vssd1 0.23f $ **FLOATING
C1547 a_15469_12559# vssd1 0.23f $ **FLOATING
C1548 cal_lut\[192\] vssd1 1.29f $ **FLOATING
C1549 a_13353_12559# vssd1 0.23f $ **FLOATING
C1550 a_9033_12559# vssd1 0.206f $ **FLOATING
C1551 _0698_ vssd1 1.87f $ **FLOATING
C1552 a_6729_12559# vssd1 0.23f $ **FLOATING
C1553 a_3335_12559# vssd1 0.253f $ **FLOATING
C1554 a_3969_12559# vssd1 0.23f $ **FLOATING
C1555 a_1761_12559# vssd1 0.23f $ **FLOATING
C1556 a_28031_12559# vssd1 0.609f $ **FLOATING
C1557 a_28199_12533# vssd1 0.817f $ **FLOATING
C1558 a_27606_12559# vssd1 0.626f $ **FLOATING
C1559 a_27774_12533# vssd1 0.581f $ **FLOATING
C1560 a_27333_12565# vssd1 1.43f $ **FLOATING
C1561 _0172_ vssd1 1.01f $ **FLOATING
C1562 a_27167_12565# vssd1 1.81f $ **FLOATING
C1563 a_26063_12559# vssd1 0.524f $ **FLOATING
C1564 a_25463_12865# vssd1 0.604f $ **FLOATING
C1565 a_25287_12533# vssd1 0.508f $ **FLOATING
C1566 _0014_ vssd1 1.36f $ **FLOATING
C1567 a_24235_12937# vssd1 0.581f $ **FLOATING
C1568 a_24306_12836# vssd1 0.626f $ **FLOATING
C1569 a_24106_12681# vssd1 1.43f $ **FLOATING
C1570 a_24099_12777# vssd1 1.81f $ **FLOATING
C1571 a_23815_12791# vssd1 0.609f $ **FLOATING
C1572 a_23719_12791# vssd1 0.817f $ **FLOATING
C1573 a_23207_12559# vssd1 0.508f $ **FLOATING
C1574 a_23027_12559# vssd1 0.604f $ **FLOATING
C1575 a_21897_12533# vssd1 0.723f $ **FLOATING
C1576 a_21095_12559# vssd1 0.524f $ **FLOATING
C1577 _0506_ vssd1 3.42f $ **FLOATING
C1578 cal_lut\[114\] vssd1 4.77f $ **FLOATING
C1579 _0535_ vssd1 3.03f $ **FLOATING
C1580 a_20325_12533# vssd1 0.672f $ **FLOATING
C1581 a_18739_12559# vssd1 0.609f $ **FLOATING
C1582 a_18907_12533# vssd1 0.817f $ **FLOATING
C1583 a_18314_12559# vssd1 0.626f $ **FLOATING
C1584 a_18482_12533# vssd1 0.581f $ **FLOATING
C1585 a_18041_12565# vssd1 1.43f $ **FLOATING
C1586 _0017_ vssd1 0.93f $ **FLOATING
C1587 a_17875_12565# vssd1 1.81f $ **FLOATING
C1588 a_17599_12559# vssd1 0.524f $ **FLOATING
C1589 _0859_ vssd1 0.986f $ **FLOATING
C1590 cal_lut\[17\] vssd1 1.94f $ **FLOATING
C1591 _0603_ vssd1 3.68f $ **FLOATING
C1592 a_16737_12533# vssd1 0.672f $ **FLOATING
C1593 a_15979_12559# vssd1 0.609f $ **FLOATING
C1594 a_16147_12533# vssd1 0.817f $ **FLOATING
C1595 a_15554_12559# vssd1 0.626f $ **FLOATING
C1596 a_15722_12533# vssd1 0.581f $ **FLOATING
C1597 a_15281_12565# vssd1 1.43f $ **FLOATING
C1598 _0016_ vssd1 0.872f $ **FLOATING
C1599 a_15115_12565# vssd1 1.81f $ **FLOATING
C1600 a_14839_12559# vssd1 0.524f $ **FLOATING
C1601 a_13863_12559# vssd1 0.609f $ **FLOATING
C1602 a_14031_12533# vssd1 0.817f $ **FLOATING
C1603 a_13438_12559# vssd1 0.626f $ **FLOATING
C1604 a_13606_12533# vssd1 0.581f $ **FLOATING
C1605 a_13165_12565# vssd1 1.43f $ **FLOATING
C1606 _0191_ vssd1 1.08f $ **FLOATING
C1607 a_12999_12565# vssd1 1.81f $ **FLOATING
C1608 _0660_ vssd1 1.55f $ **FLOATING
C1609 _0650_ vssd1 2.51f $ **FLOATING
C1610 a_11707_12559# vssd1 0.508f $ **FLOATING
C1611 a_11527_12559# vssd1 0.604f $ **FLOATING
C1612 a_9595_12559# vssd1 0.524f $ **FLOATING
C1613 a_8951_12559# vssd1 0.804f $ **FLOATING
C1614 a_7895_12778# vssd1 0.524f $ **FLOATING
C1615 a_7239_12559# vssd1 0.609f $ **FLOATING
C1616 a_7407_12533# vssd1 0.817f $ **FLOATING
C1617 a_6814_12559# vssd1 0.626f $ **FLOATING
C1618 a_6982_12533# vssd1 0.581f $ **FLOATING
C1619 a_6541_12565# vssd1 1.43f $ **FLOATING
C1620 a_6375_12565# vssd1 1.81f $ **FLOATING
C1621 net27 vssd1 9.48f $ **FLOATING
C1622 a_6007_12559# vssd1 0.524f $ **FLOATING
C1623 a_5644_12533# vssd1 0.598f $ **FLOATING
C1624 a_5404_12797# vssd1 0.62f $ **FLOATING
C1625 a_5278_12533# vssd1 0.58f $ **FLOATING
C1626 a_4479_12559# vssd1 0.609f $ **FLOATING
C1627 a_4647_12533# vssd1 0.97f $ **FLOATING
C1628 a_4054_12559# vssd1 0.626f $ **FLOATING
C1629 a_4222_12533# vssd1 0.581f $ **FLOATING
C1630 a_3781_12565# vssd1 1.43f $ **FLOATING
C1631 _0203_ vssd1 1.06f $ **FLOATING
C1632 a_3615_12565# vssd1 1.81f $ **FLOATING
C1633 _0396_ vssd1 1.19f $ **FLOATING
C1634 _0395_ vssd1 1.58f $ **FLOATING
C1635 a_3117_12533# vssd1 0.55f $ **FLOATING
C1636 a_2271_12559# vssd1 0.609f $ **FLOATING
C1637 a_2439_12533# vssd1 0.97f $ **FLOATING
C1638 a_1846_12559# vssd1 0.626f $ **FLOATING
C1639 a_2014_12533# vssd1 0.581f $ **FLOATING
C1640 a_1573_12565# vssd1 1.43f $ **FLOATING
C1641 _0200_ vssd1 1.04f $ **FLOATING
C1642 a_1407_12565# vssd1 1.81f $ **FLOATING
C1643 a_27903_13103# vssd1 0.524f $ **FLOATING
C1644 _0359_ vssd1 0.647f $ **FLOATING
C1645 a_27531_13469# vssd1 0.508f $ **FLOATING
C1646 a_27351_13469# vssd1 0.604f $ **FLOATING
C1647 a_26861_13103# vssd1 0.23f $ **FLOATING
C1648 cal_lut\[175\] vssd1 3.02f $ **FLOATING
C1649 _0174_ vssd1 1.23f $ **FLOATING
C1650 a_26443_13103# vssd1 0.581f $ **FLOATING
C1651 a_26514_13077# vssd1 0.626f $ **FLOATING
C1652 a_26307_13077# vssd1 1.81f $ **FLOATING
C1653 a_26314_13377# vssd1 1.43f $ **FLOATING
C1654 a_26023_13077# vssd1 0.609f $ **FLOATING
C1655 a_25927_13255# vssd1 0.817f $ **FLOATING
C1656 a_25389_13103# vssd1 0.23f $ **FLOATING
C1657 cal_lut\[14\] vssd1 1.82f $ **FLOATING
C1658 a_22461_13103# vssd1 0.23f $ **FLOATING
C1659 a_24971_13103# vssd1 0.581f $ **FLOATING
C1660 a_25042_13077# vssd1 0.626f $ **FLOATING
C1661 a_24835_13077# vssd1 1.81f $ **FLOATING
C1662 a_24842_13377# vssd1 1.43f $ **FLOATING
C1663 a_24551_13077# vssd1 0.609f $ **FLOATING
C1664 a_24455_13255# vssd1 0.817f $ **FLOATING
C1665 a_23759_13469# vssd1 0.508f $ **FLOATING
C1666 cal_lut\[15\] vssd1 2.82f $ **FLOATING
C1667 a_23579_13469# vssd1 0.604f $ **FLOATING
C1668 a_22971_13469# vssd1 0.609f $ **FLOATING
C1669 a_23139_13371# vssd1 0.817f $ **FLOATING
C1670 a_22546_13469# vssd1 0.626f $ **FLOATING
C1671 a_22714_13215# vssd1 0.581f $ **FLOATING
C1672 a_22273_13103# vssd1 1.43f $ **FLOATING
C1673 a_22107_13103# vssd1 1.81f $ **FLOATING
C1674 net36 vssd1 11.4f $ **FLOATING
C1675 a_20848_13353# vssd1 0.259f $ **FLOATING
C1676 _0445_ vssd1 10.3f $ **FLOATING
C1677 cal_lut\[173\] vssd1 6.36f $ **FLOATING
C1678 _0608_ vssd1 1.47f $ **FLOATING
C1679 _0604_ vssd1 0.975f $ **FLOATING
C1680 _0601_ vssd1 0.857f $ **FLOATING
C1681 _0858_ vssd1 1.09f $ **FLOATING
C1682 a_12617_13103# vssd1 0.23f $ **FLOATING
C1683 a_21735_13469# vssd1 0.508f $ **FLOATING
C1684 a_21555_13469# vssd1 0.604f $ **FLOATING
C1685 cal_lut\[18\] vssd1 2.14f $ **FLOATING
C1686 _0528_ vssd1 1.92f $ **FLOATING
C1687 a_20417_13249# vssd1 0.672f $ **FLOATING
C1688 _0538_ vssd1 0.849f $ **FLOATING
C1689 _0529_ vssd1 0.915f $ **FLOATING
C1690 _0525_ vssd1 1.06f $ **FLOATING
C1691 a_19333_13255# vssd1 0.502f $ **FLOATING
C1692 a_18597_13077# vssd1 0.713f $ **FLOATING
C1693 a_17187_13255# vssd1 0.619f $ **FLOATING
C1694 a_16373_13077# vssd1 0.858f $ **FLOATING
C1695 a_15071_13268# vssd1 0.524f $ **FLOATING
C1696 a_14604_13353# vssd1 0.502f $ **FLOATING
C1697 a_13127_13469# vssd1 0.609f $ **FLOATING
C1698 a_13295_13371# vssd1 0.817f $ **FLOATING
C1699 a_12702_13469# vssd1 0.626f $ **FLOATING
C1700 a_12870_13215# vssd1 0.581f $ **FLOATING
C1701 a_12429_13103# vssd1 1.43f $ **FLOATING
C1702 a_12263_13103# vssd1 1.81f $ **FLOATING
C1703 _0652_ vssd1 1.83f $ **FLOATING
C1704 a_11509_13353# vssd1 0.214f $ **FLOATING
C1705 a_11425_13353# vssd1 0.167f $ **FLOATING
C1706 a_10041_13103# vssd1 0.23f $ **FLOATING
C1707 a_11343_13103# vssd1 0.972f $ **FLOATING
C1708 cal_lut\[21\] vssd1 1.68f $ **FLOATING
C1709 _0651_ vssd1 2.69f $ **FLOATING
C1710 a_10551_13469# vssd1 0.609f $ **FLOATING
C1711 a_10719_13371# vssd1 0.817f $ **FLOATING
C1712 a_10126_13469# vssd1 0.626f $ **FLOATING
C1713 a_10294_13215# vssd1 0.581f $ **FLOATING
C1714 a_9853_13103# vssd1 1.43f $ **FLOATING
C1715 _0020_ vssd1 0.977f $ **FLOATING
C1716 a_9687_13103# vssd1 1.81f $ **FLOATING
C1717 _0504_ vssd1 1.58f $ **FLOATING
C1718 a_9117_13353# vssd1 0.214f $ **FLOATING
C1719 a_9033_13353# vssd1 0.167f $ **FLOATING
C1720 a_7741_13103# vssd1 0.23f $ **FLOATING
C1721 a_8951_13103# vssd1 0.972f $ **FLOATING
C1722 _0503_ vssd1 4.1f $ **FLOATING
C1723 a_8251_13469# vssd1 0.609f $ **FLOATING
C1724 a_8419_13371# vssd1 0.817f $ **FLOATING
C1725 a_7826_13469# vssd1 0.626f $ **FLOATING
C1726 a_7994_13215# vssd1 0.581f $ **FLOATING
C1727 a_7553_13103# vssd1 1.43f $ **FLOATING
C1728 _0019_ vssd1 1.11f $ **FLOATING
C1729 a_7387_13103# vssd1 1.81f $ **FLOATING
C1730 _0018_ vssd1 0.913f $ **FLOATING
C1731 a_4259_13103# vssd1 0.21f $ **FLOATING
C1732 a_5165_13103# vssd1 0.23f $ **FLOATING
C1733 _0860_ vssd1 6.34f $ **FLOATING
C1734 a_6699_13268# vssd1 0.524f $ **FLOATING
C1735 a_5675_13469# vssd1 0.609f $ **FLOATING
C1736 a_5843_13371# vssd1 0.817f $ **FLOATING
C1737 a_5250_13469# vssd1 0.626f $ **FLOATING
C1738 a_5418_13215# vssd1 0.581f $ **FLOATING
C1739 a_4977_13103# vssd1 1.43f $ **FLOATING
C1740 a_4811_13103# vssd1 1.81f $ **FLOATING
C1741 _0204_ vssd1 0.984f $ **FLOATING
C1742 a_3891_13353# vssd1 0.238f $ **FLOATING
C1743 _0389_ vssd1 2.19f $ **FLOATING
C1744 a_4487_13077# vssd1 0.446f $ **FLOATING
C1745 _0397_ vssd1 0.727f $ **FLOATING
C1746 a_2221_13255# vssd1 0.502f $ **FLOATING
C1747 a_28149_14025# vssd1 0.23f $ **FLOATING
C1748 _0360_ vssd1 1.08f $ **FLOATING
C1749 _0015_ vssd1 1.77f $ **FLOATING
C1750 a_20296_13647# vssd1 0.259f $ **FLOATING
C1751 _0013_ vssd1 1f $ **FLOATING
C1752 _0534_ vssd1 0.854f $ **FLOATING
C1753 a_17996_13647# vssd1 0.259f $ **FLOATING
C1754 a_17168_13647# vssd1 0.259f $ **FLOATING
C1755 a_18689_13647# vssd1 0.23f $ **FLOATING
C1756 _0596_ vssd1 1.21f $ **FLOATING
C1757 _0600_ vssd1 0.905f $ **FLOATING
C1758 a_14277_13647# vssd1 0.206f $ **FLOATING
C1759 a_13649_13647# vssd1 0.191f $ **FLOATING
C1760 a_15101_13647# vssd1 0.23f $ **FLOATING
C1761 _0021_ vssd1 1.26f $ **FLOATING
C1762 _0862_ vssd1 1.11f $ **FLOATING
C1763 _0861_ vssd1 1.28f $ **FLOATING
C1764 _0173_ vssd1 1.05f $ **FLOATING
C1765 a_27731_14025# vssd1 0.581f $ **FLOATING
C1766 a_27802_13924# vssd1 0.626f $ **FLOATING
C1767 a_27602_13769# vssd1 1.43f $ **FLOATING
C1768 a_27595_13865# vssd1 1.81f $ **FLOATING
C1769 a_27311_13879# vssd1 0.609f $ **FLOATING
C1770 a_27215_13879# vssd1 0.817f $ **FLOATING
C1771 a_25875_13647# vssd1 0.508f $ **FLOATING
C1772 a_25695_13647# vssd1 0.604f $ **FLOATING
C1773 a_23763_13647# vssd1 0.524f $ **FLOATING
C1774 _0857_ vssd1 0.961f $ **FLOATING
C1775 _0855_ vssd1 1.08f $ **FLOATING
C1776 a_22431_13866# vssd1 0.524f $ **FLOATING
C1777 cal_lut\[174\] vssd1 3.24f $ **FLOATING
C1778 a_21971_13879# vssd1 0.619f $ **FLOATING
C1779 a_20635_13647# vssd1 0.524f $ **FLOATING
C1780 _0530_ vssd1 3.38f $ **FLOATING
C1781 _0533_ vssd1 1.41f $ **FLOATING
C1782 a_19865_13621# vssd1 0.672f $ **FLOATING
C1783 a_19199_13647# vssd1 0.609f $ **FLOATING
C1784 a_19367_13621# vssd1 0.817f $ **FLOATING
C1785 a_18774_13647# vssd1 0.626f $ **FLOATING
C1786 a_18942_13621# vssd1 0.581f $ **FLOATING
C1787 a_18501_13653# vssd1 1.43f $ **FLOATING
C1788 a_18335_13653# vssd1 1.81f $ **FLOATING
C1789 _0593_ vssd1 3.13f $ **FLOATING
C1790 _0594_ vssd1 3.77f $ **FLOATING
C1791 a_17565_13621# vssd1 0.672f $ **FLOATING
C1792 _0597_ vssd1 1.65f $ **FLOATING
C1793 _0598_ vssd1 4.45f $ **FLOATING
C1794 a_16737_13621# vssd1 0.672f $ **FLOATING
C1795 a_15611_13647# vssd1 0.609f $ **FLOATING
C1796 a_15779_13621# vssd1 0.817f $ **FLOATING
C1797 a_15186_13647# vssd1 0.626f $ **FLOATING
C1798 a_15354_13621# vssd1 0.581f $ **FLOATING
C1799 a_14913_13653# vssd1 1.43f $ **FLOATING
C1800 _0010_ vssd1 0.961f $ **FLOATING
C1801 a_14747_13653# vssd1 1.81f $ **FLOATING
C1802 cal_lut\[16\] vssd1 6.18f $ **FLOATING
C1803 _0456_ vssd1 8.06f $ **FLOATING
C1804 a_14131_13879# vssd1 0.804f $ **FLOATING
C1805 _0575_ vssd1 0.627f $ **FLOATING
C1806 _0515_ vssd1 9.26f $ **FLOATING
C1807 a_13512_13621# vssd1 0.847f $ **FLOATING
C1808 a_11987_13647# vssd1 0.524f $ **FLOATING
C1809 _0864_ vssd1 1.05f $ **FLOATING
C1810 a_10501_13879# vssd1 0.502f $ **FLOATING
C1811 a_9131_13647# vssd1 0.508f $ **FLOATING
C1812 cal_lut\[20\] vssd1 1.46f $ **FLOATING
C1813 a_8951_13647# vssd1 0.604f $ **FLOATING
C1814 a_7751_13647# vssd1 0.508f $ **FLOATING
C1815 cal_lut\[19\] vssd1 2.28f $ **FLOATING
C1816 a_7571_13647# vssd1 0.604f $ **FLOATING
C1817 a_4491_13879# vssd1 0.619f $ **FLOATING
C1818 _0808_ vssd1 3.93f $ **FLOATING
C1819 a_2695_14013# vssd1 0.887f $ **FLOATING
C1820 a_1407_13647# vssd1 0.524f $ **FLOATING
C1821 a_27347_14557# vssd1 0.508f $ **FLOATING
C1822 cal_lut\[167\] vssd1 7.69f $ **FLOATING
C1823 a_27167_14557# vssd1 0.604f $ **FLOATING
C1824 a_26677_14191# vssd1 0.23f $ **FLOATING
C1825 cal_lut\[169\] vssd1 3f $ **FLOATING
C1826 cal_lut\[13\] vssd1 2.03f $ **FLOATING
C1827 a_21173_14191# vssd1 0.23f $ **FLOATING
C1828 a_26259_14191# vssd1 0.581f $ **FLOATING
C1829 a_26330_14165# vssd1 0.626f $ **FLOATING
C1830 a_26123_14165# vssd1 1.81f $ **FLOATING
C1831 a_26130_14465# vssd1 1.43f $ **FLOATING
C1832 a_25839_14165# vssd1 0.609f $ **FLOATING
C1833 a_25743_14343# vssd1 0.817f $ **FLOATING
C1834 a_24683_14191# vssd1 0.698f $ **FLOATING
C1835 a_23671_14191# vssd1 0.524f $ **FLOATING
C1836 _0243_ vssd1 0.647f $ **FLOATING
C1837 a_23299_14557# vssd1 0.508f $ **FLOATING
C1838 a_23119_14557# vssd1 0.604f $ **FLOATING
C1839 a_21683_14557# vssd1 0.609f $ **FLOATING
C1840 a_21851_14459# vssd1 0.817f $ **FLOATING
C1841 a_21258_14557# vssd1 0.626f $ **FLOATING
C1842 a_21426_14303# vssd1 0.581f $ **FLOATING
C1843 a_20985_14191# vssd1 1.43f $ **FLOATING
C1844 _0012_ vssd1 1.02f $ **FLOATING
C1845 a_20819_14191# vssd1 1.81f $ **FLOATING
C1846 net35 vssd1 12.1f $ **FLOATING
C1847 _0854_ vssd1 0.891f $ **FLOATING
C1848 _0532_ vssd1 0.854f $ **FLOATING
C1849 cal_lut\[12\] vssd1 1.75f $ **FLOATING
C1850 _0011_ vssd1 1.02f $ **FLOATING
C1851 cal_lut\[11\] vssd1 1.89f $ **FLOATING
C1852 _0595_ vssd1 0.949f $ **FLOATING
C1853 _0852_ vssd1 1.16f $ **FLOATING
C1854 cal_lut\[22\] vssd1 1.97f $ **FLOATING
C1855 cal_lut\[97\] vssd1 4.23f $ **FLOATING
C1856 a_12525_14191# vssd1 0.23f $ **FLOATING
C1857 a_20308_14441# vssd1 0.502f $ **FLOATING
C1858 a_19807_14191# vssd1 0.619f $ **FLOATING
C1859 a_18151_14191# vssd1 0.524f $ **FLOATING
C1860 _0853_ vssd1 0.68f $ **FLOATING
C1861 a_17732_14441# vssd1 0.502f $ **FLOATING
C1862 a_17231_14191# vssd1 0.619f $ **FLOATING
C1863 a_15575_14191# vssd1 0.524f $ **FLOATING
C1864 _0865_ vssd1 0.875f $ **FLOATING
C1865 a_15193_14343# vssd1 0.502f $ **FLOATING
C1866 a_14696_14441# vssd1 0.502f $ **FLOATING
C1867 a_13035_14557# vssd1 0.609f $ **FLOATING
C1868 a_13203_14459# vssd1 0.817f $ **FLOATING
C1869 a_12610_14557# vssd1 0.626f $ **FLOATING
C1870 a_12778_14303# vssd1 0.581f $ **FLOATING
C1871 a_12337_14191# vssd1 1.43f $ **FLOATING
C1872 a_12171_14191# vssd1 1.81f $ **FLOATING
C1873 a_10961_14191# vssd1 0.23f $ **FLOATING
C1874 a_11471_14557# vssd1 0.609f $ **FLOATING
C1875 a_11639_14459# vssd1 0.817f $ **FLOATING
C1876 a_11046_14557# vssd1 0.626f $ **FLOATING
C1877 a_11214_14303# vssd1 0.581f $ **FLOATING
C1878 a_10773_14191# vssd1 1.43f $ **FLOATING
C1879 a_10607_14191# vssd1 1.81f $ **FLOATING
C1880 net30 vssd1 12.2f $ **FLOATING
C1881 cal_lut\[80\] vssd1 1.99f $ **FLOATING
C1882 a_9305_14191# vssd1 0.23f $ **FLOATING
C1883 a_9815_14557# vssd1 0.609f $ **FLOATING
C1884 a_9983_14459# vssd1 0.817f $ **FLOATING
C1885 a_9390_14557# vssd1 0.626f $ **FLOATING
C1886 a_9558_14303# vssd1 0.581f $ **FLOATING
C1887 a_9117_14191# vssd1 1.43f $ **FLOATING
C1888 a_8951_14191# vssd1 1.81f $ **FLOATING
C1889 cal_lut\[37\] vssd1 2.77f $ **FLOATING
C1890 a_7465_14191# vssd1 0.23f $ **FLOATING
C1891 a_7975_14557# vssd1 0.609f $ **FLOATING
C1892 a_8143_14459# vssd1 0.817f $ **FLOATING
C1893 a_7550_14557# vssd1 0.626f $ **FLOATING
C1894 a_7718_14303# vssd1 0.581f $ **FLOATING
C1895 a_7277_14191# vssd1 1.43f $ **FLOATING
C1896 a_7111_14191# vssd1 1.81f $ **FLOATING
C1897 a_3981_14441# vssd1 0.203f $ **FLOATING
C1898 a_2497_14191# vssd1 0.23f $ **FLOATING
C1899 a_5179_14191# vssd1 0.698f $ **FLOATING
C1900 a_3852_14165# vssd1 0.655f $ **FLOATING
C1901 a_3007_14557# vssd1 0.609f $ **FLOATING
C1902 a_3175_14459# vssd1 0.97f $ **FLOATING
C1903 a_2582_14557# vssd1 0.626f $ **FLOATING
C1904 a_2750_14303# vssd1 0.581f $ **FLOATING
C1905 a_2309_14191# vssd1 1.43f $ **FLOATING
C1906 a_2143_14191# vssd1 1.81f $ **FLOATING
C1907 a_1651_14165# vssd1 1.2f $ **FLOATING
C1908 _0168_ vssd1 1.16f $ **FLOATING
C1909 a_23841_14735# vssd1 0.23f $ **FLOATING
C1910 cal_lut\[67\] vssd1 3.08f $ **FLOATING
C1911 a_22277_14735# vssd1 0.23f $ **FLOATING
C1912 _0527_ vssd1 1.23f $ **FLOATING
C1913 _0501_ vssd1 8.29f $ **FLOATING
C1914 a_17033_14735# vssd1 0.23f $ **FLOATING
C1915 net80 vssd1 4.06f $ **FLOATING
C1916 _0096_ vssd1 1.13f $ **FLOATING
C1917 _0080_ vssd1 0.975f $ **FLOATING
C1918 a_8477_14735# vssd1 0.23f $ **FLOATING
C1919 a_6729_14735# vssd1 0.216f $ **FLOATING
C1920 a_3151_14735# vssd1 0.253f $ **FLOATING
C1921 a_5073_14735# vssd1 0.23f $ **FLOATING
C1922 a_4437_15055# vssd1 0.21f $ **FLOATING
C1923 a_27259_14735# vssd1 0.524f $ **FLOATING
C1924 _0353_ vssd1 1f $ **FLOATING
C1925 a_26155_14735# vssd1 0.524f $ **FLOATING
C1926 _0354_ vssd1 0.647f $ **FLOATING
C1927 a_25783_14735# vssd1 0.508f $ **FLOATING
C1928 a_25603_14735# vssd1 0.604f $ **FLOATING
C1929 _0352_ vssd1 9.98f $ **FLOATING
C1930 a_25187_15041# vssd1 0.604f $ **FLOATING
C1931 cal_lut\[68\] vssd1 2.92f $ **FLOATING
C1932 a_25011_14709# vssd1 0.508f $ **FLOATING
C1933 a_24351_14735# vssd1 0.609f $ **FLOATING
C1934 a_24519_14709# vssd1 0.817f $ **FLOATING
C1935 a_23926_14735# vssd1 0.626f $ **FLOATING
C1936 a_24094_14709# vssd1 0.581f $ **FLOATING
C1937 a_23653_14741# vssd1 1.43f $ **FLOATING
C1938 _0067_ vssd1 1.01f $ **FLOATING
C1939 a_23487_14741# vssd1 1.81f $ **FLOATING
C1940 a_22787_14735# vssd1 0.609f $ **FLOATING
C1941 a_22955_14709# vssd1 0.817f $ **FLOATING
C1942 a_22362_14735# vssd1 0.626f $ **FLOATING
C1943 a_22530_14709# vssd1 0.581f $ **FLOATING
C1944 a_22089_14741# vssd1 1.43f $ **FLOATING
C1945 a_21923_14741# vssd1 1.81f $ **FLOATING
C1946 a_20775_14967# vssd1 0.619f $ **FLOATING
C1947 a_19977_14709# vssd1 0.713f $ **FLOATING
C1948 a_17543_14735# vssd1 0.609f $ **FLOATING
C1949 a_17711_14709# vssd1 0.817f $ **FLOATING
C1950 a_17118_14735# vssd1 0.626f $ **FLOATING
C1951 a_17286_14709# vssd1 0.581f $ **FLOATING
C1952 a_16845_14741# vssd1 1.43f $ **FLOATING
C1953 _0022_ vssd1 1.8f $ **FLOATING
C1954 a_16679_14741# vssd1 1.81f $ **FLOATING
C1955 a_16311_14735# vssd1 0.524f $ **FLOATING
C1956 a_14616_14709# vssd1 0.648f $ **FLOATING
C1957 a_12863_14954# vssd1 0.524f $ **FLOATING
C1958 a_12120_14851# vssd1 0.502f $ **FLOATING
C1959 cal_lut\[81\] vssd1 2.06f $ **FLOATING
C1960 a_11207_14954# vssd1 0.524f $ **FLOATING
C1961 a_10699_14735# vssd1 0.524f $ **FLOATING
C1962 _0257_ vssd1 1.24f $ **FLOATING
C1963 a_9823_15041# vssd1 0.604f $ **FLOATING
C1964 cal_lut\[79\] vssd1 2.09f $ **FLOATING
C1965 a_9647_14709# vssd1 0.508f $ **FLOATING
C1966 a_8987_14735# vssd1 0.609f $ **FLOATING
C1967 a_9155_14709# vssd1 0.817f $ **FLOATING
C1968 a_8562_14735# vssd1 0.626f $ **FLOATING
C1969 a_8730_14709# vssd1 0.581f $ **FLOATING
C1970 a_8289_14741# vssd1 1.43f $ **FLOATING
C1971 a_8123_14741# vssd1 1.81f $ **FLOATING
C1972 net28 vssd1 5.21f $ **FLOATING
C1973 a_7239_14735# vssd1 0.599f $ **FLOATING
C1974 a_7410_14709# vssd1 1.41f $ **FLOATING
C1975 a_6823_14735# vssd1 0.627f $ **FLOATING
C1976 a_6982_14709# vssd1 0.587f $ **FLOATING
C1977 a_6541_14741# vssd1 1.39f $ **FLOATING
C1978 a_6375_14741# vssd1 1.77f $ **FLOATING
C1979 a_5583_14735# vssd1 0.609f $ **FLOATING
C1980 a_5751_14709# vssd1 0.97f $ **FLOATING
C1981 a_5158_14735# vssd1 0.626f $ **FLOATING
C1982 a_5326_14709# vssd1 0.581f $ **FLOATING
C1983 a_4885_14741# vssd1 1.43f $ **FLOATING
C1984 _0205_ vssd1 1.01f $ **FLOATING
C1985 a_4719_14741# vssd1 1.81f $ **FLOATING
C1986 _0398_ vssd1 1.07f $ **FLOATING
C1987 a_4245_14796# vssd1 0.446f $ **FLOATING
C1988 _0202_ vssd1 1.19f $ **FLOATING
C1989 ctr\[0\] vssd1 1.9f $ **FLOATING
C1990 a_1761_14735# vssd1 0.23f $ **FLOATING
C1991 _0394_ vssd1 1f $ **FLOATING
C1992 _0393_ vssd1 1.2f $ **FLOATING
C1993 a_2933_14709# vssd1 0.55f $ **FLOATING
C1994 a_2271_14735# vssd1 0.609f $ **FLOATING
C1995 a_2439_14709# vssd1 0.817f $ **FLOATING
C1996 a_1846_14735# vssd1 0.626f $ **FLOATING
C1997 a_2014_14709# vssd1 0.581f $ **FLOATING
C1998 a_1573_14741# vssd1 1.43f $ **FLOATING
C1999 a_1407_14741# vssd1 1.81f $ **FLOATING
C2000 a_28057_15279# vssd1 0.23f $ **FLOATING
C2001 _0167_ vssd1 1.23f $ **FLOATING
C2002 a_27639_15279# vssd1 0.581f $ **FLOATING
C2003 a_27710_15253# vssd1 0.626f $ **FLOATING
C2004 a_27503_15253# vssd1 1.81f $ **FLOATING
C2005 a_27510_15553# vssd1 1.43f $ **FLOATING
C2006 a_27219_15253# vssd1 0.609f $ **FLOATING
C2007 a_27123_15431# vssd1 0.817f $ **FLOATING
C2008 _0244_ vssd1 0.81f $ **FLOATING
C2009 a_24823_15444# vssd1 0.524f $ **FLOATING
C2010 a_24407_15279# vssd1 0.648f $ **FLOATING
C2011 _0656_ vssd1 3.26f $ **FLOATING
C2012 _0537_ vssd1 2.89f $ **FLOATING
C2013 net37 vssd1 8.38f $ **FLOATING
C2014 _0066_ vssd1 1.26f $ **FLOATING
C2015 a_19609_15279# vssd1 0.23f $ **FLOATING
C2016 a_23811_15431# vssd1 0.619f $ **FLOATING
C2017 a_22983_15431# vssd1 0.619f $ **FLOATING
C2018 a_22619_15253# vssd1 0.698f $ **FLOATING
C2019 a_21739_15279# vssd1 0.524f $ **FLOATING
C2020 _0242_ vssd1 0.719f $ **FLOATING
C2021 a_21228_15529# vssd1 0.502f $ **FLOATING
C2022 a_20779_15253# vssd1 0.698f $ **FLOATING
C2023 a_20119_15645# vssd1 0.609f $ **FLOATING
C2024 a_20287_15547# vssd1 0.817f $ **FLOATING
C2025 a_19694_15645# vssd1 0.626f $ **FLOATING
C2026 a_19862_15391# vssd1 0.581f $ **FLOATING
C2027 a_19421_15279# vssd1 1.43f $ **FLOATING
C2028 a_19255_15279# vssd1 1.81f $ **FLOATING
C2029 net38 vssd1 12.5f $ **FLOATING
C2030 _0023_ vssd1 1.03f $ **FLOATING
C2031 cal_lut\[23\] vssd1 1.84f $ **FLOATING
C2032 a_17812_15529# vssd1 0.259f $ **FLOATING
C2033 _0599_ vssd1 1.58f $ **FLOATING
C2034 _0549_ vssd1 2.8f $ **FLOATING
C2035 _0275_ vssd1 0.863f $ **FLOATING
C2036 a_11421_15279# vssd1 0.23f $ **FLOATING
C2037 a_18611_15279# vssd1 0.524f $ **FLOATING
C2038 _0866_ vssd1 0.68f $ **FLOATING
C2039 a_18192_15529# vssd1 0.502f $ **FLOATING
C2040 a_17381_15425# vssd1 0.672f $ **FLOATING
C2041 a_16035_15279# vssd1 0.619f $ **FLOATING
C2042 a_15623_15431# vssd1 0.619f $ **FLOATING
C2043 a_15193_15431# vssd1 0.502f $ **FLOATING
C2044 a_14733_15431# vssd1 0.502f $ **FLOATING
C2045 a_14273_15431# vssd1 0.502f $ **FLOATING
C2046 a_13537_15431# vssd1 0.502f $ **FLOATING
C2047 a_13135_15253# vssd1 0.604f $ **FLOATING
C2048 a_12959_15253# vssd1 0.508f $ **FLOATING
C2049 a_11931_15645# vssd1 0.609f $ **FLOATING
C2050 a_12099_15547# vssd1 0.817f $ **FLOATING
C2051 a_11506_15645# vssd1 0.626f $ **FLOATING
C2052 a_11674_15391# vssd1 0.581f $ **FLOATING
C2053 a_11233_15279# vssd1 1.43f $ **FLOATING
C2054 _0004_ vssd1 0.977f $ **FLOATING
C2055 a_11067_15279# vssd1 1.81f $ **FLOATING
C2056 net29 vssd1 13.2f $ **FLOATING
C2057 _0079_ vssd1 1.19f $ **FLOATING
C2058 _0078_ vssd1 1f $ **FLOATING
C2059 _0036_ vssd1 1.23f $ **FLOATING
C2060 net77 vssd1 1.5f $ **FLOATING
C2061 _0810_ vssd1 1.14f $ **FLOATING
C2062 _0809_ vssd1 2.66f $ **FLOATING
C2063 a_4091_15529# vssd1 0.224f $ **FLOATING
C2064 _0199_ vssd1 0.967f $ **FLOATING
C2065 _0661_ vssd1 2.44f $ **FLOATING
C2066 a_10839_15444# vssd1 0.524f $ **FLOATING
C2067 a_9595_15279# vssd1 0.524f $ **FLOATING
C2068 _0256_ vssd1 0.895f $ **FLOATING
C2069 a_9275_15444# vssd1 0.524f $ **FLOATING
C2070 _0255_ vssd1 2.85f $ **FLOATING
C2071 a_8263_15444# vssd1 0.524f $ **FLOATING
C2072 _0880_ vssd1 3.72f $ **FLOATING
C2073 a_7527_15444# vssd1 0.524f $ **FLOATING
C2074 a_5971_15253# vssd1 0.788f $ **FLOATING
C2075 a_5713_15253# vssd1 0.794f $ **FLOATING
C2076 a_5617_15431# vssd1 0.553f $ **FLOATING
C2077 a_4843_15307# vssd1 0.56f $ **FLOATING
C2078 net68 vssd1 0.874f $ **FLOATING
C2079 a_3851_15253# vssd1 1.12f $ **FLOATING
C2080 clknet_1_0__leaf_net67 vssd1 6.71f $ **FLOATING
C2081 a_1945_15431# vssd1 0.502f $ **FLOATING
C2082 _0388_ vssd1 0.68f $ **FLOATING
C2083 a_1639_15444# vssd1 0.524f $ **FLOATING
C2084 a_27521_15823# vssd1 0.23f $ **FLOATING
C2085 a_24853_15823# vssd1 0.23f $ **FLOATING
C2086 _0551_ vssd1 2.53f $ **FLOATING
C2087 a_18029_16201# vssd1 0.23f $ **FLOATING
C2088 a_16156_15823# vssd1 0.259f $ **FLOATING
C2089 cal_lut\[78\] vssd1 3.53f $ **FLOATING
C2090 cal_lut\[36\] vssd1 1.81f $ **FLOATING
C2091 a_13997_15823# vssd1 0.23f $ **FLOATING
C2092 _0844_ vssd1 1.26f $ **FLOATING
C2093 a_9949_15823# vssd1 0.23f $ **FLOATING
C2094 a_8293_15823# vssd1 0.23f $ **FLOATING
C2095 a_5825_15823# vssd1 0.325f $ **FLOATING
C2096 a_5460_15823# vssd1 0.429f $ **FLOATING
C2097 a_4624_15823# vssd1 0.237f $ **FLOATING
C2098 _0192_ vssd1 1.57f $ **FLOATING
C2099 a_5377_16143# vssd1 0.267f $ **FLOATING
C2100 _0387_ vssd1 0.918f $ **FLOATING
C2101 a_2313_15823# vssd1 0.23f $ **FLOATING
C2102 a_28031_15823# vssd1 0.609f $ **FLOATING
C2103 a_28199_15797# vssd1 0.817f $ **FLOATING
C2104 a_27606_15823# vssd1 0.626f $ **FLOATING
C2105 a_27774_15797# vssd1 0.581f $ **FLOATING
C2106 a_27333_15829# vssd1 1.43f $ **FLOATING
C2107 a_27167_15829# vssd1 1.81f $ **FLOATING
C2108 _0249_ vssd1 0.758f $ **FLOATING
C2109 a_26479_16042# vssd1 0.524f $ **FLOATING
C2110 a_26012_15939# vssd1 0.502f $ **FLOATING
C2111 cal_lut\[72\] vssd1 3.56f $ **FLOATING
C2112 a_25363_15823# vssd1 0.609f $ **FLOATING
C2113 a_25531_15797# vssd1 0.817f $ **FLOATING
C2114 a_24938_15823# vssd1 0.626f $ **FLOATING
C2115 a_25106_15797# vssd1 0.581f $ **FLOATING
C2116 a_24665_15829# vssd1 1.43f $ **FLOATING
C2117 _0068_ vssd1 0.961f $ **FLOATING
C2118 a_24499_15829# vssd1 1.81f $ **FLOATING
C2119 _0505_ vssd1 16.9f $ **FLOATING
C2120 cal_lut\[168\] vssd1 4.08f $ **FLOATING
C2121 a_21879_16055# vssd1 0.619f $ **FLOATING
C2122 _0850_ vssd1 23.1f $ **FLOATING
C2123 a_20963_15797# vssd1 0.698f $ **FLOATING
C2124 a_20400_15939# vssd1 0.502f $ **FLOATING
C2125 cal_lut\[24\] vssd1 2f $ **FLOATING
C2126 a_17611_16201# vssd1 0.581f $ **FLOATING
C2127 a_17682_16100# vssd1 0.626f $ **FLOATING
C2128 a_17482_15945# vssd1 1.43f $ **FLOATING
C2129 a_17475_16041# vssd1 1.81f $ **FLOATING
C2130 a_17191_16055# vssd1 0.609f $ **FLOATING
C2131 a_17095_16055# vssd1 0.817f $ **FLOATING
C2132 _0541_ vssd1 6.5f $ **FLOATING
C2133 _0542_ vssd1 4.54f $ **FLOATING
C2134 a_15725_15797# vssd1 0.672f $ **FLOATING
C2135 _0543_ vssd1 0.636f $ **FLOATING
C2136 _0546_ vssd1 4.09f $ **FLOATING
C2137 _0550_ vssd1 2.98f $ **FLOATING
C2138 _0554_ vssd1 1.75f $ **FLOATING
C2139 a_14507_15823# vssd1 0.609f $ **FLOATING
C2140 a_14675_15797# vssd1 0.817f $ **FLOATING
C2141 a_14082_15823# vssd1 0.626f $ **FLOATING
C2142 a_14250_15797# vssd1 0.581f $ **FLOATING
C2143 a_13809_15829# vssd1 1.43f $ **FLOATING
C2144 a_13643_15829# vssd1 1.81f $ **FLOATING
C2145 _0518_ vssd1 1.74f $ **FLOATING
C2146 a_13052_15797# vssd1 0.648f $ **FLOATING
C2147 a_11605_16055# vssd1 0.502f $ **FLOATING
C2148 a_10459_15823# vssd1 0.609f $ **FLOATING
C2149 a_10627_15797# vssd1 0.817f $ **FLOATING
C2150 a_10034_15823# vssd1 0.626f $ **FLOATING
C2151 a_10202_15797# vssd1 0.581f $ **FLOATING
C2152 a_9761_15829# vssd1 1.43f $ **FLOATING
C2153 _0003_ vssd1 1.01f $ **FLOATING
C2154 a_9595_15829# vssd1 1.81f $ **FLOATING
C2155 a_8803_15823# vssd1 0.609f $ **FLOATING
C2156 a_8971_15797# vssd1 0.817f $ **FLOATING
C2157 a_8378_15823# vssd1 0.626f $ **FLOATING
C2158 a_8546_15797# vssd1 0.581f $ **FLOATING
C2159 a_8105_15829# vssd1 1.43f $ **FLOATING
C2160 a_7939_15829# vssd1 1.81f $ **FLOATING
C2161 a_7387_15823# vssd1 0.524f $ **FLOATING
C2162 _0840_ vssd1 0.803f $ **FLOATING
C2163 a_7072_15797# vssd1 0.648f $ **FLOATING
C2164 a_6647_15823# vssd1 0.508f $ **FLOATING
C2165 a_6467_15823# vssd1 0.604f $ **FLOATING
C2166 a_4351_15823# vssd1 0.569f $ **FLOATING
C2167 temp_delay_last vssd1 1.61f $ **FLOATING
C2168 a_4027_16144# vssd1 0.604f $ **FLOATING
C2169 a_3575_15797# vssd1 0.85f $ **FLOATING
C2170 a_2823_15823# vssd1 0.609f $ **FLOATING
C2171 a_2991_15797# vssd1 0.817f $ **FLOATING
C2172 a_2398_15823# vssd1 0.626f $ **FLOATING
C2173 a_2566_15797# vssd1 0.581f $ **FLOATING
C2174 a_2125_15829# vssd1 1.43f $ **FLOATING
C2175 _0198_ vssd1 1.68f $ **FLOATING
C2176 a_1959_15829# vssd1 1.81f $ **FLOATING
C2177 a_1407_15823# vssd1 0.698f $ **FLOATING
C2178 _0071_ vssd1 0.96f $ **FLOATING
C2179 a_26233_16367# vssd1 0.23f $ **FLOATING
C2180 a_27351_16367# vssd1 0.524f $ **FLOATING
C2181 a_26743_16733# vssd1 0.609f $ **FLOATING
C2182 a_26911_16635# vssd1 0.817f $ **FLOATING
C2183 a_26318_16733# vssd1 0.626f $ **FLOATING
C2184 a_26486_16479# vssd1 0.581f $ **FLOATING
C2185 a_26045_16367# vssd1 1.43f $ **FLOATING
C2186 _0072_ vssd1 1.03f $ **FLOATING
C2187 a_25879_16367# vssd1 1.81f $ **FLOATING
C2188 a_23223_16617# vssd1 0.167f $ **FLOATING
C2189 a_23021_16617# vssd1 0.214f $ **FLOATING
C2190 a_21725_16367# vssd1 0.23f $ **FLOATING
C2191 a_25047_16733# vssd1 0.508f $ **FLOATING
C2192 cal_lut\[69\] vssd1 2.66f $ **FLOATING
C2193 a_24867_16733# vssd1 0.604f $ **FLOATING
C2194 a_23759_16733# vssd1 0.508f $ **FLOATING
C2195 a_23579_16733# vssd1 0.604f $ **FLOATING
C2196 _0688_ vssd1 5.83f $ **FLOATING
C2197 cal_lut\[25\] vssd1 1.71f $ **FLOATING
C2198 a_22895_16519# vssd1 0.972f $ **FLOATING
C2199 a_22235_16733# vssd1 0.609f $ **FLOATING
C2200 a_22403_16635# vssd1 0.817f $ **FLOATING
C2201 a_21810_16733# vssd1 0.626f $ **FLOATING
C2202 a_21978_16479# vssd1 0.581f $ **FLOATING
C2203 a_21537_16367# vssd1 1.43f $ **FLOATING
C2204 a_21371_16367# vssd1 1.81f $ **FLOATING
C2205 _0024_ vssd1 0.872f $ **FLOATING
C2206 _0540_ vssd1 2.78f $ **FLOATING
C2207 _0606_ vssd1 2.9f $ **FLOATING
C2208 _0077_ vssd1 1.31f $ **FLOATING
C2209 a_11895_16367# vssd1 0.554f $ **FLOATING
C2210 a_11439_16367# vssd1 0.275f $ **FLOATING
C2211 a_21095_16367# vssd1 0.524f $ **FLOATING
C2212 _0867_ vssd1 1.04f $ **FLOATING
C2213 a_20407_16519# vssd1 0.619f $ **FLOATING
C2214 a_19756_16617# vssd1 0.502f $ **FLOATING
C2215 a_19303_16519# vssd1 0.619f $ **FLOATING
C2216 a_18611_16367# vssd1 0.524f $ **FLOATING
C2217 a_18291_16532# vssd1 0.524f $ **FLOATING
C2218 a_17875_16367# vssd1 0.648f $ **FLOATING
C2219 _0254_ vssd1 0.945f $ **FLOATING
C2220 _0624_ vssd1 3f $ **FLOATING
C2221 _0617_ vssd1 5.29f $ **FLOATING
C2222 a_9595_16367# vssd1 0.275f $ **FLOATING
C2223 _0035_ vssd1 1.04f $ **FLOATING
C2224 a_12343_16617# vssd1 0.381f $ **FLOATING
C2225 a_11895_16617# vssd1 0.381f $ **FLOATING
C2226 cal_lut\[4\] vssd1 1.41f $ **FLOATING
C2227 _0843_ vssd1 1.1f $ **FLOATING
C2228 a_7741_16367# vssd1 0.23f $ **FLOATING
C2229 a_17456_16617# vssd1 0.502f $ **FLOATING
C2230 a_16373_16341# vssd1 0.858f $ **FLOATING
C2231 _0879_ vssd1 1.21f $ **FLOATING
C2232 a_14243_16532# vssd1 0.524f $ **FLOATING
C2233 a_12856_16617# vssd1 0.502f $ **FLOATING
C2234 cal_lut\[5\] vssd1 2.37f $ **FLOATING
C2235 _0625_ vssd1 3.18f $ **FLOATING
C2236 _0609_ vssd1 4.59f $ **FLOATING
C2237 a_11302_16519# vssd1 0.597f $ **FLOATING
C2238 a_10832_16617# vssd1 0.502f $ **FLOATING
C2239 a_9749_16617# vssd1 0.597f $ **FLOATING
C2240 _0702_ vssd1 3.36f $ **FLOATING
C2241 cal_lut\[1\] vssd1 5.59f $ **FLOATING
C2242 a_9223_16733# vssd1 0.508f $ **FLOATING
C2243 a_9043_16733# vssd1 0.604f $ **FLOATING
C2244 a_8251_16733# vssd1 0.609f $ **FLOATING
C2245 a_8419_16635# vssd1 0.817f $ **FLOATING
C2246 a_7826_16733# vssd1 0.626f $ **FLOATING
C2247 a_7994_16479# vssd1 0.581f $ **FLOATING
C2248 a_7553_16367# vssd1 1.43f $ **FLOATING
C2249 _0001_ vssd1 0.954f $ **FLOATING
C2250 a_7387_16367# vssd1 1.81f $ **FLOATING
C2251 a_4733_16367# vssd1 0.267f $ **FLOATING
C2252 a_5993_16367# vssd1 0.216f $ **FLOATING
C2253 a_6503_16733# vssd1 0.599f $ **FLOATING
C2254 a_6674_16620# vssd1 1.41f $ **FLOATING
C2255 a_6087_16733# vssd1 0.627f $ **FLOATING
C2256 a_6246_16503# vssd1 0.587f $ **FLOATING
C2257 a_5805_16367# vssd1 1.39f $ **FLOATING
C2258 a_5639_16367# vssd1 1.77f $ **FLOATING
C2259 _0193_ vssd1 1.08f $ **FLOATING
C2260 a_5181_16617# vssd1 0.325f $ **FLOATING
C2261 a_4816_16617# vssd1 0.429f $ **FLOATING
C2262 net69 vssd1 1.1f $ **FLOATING
C2263 a_4167_16367# vssd1 1.2f $ **FLOATING
C2264 a_24469_17289# vssd1 0.23f $ **FLOATING
C2265 _0250_ vssd1 0.758f $ **FLOATING
C2266 a_27491_17130# vssd1 0.524f $ **FLOATING
C2267 a_27024_17027# vssd1 0.502f $ **FLOATING
C2268 cal_lut\[73\] vssd1 2.97f $ **FLOATING
C2269 a_25327_16911# vssd1 0.524f $ **FLOATING
C2270 _0245_ vssd1 1.08f $ **FLOATING
C2271 a_24051_17289# vssd1 0.581f $ **FLOATING
C2272 a_24122_17188# vssd1 0.626f $ **FLOATING
C2273 a_23922_17033# vssd1 1.43f $ **FLOATING
C2274 a_23915_17129# vssd1 1.81f $ **FLOATING
C2275 a_23631_17143# vssd1 0.609f $ **FLOATING
C2276 a_23535_17143# vssd1 0.817f $ **FLOATING
C2277 a_22875_17249# vssd1 0.56f $ **FLOATING
C2278 _0689_ vssd1 1.12f $ **FLOATING
C2279 _0684_ vssd1 3.44f $ **FLOATING
C2280 _0692_ vssd1 6.02f $ **FLOATING
C2281 a_20345_16911# vssd1 0.23f $ **FLOATING
C2282 cal_lut\[29\] vssd1 1.46f $ **FLOATING
C2283 a_18873_16911# vssd1 0.23f $ **FLOATING
C2284 _0871_ vssd1 1.07f $ **FLOATING
C2285 _0477_ vssd1 16.2f $ **FLOATING
C2286 _0455_ vssd1 2.84f $ **FLOATING
C2287 _0002_ vssd1 1.32f $ **FLOATING
C2288 a_6391_16911# vssd1 0.388f $ **FLOATING
C2289 a_5639_16911# vssd1 0.388f $ **FLOATING
C2290 _0382_ vssd1 1.64f $ **FLOATING
C2291 _0381_ vssd1 1.37f $ **FLOATING
C2292 a_21878_17143# vssd1 0.702f $ **FLOATING
C2293 a_20855_16911# vssd1 0.609f $ **FLOATING
C2294 a_21023_16885# vssd1 0.817f $ **FLOATING
C2295 a_20430_16911# vssd1 0.626f $ **FLOATING
C2296 a_20598_16885# vssd1 0.581f $ **FLOATING
C2297 a_20157_16917# vssd1 1.43f $ **FLOATING
C2298 a_19991_16917# vssd1 1.81f $ **FLOATING
C2299 a_19383_16911# vssd1 0.609f $ **FLOATING
C2300 a_19551_16885# vssd1 0.817f $ **FLOATING
C2301 a_18958_16911# vssd1 0.626f $ **FLOATING
C2302 a_19126_16885# vssd1 0.581f $ **FLOATING
C2303 a_18685_16917# vssd1 1.43f $ **FLOATING
C2304 _0028_ vssd1 0.961f $ **FLOATING
C2305 a_18519_16917# vssd1 1.81f $ **FLOATING
C2306 a_18100_17027# vssd1 0.502f $ **FLOATING
C2307 _0851_ vssd1 12.3f $ **FLOATING
C2308 a_15439_17130# vssd1 0.524f $ **FLOATING
C2309 a_14523_16885# vssd1 0.698f $ **FLOATING
C2310 a_13751_16911# vssd1 0.795f $ **FLOATING
C2311 a_13968_17218# vssd1 0.788f $ **FLOATING
C2312 a_13551_16911# vssd1 0.696f $ **FLOATING
C2313 a_12950_16988# vssd1 0.658f $ **FLOATING
C2314 _0845_ vssd1 1.27f $ **FLOATING
C2315 a_12219_17130# vssd1 0.524f $ **FLOATING
C2316 _0842_ vssd1 0.725f $ **FLOATING
C2317 a_8723_17130# vssd1 0.524f $ **FLOATING
C2318 a_8303_16911# vssd1 0.508f $ **FLOATING
C2319 a_8123_16911# vssd1 0.604f $ **FLOATING
C2320 a_7631_17171# vssd1 1.2f $ **FLOATING
C2321 a_6927_16911# vssd1 0.698f $ **FLOATING
C2322 net2 vssd1 8.31f $ **FLOATING
C2323 a_3882_16911# vssd1 4.03f $ **FLOATING
C2324 net67 vssd1 5.4f $ **FLOATING
C2325 a_3155_16911# vssd1 1.2f $ **FLOATING
C2326 a_2879_16911# vssd1 0.524f $ **FLOATING
C2327 _0379_ vssd1 1.44f $ **FLOATING
C2328 a_2417_17027# vssd1 0.601f $ **FLOATING
C2329 a_2317_16911# vssd1 0.488f $ **FLOATING
C2330 a_1773_17027# vssd1 0.601f $ **FLOATING
C2331 a_1673_16911# vssd1 0.488f $ **FLOATING
C2332 a_27521_17455# vssd1 0.23f $ **FLOATING
C2333 a_28031_17821# vssd1 0.609f $ **FLOATING
C2334 a_28199_17723# vssd1 0.817f $ **FLOATING
C2335 a_27606_17821# vssd1 0.626f $ **FLOATING
C2336 a_27774_17567# vssd1 0.581f $ **FLOATING
C2337 a_27333_17455# vssd1 1.43f $ **FLOATING
C2338 _0073_ vssd1 0.908f $ **FLOATING
C2339 a_27167_17455# vssd1 1.81f $ **FLOATING
C2340 _0248_ vssd1 1.24f $ **FLOATING
C2341 a_25589_17455# vssd1 0.23f $ **FLOATING
C2342 a_26748_17705# vssd1 0.502f $ **FLOATING
C2343 a_26099_17821# vssd1 0.609f $ **FLOATING
C2344 a_26267_17723# vssd1 0.817f $ **FLOATING
C2345 a_25674_17821# vssd1 0.626f $ **FLOATING
C2346 a_25842_17567# vssd1 0.581f $ **FLOATING
C2347 a_25401_17455# vssd1 1.43f $ **FLOATING
C2348 _0069_ vssd1 0.908f $ **FLOATING
C2349 a_25235_17455# vssd1 1.81f $ **FLOATING
C2350 _0025_ vssd1 1.3f $ **FLOATING
C2351 a_23407_17705# vssd1 0.167f $ **FLOATING
C2352 a_23205_17705# vssd1 0.214f $ **FLOATING
C2353 a_24485_17607# vssd1 0.502f $ **FLOATING
C2354 a_23763_17455# vssd1 0.524f $ **FLOATING
C2355 _0868_ vssd1 1.15f $ **FLOATING
C2356 _0479_ vssd1 6.08f $ **FLOATING
C2357 cal_lut\[74\] vssd1 3.18f $ **FLOATING
C2358 _0473_ vssd1 1.45f $ **FLOATING
C2359 a_23079_17607# vssd1 0.972f $ **FLOATING
C2360 a_21371_17455# vssd1 0.648f $ **FLOATING
C2361 _0029_ vssd1 0.985f $ **FLOATING
C2362 _0613_ vssd1 1.26f $ **FLOATING
C2363 a_16404_17705# vssd1 0.259f $ **FLOATING
C2364 cal_lut\[96\] vssd1 3.4f $ **FLOATING
C2365 a_15285_17455# vssd1 0.23f $ **FLOATING
C2366 a_19991_17455# vssd1 0.524f $ **FLOATING
C2367 _0873_ vssd1 1.13f $ **FLOATING
C2368 a_19303_17607# vssd1 0.619f $ **FLOATING
C2369 a_16574_17455# vssd1 0.672f $ **FLOATING
C2370 _0610_ vssd1 1.71f $ **FLOATING
C2371 cal_lut\[101\] vssd1 4.4f $ **FLOATING
C2372 a_15795_17821# vssd1 0.609f $ **FLOATING
C2373 a_15963_17723# vssd1 0.817f $ **FLOATING
C2374 a_15370_17821# vssd1 0.626f $ **FLOATING
C2375 a_15538_17567# vssd1 0.581f $ **FLOATING
C2376 a_15097_17455# vssd1 1.43f $ **FLOATING
C2377 _0095_ vssd1 0.994f $ **FLOATING
C2378 a_14931_17455# vssd1 1.81f $ **FLOATING
C2379 a_10423_17455# vssd1 0.171f $ **FLOATING
C2380 a_10055_17455# vssd1 0.18f $ **FLOATING
C2381 a_9687_17455# vssd1 0.18f $ **FLOATING
C2382 a_12249_17455# vssd1 0.23f $ **FLOATING
C2383 _0555_ vssd1 1.65f $ **FLOATING
C2384 a_14705_17620# vssd1 0.524f $ **FLOATING
C2385 a_14103_17455# vssd1 1.2f $ **FLOATING
C2386 a_13459_17455# vssd1 1.2f $ **FLOATING
C2387 a_12759_17821# vssd1 0.609f $ **FLOATING
C2388 a_12927_17723# vssd1 0.817f $ **FLOATING
C2389 a_12334_17821# vssd1 0.626f $ **FLOATING
C2390 a_12502_17567# vssd1 0.581f $ **FLOATING
C2391 a_12061_17455# vssd1 1.43f $ **FLOATING
C2392 _0005_ vssd1 0.908f $ **FLOATING
C2393 a_11895_17455# vssd1 1.81f $ **FLOATING
C2394 a_11199_17607# vssd1 0.478f $ **FLOATING
C2395 a_11029_17429# vssd1 0.485f $ **FLOATING
C2396 a_10596_17705# vssd1 0.546f $ **FLOATING
C2397 _0663_ vssd1 1.12f $ **FLOATING
C2398 _0662_ vssd1 1.24f $ **FLOATING
C2399 net12 vssd1 2f $ **FLOATING
C2400 cal_lut\[3\] vssd1 1.84f $ **FLOATING
C2401 a_2931_17455# vssd1 0.45f $ **FLOATING
C2402 a_2489_17455# vssd1 0.361f $ **FLOATING
C2403 a_4811_17705# vssd1 0.388f $ **FLOATING
C2404 a_4531_17705# vssd1 0.253f $ **FLOATING
C2405 a_8544_17429# vssd1 0.648f $ **FLOATING
C2406 a_7111_17455# vssd1 0.698f $ **FLOATING
C2407 a_5341_17429# vssd1 4.03f $ **FLOATING
C2408 _0476_ vssd1 24.1f $ **FLOATING
C2409 a_4313_17429# vssd1 0.55f $ **FLOATING
C2410 a_3891_17455# vssd1 0.648f $ **FLOATING
C2411 _0754_ vssd1 1.38f $ **FLOATING
C2412 _0436_ vssd1 2.85f $ **FLOATING
C2413 net6 vssd1 4.12f $ **FLOATING
C2414 a_1683_17455# vssd1 0.619f $ **FLOATING
C2415 cal_lut\[71\] vssd1 5.09f $ **FLOATING
C2416 a_27337_17999# vssd1 0.23f $ **FLOATING
C2417 a_23056_17999# vssd1 0.259f $ **FLOATING
C2418 a_24945_17999# vssd1 0.23f $ **FLOATING
C2419 a_27847_17999# vssd1 0.609f $ **FLOATING
C2420 a_28015_17973# vssd1 0.817f $ **FLOATING
C2421 a_27422_17999# vssd1 0.626f $ **FLOATING
C2422 a_27590_17973# vssd1 0.581f $ **FLOATING
C2423 a_27149_18005# vssd1 1.43f $ **FLOATING
C2424 _0070_ vssd1 1.15f $ **FLOATING
C2425 a_26983_18005# vssd1 1.81f $ **FLOATING
C2426 a_26417_18231# vssd1 0.502f $ **FLOATING
C2427 a_26063_17999# vssd1 0.524f $ **FLOATING
C2428 _0247_ vssd1 0.758f $ **FLOATING
C2429 a_25455_17999# vssd1 0.609f $ **FLOATING
C2430 a_25623_17973# vssd1 0.817f $ **FLOATING
C2431 a_25030_17999# vssd1 0.626f $ **FLOATING
C2432 a_25198_17973# vssd1 0.581f $ **FLOATING
C2433 a_24757_18005# vssd1 1.43f $ **FLOATING
C2434 _0074_ vssd1 0.872f $ **FLOATING
C2435 a_24591_18005# vssd1 1.81f $ **FLOATING
C2436 a_24315_17999# vssd1 0.524f $ **FLOATING
C2437 _0251_ vssd1 0.947f $ **FLOATING
C2438 _0640_ vssd1 4.92f $ **FLOATING
C2439 _0641_ vssd1 4.43f $ **FLOATING
C2440 a_22625_17973# vssd1 0.672f $ **FLOATING
C2441 _0480_ vssd1 1.16f $ **FLOATING
C2442 _0458_ vssd1 3.86f $ **FLOATING
C2443 _0526_ vssd1 3.24f $ **FLOATING
C2444 _0508_ vssd1 14f $ **FLOATING
C2445 _0475_ vssd1 7.33f $ **FLOATING
C2446 cal_lut\[77\] vssd1 3.06f $ **FLOATING
C2447 a_17217_17999# vssd1 0.23f $ **FLOATING
C2448 _0611_ vssd1 0.964f $ **FLOATING
C2449 _0274_ vssd1 1.49f $ **FLOATING
C2450 a_21970_18231# vssd1 0.702f $ **FLOATING
C2451 a_20775_18231# vssd1 0.619f $ **FLOATING
C2452 a_19308_17973# vssd1 0.648f $ **FLOATING
C2453 a_18369_18337# vssd1 0.713f $ **FLOATING
C2454 a_17727_17999# vssd1 0.609f $ **FLOATING
C2455 a_17895_17973# vssd1 0.817f $ **FLOATING
C2456 a_17302_17999# vssd1 0.626f $ **FLOATING
C2457 a_17470_17973# vssd1 0.581f $ **FLOATING
C2458 a_17029_18005# vssd1 1.43f $ **FLOATING
C2459 a_16863_18005# vssd1 1.81f $ **FLOATING
C2460 a_16035_18112# vssd1 0.619f $ **FLOATING
C2461 a_15561_18231# vssd1 0.502f $ **FLOATING
C2462 a_14655_18115# vssd1 0.858f $ **FLOATING
C2463 a_11950_18319# vssd1 0.2f $ **FLOATING
C2464 a_9135_18319# vssd1 0.18f $ **FLOATING
C2465 a_8491_18319# vssd1 0.275f $ **FLOATING
C2466 a_5825_17999# vssd1 0.325f $ **FLOATING
C2467 a_5460_17999# vssd1 0.429f $ **FLOATING
C2468 a_4143_17999# vssd1 0.495f $ **FLOATING
C2469 a_3785_17999# vssd1 0.422f $ **FLOATING
C2470 a_6729_17999# vssd1 0.216f $ **FLOATING
C2471 a_5377_18319# vssd1 0.267f $ **FLOATING
C2472 a_14287_17999# vssd1 0.698f $ **FLOATING
C2473 _0539_ vssd1 5.69f $ **FLOATING
C2474 a_13969_18218# vssd1 0.524f $ **FLOATING
C2475 _0836_ vssd1 13.5f $ **FLOATING
C2476 a_12525_18231# vssd1 0.502f $ **FLOATING
C2477 _0588_ vssd1 1.71f $ **FLOATING
C2478 _0576_ vssd1 3.02f $ **FLOATING
C2479 _0574_ vssd1 5f $ **FLOATING
C2480 a_11765_17973# vssd1 0.888f $ **FLOATING
C2481 _0490_ vssd1 6.03f $ **FLOATING
C2482 _0516_ vssd1 3.78f $ **FLOATING
C2483 cal_lut\[2\] vssd1 2.14f $ **FLOATING
C2484 a_8645_17999# vssd1 0.597f $ **FLOATING
C2485 a_7239_17999# vssd1 0.599f $ **FLOATING
C2486 a_7410_17973# vssd1 1.41f $ **FLOATING
C2487 a_6823_17999# vssd1 0.627f $ **FLOATING
C2488 a_6982_17973# vssd1 0.587f $ **FLOATING
C2489 a_6541_18005# vssd1 1.39f $ **FLOATING
C2490 _0195_ vssd1 1.09f $ **FLOATING
C2491 a_6375_18005# vssd1 1.77f $ **FLOATING
C2492 _0384_ vssd1 1.54f $ **FLOATING
C2493 net72 vssd1 4.29f $ **FLOATING
C2494 a_4995_17999# vssd1 0.698f $ **FLOATING
C2495 _0741_ vssd1 2.27f $ **FLOATING
C2496 a_3615_17999# vssd1 1.45f $ **FLOATING
C2497 a_2742_18082# vssd1 0.611f $ **FLOATING
C2498 net7 vssd1 4.44f $ **FLOATING
C2499 a_2288_17973# vssd1 0.648f $ **FLOATING
C2500 net5 vssd1 4.67f $ **FLOATING
C2501 a_1743_18259# vssd1 1.2f $ **FLOATING
C2502 a_26325_18543# vssd1 0.23f $ **FLOATING
C2503 a_26835_18909# vssd1 0.609f $ **FLOATING
C2504 a_27003_18811# vssd1 0.817f $ **FLOATING
C2505 a_26410_18909# vssd1 0.626f $ **FLOATING
C2506 a_26578_18655# vssd1 0.581f $ **FLOATING
C2507 a_26137_18543# vssd1 1.43f $ **FLOATING
C2508 a_25971_18543# vssd1 1.81f $ **FLOATING
C2509 cal_lut\[75\] vssd1 2.59f $ **FLOATING
C2510 _0246_ vssd1 15.3f $ **FLOATING
C2511 _0642_ vssd1 1.36f $ **FLOATING
C2512 _0648_ vssd1 7.81f $ **FLOATING
C2513 _0635_ vssd1 3.99f $ **FLOATING
C2514 _0643_ vssd1 0.843f $ **FLOATING
C2515 _0612_ vssd1 2.42f $ **FLOATING
C2516 _0605_ vssd1 3.37f $ **FLOATING
C2517 _0076_ vssd1 0.913f $ **FLOATING
C2518 _0492_ vssd1 10.2f $ **FLOATING
C2519 a_15959_18793# vssd1 0.388f $ **FLOATING
C2520 _0472_ vssd1 7.68f $ **FLOATING
C2521 a_14550_18793# vssd1 0.36f $ **FLOATING
C2522 a_14353_18793# vssd1 0.247f $ **FLOATING
C2523 a_14103_18793# vssd1 0.393f $ **FLOATING
C2524 a_8979_18543# vssd1 0.554f $ **FLOATING
C2525 a_12455_18793# vssd1 0.436f $ **FLOATING
C2526 a_12075_18793# vssd1 0.253f $ **FLOATING
C2527 a_9423_18793# vssd1 0.381f $ **FLOATING
C2528 a_8975_18793# vssd1 0.381f $ **FLOATING
C2529 a_7465_18543# vssd1 0.216f $ **FLOATING
C2530 a_25552_18793# vssd1 0.502f $ **FLOATING
C2531 a_23903_18695# vssd1 0.619f $ **FLOATING
C2532 a_23483_18909# vssd1 0.508f $ **FLOATING
C2533 cal_lut\[26\] vssd1 1.98f $ **FLOATING
C2534 a_23303_18909# vssd1 0.604f $ **FLOATING
C2535 a_22383_18793# vssd1 0.702f $ **FLOATING
C2536 a_21721_18909# vssd1 0.85f $ **FLOATING
C2537 a_21555_18909# vssd1 0.604f $ **FLOATING
C2538 a_20543_18543# vssd1 0.905f $ **FLOATING
C2539 a_20690_18517# vssd1 1.31f $ **FLOATING
C2540 a_20039_18695# vssd1 0.619f $ **FLOATING
C2541 a_19667_18517# vssd1 0.641f $ **FLOATING
C2542 a_19303_18695# vssd1 0.673f $ **FLOATING
C2543 a_18475_18695# vssd1 0.619f $ **FLOATING
C2544 a_17187_18708# vssd1 0.524f $ **FLOATING
C2545 _0491_ vssd1 4.84f $ **FLOATING
C2546 a_15207_18543# vssd1 0.887f $ **FLOATING
C2547 a_14770_18517# vssd1 0.649f $ **FLOATING
C2548 a_13291_18909# vssd1 0.795f $ **FLOATING
C2549 a_13508_18517# vssd1 0.788f $ **FLOATING
C2550 a_13091_18543# vssd1 0.696f $ **FLOATING
C2551 net15 vssd1 2.69f $ **FLOATING
C2552 net16 vssd1 2.01f $ **FLOATING
C2553 a_11857_18517# vssd1 0.55f $ **FLOATING
C2554 _0517_ vssd1 1.78f $ **FLOATING
C2555 _0520_ vssd1 1.58f $ **FLOATING
C2556 a_7975_18909# vssd1 0.599f $ **FLOATING
C2557 a_8146_18796# vssd1 1.41f $ **FLOATING
C2558 a_7559_18909# vssd1 0.627f $ **FLOATING
C2559 a_7718_18679# vssd1 0.587f $ **FLOATING
C2560 a_7277_18543# vssd1 1.39f $ **FLOATING
C2561 a_7111_18543# vssd1 1.77f $ **FLOATING
C2562 clknet_1_0__leaf_io_in[0] vssd1 15.5f $ **FLOATING
C2563 _0194_ vssd1 1.03f $ **FLOATING
C2564 a_6651_18793# vssd1 0.388f $ **FLOATING
C2565 a_4443_18793# vssd1 0.388f $ **FLOATING
C2566 a_2371_18523# vssd1 0.429f $ **FLOATING
C2567 _0426_ vssd1 1.83f $ **FLOATING
C2568 a_3995_18793# vssd1 0.642f $ **FLOATING
C2569 a_2747_18517# vssd1 0.698f $ **FLOATING
C2570 a_2099_18695# vssd1 0.67f $ **FLOATING
C2571 _0743_ vssd1 0.697f $ **FLOATING
C2572 a_1736_18517# vssd1 0.648f $ **FLOATING
C2573 _0075_ vssd1 0.975f $ **FLOATING
C2574 a_23565_19087# vssd1 0.23f $ **FLOATING
C2575 a_26063_19087# vssd1 0.524f $ **FLOATING
C2576 _0252_ vssd1 0.986f $ **FLOATING
C2577 a_25235_19087# vssd1 0.524f $ **FLOATING
C2578 _0870_ vssd1 0.675f $ **FLOATING
C2579 a_24863_19087# vssd1 0.508f $ **FLOATING
C2580 cal_lut\[27\] vssd1 1.67f $ **FLOATING
C2581 a_24683_19087# vssd1 0.604f $ **FLOATING
C2582 a_24075_19087# vssd1 0.609f $ **FLOATING
C2583 a_24243_19061# vssd1 0.817f $ **FLOATING
C2584 a_23650_19087# vssd1 0.626f $ **FLOATING
C2585 a_23818_19061# vssd1 0.581f $ **FLOATING
C2586 a_23377_19093# vssd1 1.43f $ **FLOATING
C2587 a_23211_19093# vssd1 1.81f $ **FLOATING
C2588 net42 vssd1 11.2f $ **FLOATING
C2589 a_19915_19087# vssd1 0.795f $ **FLOATING
C2590 a_20132_19394# vssd1 0.788f $ **FLOATING
C2591 a_19715_19087# vssd1 0.696f $ **FLOATING
C2592 a_19167_19061# vssd1 0.74f $ **FLOATING
C2593 a_19057_19319# vssd1 0.768f $ **FLOATING
C2594 _0253_ vssd1 0.883f $ **FLOATING
C2595 a_9503_19087# vssd1 0.238f $ **FLOATING
C2596 a_12437_19407# vssd1 0.18f $ **FLOATING
C2597 _0556_ vssd1 1.5f $ **FLOATING
C2598 a_11067_19407# vssd1 0.18f $ **FLOATING
C2599 a_18698_19319# vssd1 0.711f $ **FLOATING
C2600 a_18243_19200# vssd1 0.619f $ **FLOATING
C2601 _0507_ vssd1 2.02f $ **FLOATING
C2602 cal_lut\[70\] vssd1 5.25f $ **FLOATING
C2603 _0474_ vssd1 15.1f $ **FLOATING
C2604 a_17555_19319# vssd1 0.619f $ **FLOATING
C2605 a_17135_19087# vssd1 0.508f $ **FLOATING
C2606 cal_lut\[76\] vssd1 5.63f $ **FLOATING
C2607 a_16955_19087# vssd1 0.604f $ **FLOATING
C2608 a_15370_19407# vssd1 1.24f $ **FLOATING
C2609 a_15494_19319# vssd1 0.897f $ **FLOATING
C2610 a_15115_19087# vssd1 0.619f $ **FLOATING
C2611 a_13714_19407# vssd1 1.24f $ **FLOATING
C2612 a_13838_19319# vssd1 0.897f $ **FLOATING
C2613 a_13459_19087# vssd1 0.619f $ **FLOATING
C2614 cal_lut\[6\] vssd1 1.84f $ **FLOATING
C2615 _0519_ vssd1 7.15f $ **FLOATING
C2616 net4 vssd1 10.9f $ **FLOATING
C2617 a_10562_19319# vssd1 0.702f $ **FLOATING
C2618 _0590_ vssd1 2.61f $ **FLOATING
C2619 _0589_ vssd1 3.07f $ **FLOATING
C2620 a_5007_19087# vssd1 0.167f $ **FLOATING
C2621 a_4805_19087# vssd1 0.214f $ **FLOATING
C2622 a_4253_19087# vssd1 0.238f $ **FLOATING
C2623 a_2447_19087# vssd1 0.557f $ **FLOATING
C2624 _0383_ vssd1 1.03f $ **FLOATING
C2625 a_3435_19407# vssd1 0.211f $ **FLOATING
C2626 a_9933_19061# vssd1 0.858f $ **FLOATING
C2627 _0628_ vssd1 2.53f $ **FLOATING
C2628 _0439_ vssd1 3.12f $ **FLOATING
C2629 a_7157_19319# vssd1 0.767f $ **FLOATING
C2630 a_6979_19061# vssd1 0.83f $ **FLOATING
C2631 a_6375_19095# vssd1 0.648f $ **FLOATING
C2632 _0430_ vssd1 0.997f $ **FLOATING
C2633 a_4679_19319# vssd1 0.972f $ **FLOATING
C2634 _0742_ vssd1 0.954f $ **FLOATING
C2635 a_3299_19061# vssd1 0.791f $ **FLOATING
C2636 _0423_ vssd1 2.45f $ **FLOATING
C2637 _0745_ vssd1 1.1f $ **FLOATING
C2638 a_2023_19319# vssd1 1.33f $ **FLOATING
C2639 a_1471_19319# vssd1 0.611f $ **FLOATING
C2640 a_25389_19631# vssd1 0.23f $ **FLOATING
C2641 _0026_ vssd1 0.96f $ **FLOATING
C2642 _0027_ vssd1 0.955f $ **FLOATING
C2643 a_24971_19631# vssd1 0.581f $ **FLOATING
C2644 a_25042_19605# vssd1 0.626f $ **FLOATING
C2645 a_24835_19605# vssd1 1.81f $ **FLOATING
C2646 a_24842_19905# vssd1 1.43f $ **FLOATING
C2647 a_24551_19605# vssd1 0.609f $ **FLOATING
C2648 a_24455_19783# vssd1 0.817f $ **FLOATING
C2649 _0869_ vssd1 1.02f $ **FLOATING
C2650 a_23627_19796# vssd1 0.524f $ **FLOATING
C2651 a_22813_19631# vssd1 0.23f $ **FLOATING
C2652 a_20713_19631# vssd1 0.23f $ **FLOATING
C2653 a_22395_19631# vssd1 0.581f $ **FLOATING
C2654 a_22466_19605# vssd1 0.626f $ **FLOATING
C2655 a_22259_19605# vssd1 1.81f $ **FLOATING
C2656 a_22266_19905# vssd1 1.43f $ **FLOATING
C2657 a_21975_19605# vssd1 0.609f $ **FLOATING
C2658 a_21879_19783# vssd1 0.817f $ **FLOATING
C2659 a_21223_19997# vssd1 0.609f $ **FLOATING
C2660 a_21391_19899# vssd1 0.817f $ **FLOATING
C2661 a_20798_19997# vssd1 0.626f $ **FLOATING
C2662 a_20966_19743# vssd1 0.581f $ **FLOATING
C2663 a_20525_19631# vssd1 1.43f $ **FLOATING
C2664 a_20359_19631# vssd1 1.81f $ **FLOATING
C2665 cal_lut\[59\] vssd1 2.8f $ **FLOATING
C2666 a_19940_19881# vssd1 0.502f $ **FLOATING
C2667 a_19255_19631# vssd1 0.648f $ **FLOATING
C2668 net18 vssd1 9.68f $ **FLOATING
C2669 cal_lut\[28\] vssd1 5.19f $ **FLOATING
C2670 _0467_ vssd1 16.4f $ **FLOATING
C2671 a_17628_19881# vssd1 0.259f $ **FLOATING
C2672 cal_lut\[35\] vssd1 3.76f $ **FLOATING
C2673 a_15377_19631# vssd1 0.23f $ **FLOATING
C2674 a_18475_19783# vssd1 0.619f $ **FLOATING
C2675 a_18027_19783# vssd1 0.56f $ **FLOATING
C2676 _0579_ vssd1 0.974f $ **FLOATING
C2677 _0580_ vssd1 0.854f $ **FLOATING
C2678 a_17197_19777# vssd1 0.672f $ **FLOATING
C2679 a_15887_19997# vssd1 0.609f $ **FLOATING
C2680 a_16055_19899# vssd1 0.817f $ **FLOATING
C2681 a_15462_19997# vssd1 0.626f $ **FLOATING
C2682 a_15630_19743# vssd1 0.581f $ **FLOATING
C2683 a_15189_19631# vssd1 1.43f $ **FLOATING
C2684 a_15023_19631# vssd1 1.81f $ **FLOATING
C2685 _0034_ vssd1 0.872f $ **FLOATING
C2686 _0442_ vssd1 9.74f $ **FLOATING
C2687 a_10809_19605# vssd1 0.607f $ **FLOATING
C2688 _0629_ vssd1 3.41f $ **FLOATING
C2689 a_9429_19605# vssd1 0.607f $ **FLOATING
C2690 _0703_ vssd1 2.41f $ **FLOATING
C2691 a_8309_19881# vssd1 0.253f $ **FLOATING
C2692 clknet_1_0__leaf__0380_ vssd1 8.95f $ **FLOATING
C2693 a_4627_19631# vssd1 0.18f $ **FLOATING
C2694 a_4180_19631# vssd1 0.238f $ **FLOATING
C2695 a_3990_19631# vssd1 0.217f $ **FLOATING
C2696 a_5841_19605# vssd1 0.607f $ **FLOATING
C2697 a_5081_19881# vssd1 0.238f $ **FLOATING
C2698 _0740_ vssd1 0.856f $ **FLOATING
C2699 a_2614_19631# vssd1 0.255f $ **FLOATING
C2700 a_2107_19631# vssd1 0.19f $ **FLOATING
C2701 a_1917_19631# vssd1 0.19f $ **FLOATING
C2702 a_3112_19783# vssd1 0.732f $ **FLOATING
C2703 a_1917_19881# vssd1 0.667f $ **FLOATING
C2704 a_14747_19631# vssd1 0.524f $ **FLOATING
C2705 a_14167_19783# vssd1 0.658f $ **FLOATING
C2706 a_11191_19659# vssd1 0.56f $ **FLOATING
C2707 a_10380_19783# vssd1 0.59f $ **FLOATING
C2708 _0668_ vssd1 1.78f $ **FLOATING
C2709 a_9000_19783# vssd1 0.59f $ **FLOATING
C2710 a_8478_19631# vssd1 0.55f $ **FLOATING
C2711 _0764_ vssd1 0.907f $ **FLOATING
C2712 a_6537_19605# vssd1 4.03f $ **FLOATING
C2713 a_5412_19783# vssd1 0.59f $ **FLOATING
C2714 _0739_ vssd1 0.674f $ **FLOATING
C2715 _0738_ vssd1 0.894f $ **FLOATING
C2716 a_3799_19631# vssd1 0.893f $ **FLOATING
C2717 a_3072_19637# vssd1 0.719f $ **FLOATING
C2718 _0428_ vssd1 5.1f $ **FLOATING
C2719 a_1551_19605# vssd1 1.57f $ **FLOATING
C2720 a_26309_20553# vssd1 0.23f $ **FLOATING
C2721 a_24377_20553# vssd1 0.23f $ **FLOATING
C2722 _0058_ vssd1 1.02f $ **FLOATING
C2723 _0059_ vssd1 1.05f $ **FLOATING
C2724 a_25891_20553# vssd1 0.581f $ **FLOATING
C2725 a_25962_20452# vssd1 0.626f $ **FLOATING
C2726 a_25762_20297# vssd1 1.43f $ **FLOATING
C2727 a_25755_20393# vssd1 1.81f $ **FLOATING
C2728 a_25471_20407# vssd1 0.609f $ **FLOATING
C2729 a_25375_20407# vssd1 0.817f $ **FLOATING
C2730 a_23959_20553# vssd1 0.581f $ **FLOATING
C2731 a_24030_20452# vssd1 0.626f $ **FLOATING
C2732 a_23830_20297# vssd1 1.43f $ **FLOATING
C2733 a_23823_20393# vssd1 1.81f $ **FLOATING
C2734 a_23539_20407# vssd1 0.609f $ **FLOATING
C2735 a_23443_20407# vssd1 0.817f $ **FLOATING
C2736 a_22659_20175# vssd1 0.524f $ **FLOATING
C2737 _0233_ vssd1 0.867f $ **FLOATING
C2738 a_22291_20175# vssd1 0.698f $ **FLOATING
C2739 a_21872_20291# vssd1 0.502f $ **FLOATING
C2740 a_20359_20175# vssd1 0.524f $ **FLOATING
C2741 _0234_ vssd1 1.19f $ **FLOATING
C2742 a_18611_20288# vssd1 0.619f $ **FLOATING
C2743 _0461_ vssd1 2.17f $ **FLOATING
C2744 cal_lut\[58\] vssd1 3.02f $ **FLOATING
C2745 _0586_ vssd1 7.53f $ **FLOATING
C2746 _0582_ vssd1 0.927f $ **FLOATING
C2747 _0587_ vssd1 3.71f $ **FLOATING
C2748 _0602_ vssd1 3.85f $ **FLOATING
C2749 _0878_ vssd1 1.19f $ **FLOATING
C2750 a_13722_20175# vssd1 0.36f $ **FLOATING
C2751 a_13525_20175# vssd1 0.247f $ **FLOATING
C2752 a_13275_20175# vssd1 0.393f $ **FLOATING
C2753 a_5915_20175# vssd1 0.238f $ **FLOATING
C2754 a_4265_20175# vssd1 0.191f $ **FLOATING
C2755 net20 vssd1 13.2f $ **FLOATING
C2756 a_4719_20495# vssd1 0.171f $ **FLOATING
C2757 _0761_ vssd1 1.61f $ **FLOATING
C2758 a_17094_20407# vssd1 0.702f $ **FLOATING
C2759 a_16127_20288# vssd1 0.619f $ **FLOATING
C2760 cal_lut\[34\] vssd1 5.79f $ **FLOATING
C2761 a_15469_20407# vssd1 0.502f $ **FLOATING
C2762 a_14747_20175# vssd1 0.698f $ **FLOATING
C2763 a_13942_20149# vssd1 0.649f $ **FLOATING
C2764 a_12263_20495# vssd1 1.31f $ **FLOATING
C2765 a_12258_20407# vssd1 0.905f $ **FLOATING
C2766 _0666_ vssd1 2.45f $ **FLOATING
C2767 _0667_ vssd1 1.71f $ **FLOATING
C2768 a_6458_20175# vssd1 4.03f $ **FLOATING
C2769 a_4892_20175# vssd1 0.546f $ **FLOATING
C2770 _0447_ vssd1 13.2f $ **FLOATING
C2771 a_4128_20149# vssd1 0.847f $ **FLOATING
C2772 a_3525_20291# vssd1 0.665f $ **FLOATING
C2773 _0421_ vssd1 9.34f $ **FLOATING
C2774 a_2722_20175# vssd1 1.17f $ **FLOATING
C2775 _0420_ vssd1 7.48f $ **FLOATING
C2776 _0422_ vssd1 8.42f $ **FLOATING
C2777 a_2750_20407# vssd1 0.786f $ **FLOATING
C2778 _0033_ vssd1 1.35f $ **FLOATING
C2779 _0057_ vssd1 1.23f $ **FLOATING
C2780 cal_lut\[30\] vssd1 3.07f $ **FLOATING
C2781 _0536_ vssd1 4.33f $ **FLOATING
C2782 _0561_ vssd1 8.33f $ **FLOATING
C2783 a_19256_20969# vssd1 0.259f $ **FLOATING
C2784 _0552_ vssd1 2.87f $ **FLOATING
C2785 _0581_ vssd1 1.65f $ **FLOATING
C2786 _0495_ vssd1 19.4f $ **FLOATING
C2787 a_11508_20719# vssd1 0.337f $ **FLOATING
C2788 a_10975_20719# vssd1 0.28f $ **FLOATING
C2789 net17 vssd1 8.32f $ **FLOATING
C2790 a_11422_20969# vssd1 0.324f $ **FLOATING
C2791 a_10413_20969# vssd1 0.206f $ **FLOATING
C2792 a_6929_20719# vssd1 0.186f $ **FLOATING
C2793 a_9613_20693# vssd1 0.607f $ **FLOATING
C2794 _0626_ vssd1 4.92f $ **FLOATING
C2795 a_25235_20719# vssd1 0.524f $ **FLOATING
C2796 _0877_ vssd1 0.686f $ **FLOATING
C2797 a_24771_21085# vssd1 0.508f $ **FLOATING
C2798 a_24591_21085# vssd1 0.604f $ **FLOATING
C2799 a_23579_20719# vssd1 0.524f $ **FLOATING
C2800 a_22891_20871# vssd1 0.619f $ **FLOATING
C2801 a_21279_20719# vssd1 0.524f $ **FLOATING
C2802 _0874_ vssd1 0.68f $ **FLOATING
C2803 a_20860_20969# vssd1 0.502f $ **FLOATING
C2804 a_20359_20719# vssd1 0.619f $ **FLOATING
C2805 a_19426_20719# vssd1 0.672f $ **FLOATING
C2806 _0560_ vssd1 1.19f $ **FLOATING
C2807 _0559_ vssd1 1.88f $ **FLOATING
C2808 a_18763_20871# vssd1 0.56f $ **FLOATING
C2809 a_16955_20719# vssd1 0.619f $ **FLOATING
C2810 a_15667_20719# vssd1 0.619f $ **FLOATING
C2811 a_15023_20719# vssd1 0.524f $ **FLOATING
C2812 _0448_ vssd1 2.05f $ **FLOATING
C2813 a_14604_20969# vssd1 0.502f $ **FLOATING
C2814 _0485_ vssd1 6.49f $ **FLOATING
C2815 a_14153_20884# vssd1 0.524f $ **FLOATING
C2816 _0883_ vssd1 5.06f $ **FLOATING
C2817 a_13415_20884# vssd1 0.524f $ **FLOATING
C2818 a_12815_20719# vssd1 1.2f $ **FLOATING
C2819 a_10975_20969# vssd1 1.14f $ **FLOATING
C2820 _0676_ vssd1 1.56f $ **FLOATING
C2821 _0678_ vssd1 1.46f $ **FLOATING
C2822 a_10331_20969# vssd1 0.804f $ **FLOATING
C2823 a_9184_20871# vssd1 0.59f $ **FLOATING
C2824 a_8397_20983# vssd1 0.601f $ **FLOATING
C2825 a_8297_20765# vssd1 0.488f $ **FLOATING
C2826 a_7583_20969# vssd1 0.167f $ **FLOATING
C2827 a_7381_20969# vssd1 0.214f $ **FLOATING
C2828 a_6646_21041# vssd1 0.538f $ **FLOATING
C2829 _0425_ vssd1 14.2f $ **FLOATING
C2830 a_2137_20719# vssd1 0.171f $ **FLOATING
C2831 _0736_ vssd1 1.58f $ **FLOATING
C2832 a_5099_20969# vssd1 0.167f $ **FLOATING
C2833 a_4897_20969# vssd1 0.214f $ **FLOATING
C2834 a_2695_20969# vssd1 0.436f $ **FLOATING
C2835 _0762_ vssd1 1.64f $ **FLOATING
C2836 _0433_ vssd1 11f $ **FLOATING
C2837 _0767_ vssd1 1.56f $ **FLOATING
C2838 _0766_ vssd1 1.48f $ **FLOATING
C2839 a_7255_20871# vssd1 0.972f $ **FLOATING
C2840 a_6516_20871# vssd1 0.645f $ **FLOATING
C2841 _0769_ vssd1 0.769f $ **FLOATING
C2842 _0768_ vssd1 1.54f $ **FLOATING
C2843 _0438_ vssd1 12.9f $ **FLOATING
C2844 a_4771_20871# vssd1 0.972f $ **FLOATING
C2845 ctr\[2\] vssd1 10.6f $ **FLOATING
C2846 a_1919_20693# vssd1 0.546f $ **FLOATING
C2847 _0232_ vssd1 0.892f $ **FLOATING
C2848 a_22872_21263# vssd1 0.259f $ **FLOATING
C2849 _0639_ vssd1 1.75f $ **FLOATING
C2850 cal_lut\[66\] vssd1 3.91f $ **FLOATING
C2851 a_20437_21263# vssd1 0.23f $ **FLOATING
C2852 _0558_ vssd1 0.889f $ **FLOATING
C2853 a_14917_21263# vssd1 0.23f $ **FLOATING
C2854 cal_lut\[40\] vssd1 1.98f $ **FLOATING
C2855 a_13261_21263# vssd1 0.23f $ **FLOATING
C2856 a_10715_21263# vssd1 0.386f $ **FLOATING
C2857 a_10521_21263# vssd1 0.23f $ **FLOATING
C2858 a_25787_21263# vssd1 0.524f $ **FLOATING
C2859 a_23391_21263# vssd1 0.508f $ **FLOATING
C2860 a_23211_21263# vssd1 0.604f $ **FLOATING
C2861 _0636_ vssd1 0.804f $ **FLOATING
C2862 _0637_ vssd1 0.815f $ **FLOATING
C2863 a_22441_21237# vssd1 0.672f $ **FLOATING
C2864 a_21923_21376# vssd1 0.619f $ **FLOATING
C2865 a_20947_21263# vssd1 0.609f $ **FLOATING
C2866 a_21115_21237# vssd1 0.817f $ **FLOATING
C2867 a_20522_21263# vssd1 0.626f $ **FLOATING
C2868 a_20690_21237# vssd1 0.581f $ **FLOATING
C2869 a_20249_21269# vssd1 1.43f $ **FLOATING
C2870 a_20083_21269# vssd1 1.81f $ **FLOATING
C2871 a_19439_21263# vssd1 0.698f $ **FLOATING
C2872 a_18979_21376# vssd1 0.619f $ **FLOATING
C2873 a_18519_21263# vssd1 0.698f $ **FLOATING
C2874 a_18151_21271# vssd1 0.648f $ **FLOATING
C2875 a_17783_21271# vssd1 0.648f $ **FLOATING
C2876 _0453_ vssd1 5.95f $ **FLOATING
C2877 _0214_ vssd1 0.836f $ **FLOATING
C2878 a_16727_21482# vssd1 0.524f $ **FLOATING
C2879 a_16076_21379# vssd1 0.502f $ **FLOATING
C2880 cal_lut\[41\] vssd1 1.75f $ **FLOATING
C2881 a_15427_21263# vssd1 0.609f $ **FLOATING
C2882 a_15595_21237# vssd1 0.817f $ **FLOATING
C2883 a_15002_21263# vssd1 0.626f $ **FLOATING
C2884 a_15170_21237# vssd1 0.581f $ **FLOATING
C2885 a_14729_21269# vssd1 1.43f $ **FLOATING
C2886 a_14563_21269# vssd1 1.81f $ **FLOATING
C2887 a_13771_21263# vssd1 0.609f $ **FLOATING
C2888 a_13939_21237# vssd1 0.817f $ **FLOATING
C2889 a_13346_21263# vssd1 0.626f $ **FLOATING
C2890 a_13514_21237# vssd1 0.581f $ **FLOATING
C2891 a_13073_21269# vssd1 1.43f $ **FLOATING
C2892 _0039_ vssd1 1.05f $ **FLOATING
C2893 a_12907_21269# vssd1 1.81f $ **FLOATING
C2894 a_12355_21271# vssd1 0.648f $ **FLOATING
C2895 a_11715_21379# vssd1 0.67f $ **FLOATING
C2896 a_11609_21379# vssd1 0.429f $ **FLOATING
C2897 a_10247_21583# vssd1 0.59f $ **FLOATING
C2898 a_9821_21583# vssd1 0.187f $ **FLOATING
C2899 a_8025_21263# vssd1 0.238f $ **FLOATING
C2900 a_7393_21263# vssd1 0.191f $ **FLOATING
C2901 a_6847_21263# vssd1 0.167f $ **FLOATING
C2902 a_6645_21263# vssd1 0.214f $ **FLOATING
C2903 a_5915_21263# vssd1 0.238f $ **FLOATING
C2904 a_5547_21263# vssd1 0.238f $ **FLOATING
C2905 a_4087_21263# vssd1 0.167f $ **FLOATING
C2906 a_3885_21263# vssd1 0.214f $ **FLOATING
C2907 a_2605_21263# vssd1 0.203f $ **FLOATING
C2908 _0670_ vssd1 3.54f $ **FLOATING
C2909 _0677_ vssd1 1.75f $ **FLOATING
C2910 a_4713_21583# vssd1 0.171f $ **FLOATING
C2911 a_9671_21495# vssd1 0.743f $ **FLOATING
C2912 a_9167_21601# vssd1 0.56f $ **FLOATING
C2913 _0557_ vssd1 4.34f $ **FLOATING
C2914 _0591_ vssd1 4.83f $ **FLOATING
C2915 _0627_ vssd1 2.72f $ **FLOATING
C2916 a_7256_21237# vssd1 0.847f $ **FLOATING
C2917 _0779_ vssd1 0.933f $ **FLOATING
C2918 _0778_ vssd1 0.713f $ **FLOATING
C2919 a_6519_21495# vssd1 0.972f $ **FLOATING
C2920 a_4495_21495# vssd1 0.546f $ **FLOATING
C2921 _0781_ vssd1 0.625f $ **FLOATING
C2922 _0780_ vssd1 1.96f $ **FLOATING
C2923 _0446_ vssd1 16.1f $ **FLOATING
C2924 _0427_ vssd1 5.1f $ **FLOATING
C2925 a_3759_21495# vssd1 0.972f $ **FLOATING
C2926 a_2511_21263# vssd1 0.796f $ **FLOATING
C2927 _0771_ vssd1 0.744f $ **FLOATING
C2928 _0770_ vssd1 1.68f $ **FLOATING
C2929 _0772_ vssd1 0.638f $ **FLOATING
C2930 a_1963_21365# vssd1 0.753f $ **FLOATING
C2931 a_1857_21365# vssd1 0.454f $ **FLOATING
C2932 a_26693_21807# vssd1 0.23f $ **FLOATING
C2933 a_27203_22173# vssd1 0.609f $ **FLOATING
C2934 a_27371_22075# vssd1 0.817f $ **FLOATING
C2935 a_26778_22173# vssd1 0.626f $ **FLOATING
C2936 a_26946_21919# vssd1 0.581f $ **FLOATING
C2937 a_26505_21807# vssd1 1.43f $ **FLOATING
C2938 _0063_ vssd1 1.18f $ **FLOATING
C2939 a_26339_21807# vssd1 1.81f $ **FLOATING
C2940 a_25849_21807# vssd1 0.23f $ **FLOATING
C2941 cal_lut\[33\] vssd1 2.44f $ **FLOATING
C2942 _0638_ vssd1 1.22f $ **FLOATING
C2943 _0462_ vssd1 17.1f $ **FLOATING
C2944 a_21725_21807# vssd1 0.23f $ **FLOATING
C2945 _0032_ vssd1 1.24f $ **FLOATING
C2946 a_25431_21807# vssd1 0.581f $ **FLOATING
C2947 a_25502_21781# vssd1 0.626f $ **FLOATING
C2948 a_25295_21781# vssd1 1.81f $ **FLOATING
C2949 a_25302_22081# vssd1 1.43f $ **FLOATING
C2950 a_25011_21781# vssd1 0.609f $ **FLOATING
C2951 a_24915_21959# vssd1 0.817f $ **FLOATING
C2952 a_24591_21807# vssd1 0.524f $ **FLOATING
C2953 a_23351_21959# vssd1 0.619f $ **FLOATING
C2954 a_22903_21959# vssd1 0.56f $ **FLOATING
C2955 a_22235_22173# vssd1 0.609f $ **FLOATING
C2956 a_22403_22075# vssd1 0.817f $ **FLOATING
C2957 a_21810_22173# vssd1 0.626f $ **FLOATING
C2958 a_21978_21919# vssd1 0.581f $ **FLOATING
C2959 a_21537_21807# vssd1 1.43f $ **FLOATING
C2960 _0030_ vssd1 1.19f $ **FLOATING
C2961 a_21371_21807# vssd1 1.81f $ **FLOATING
C2962 net43 vssd1 9.43f $ **FLOATING
C2963 _0065_ vssd1 1.03f $ **FLOATING
C2964 cal_lut\[64\] vssd1 5.22f $ **FLOATING
C2965 _0443_ vssd1 15.2f $ **FLOATING
C2966 _0553_ vssd1 3.19f $ **FLOATING
C2967 a_16481_21807# vssd1 0.23f $ **FLOATING
C2968 _0241_ vssd1 0.758f $ **FLOATING
C2969 a_20683_21972# vssd1 0.524f $ **FLOATING
C2970 a_20216_22057# vssd1 0.502f $ **FLOATING
C2971 a_19793_21959# vssd1 0.502f $ **FLOATING
C2972 a_19287_21835# vssd1 0.56f $ **FLOATING
C2973 a_17739_21959# vssd1 0.619f $ **FLOATING
C2974 a_16991_22173# vssd1 0.609f $ **FLOATING
C2975 a_17159_22075# vssd1 0.817f $ **FLOATING
C2976 a_16566_22173# vssd1 0.626f $ **FLOATING
C2977 a_16734_21919# vssd1 0.581f $ **FLOATING
C2978 a_16293_21807# vssd1 1.43f $ **FLOATING
C2979 _0041_ vssd1 1.03f $ **FLOATING
C2980 a_16127_21807# vssd1 1.81f $ **FLOATING
C2981 _0040_ vssd1 0.977f $ **FLOATING
C2982 a_15727_21959# vssd1 0.56f $ **FLOATING
C2983 _0213_ vssd1 1.22f $ **FLOATING
C2984 a_14703_21972# vssd1 0.524f $ **FLOATING
C2985 a_13459_21807# vssd1 0.648f $ **FLOATING
C2986 a_11799_22057# vssd1 0.253f $ **FLOATING
C2987 a_11014_22057# vssd1 0.333f $ **FLOATING
C2988 a_4472_21807# vssd1 0.215f $ **FLOATING
C2989 a_4381_21807# vssd1 0.118f $ **FLOATING
C2990 _0630_ vssd1 2.78f $ **FLOATING
C2991 _0669_ vssd1 4.89f $ **FLOATING
C2992 a_6463_22057# vssd1 0.253f $ **FLOATING
C2993 a_5911_22057# vssd1 0.253f $ **FLOATING
C2994 a_5359_22057# vssd1 0.253f $ **FLOATING
C2995 _0760_ vssd1 1.47f $ **FLOATING
C2996 a_3891_22057# vssd1 0.238f $ **FLOATING
C2997 a_1679_22057# vssd1 0.253f $ **FLOATING
C2998 a_12723_21807# vssd1 1.2f $ **FLOATING
C2999 a_12127_21959# vssd1 0.619f $ **FLOATING
C3000 _0673_ vssd1 2.36f $ **FLOATING
C3001 a_11581_21781# vssd1 0.55f $ **FLOATING
C3002 _0521_ vssd1 4.82f $ **FLOATING
C3003 a_10857_21781# vssd1 0.723f $ **FLOATING
C3004 a_10372_22057# vssd1 0.502f $ **FLOATING
C3005 a_7102_21807# vssd1 4.03f $ **FLOATING
C3006 _0380_ vssd1 4.92f $ **FLOATING
C3007 a_6245_21781# vssd1 0.55f $ **FLOATING
C3008 a_5693_21781# vssd1 0.55f $ **FLOATING
C3009 a_5141_21781# vssd1 0.55f $ **FLOATING
C3010 a_4283_22057# vssd1 0.869f $ **FLOATING
C3011 _0758_ vssd1 1.02f $ **FLOATING
C3012 _0757_ vssd1 0.714f $ **FLOATING
C3013 _0756_ vssd1 0.944f $ **FLOATING
C3014 a_2419_21807# vssd1 1.2f $ **FLOATING
C3015 a_1959_21807# vssd1 0.698f $ **FLOATING
C3016 _0763_ vssd1 0.844f $ **FLOATING
C3017 a_1461_21781# vssd1 0.55f $ **FLOATING
C3018 _0239_ vssd1 1.06f $ **FLOATING
C3019 _0876_ vssd1 1f $ **FLOATING
C3020 a_19100_22351# vssd1 0.259f $ **FLOATING
C3021 a_20161_22351# vssd1 0.23f $ **FLOATING
C3022 _0621_ vssd1 3.77f $ **FLOATING
C3023 a_7853_22351# vssd1 0.191f $ **FLOATING
C3024 a_6939_22351# vssd1 0.167f $ **FLOATING
C3025 a_6737_22351# vssd1 0.214f $ **FLOATING
C3026 a_2485_22351# vssd1 0.203f $ **FLOATING
C3027 a_11756_22671# vssd1 0.206f $ **FLOATING
C3028 a_8533_22671# vssd1 0.187f $ **FLOATING
C3029 _0777_ vssd1 1.44f $ **FLOATING
C3030 a_5643_22671# vssd1 0.211f $ **FLOATING
C3031 a_3067_22671# vssd1 0.211f $ **FLOATING
C3032 _0413_ vssd1 0.995f $ **FLOATING
C3033 a_25415_22351# vssd1 0.508f $ **FLOATING
C3034 a_25235_22351# vssd1 0.604f $ **FLOATING
C3035 a_24679_22351# vssd1 0.508f $ **FLOATING
C3036 a_24499_22351# vssd1 0.604f $ **FLOATING
C3037 a_23763_22351# vssd1 0.524f $ **FLOATING
C3038 _0875_ vssd1 0.647f $ **FLOATING
C3039 a_23391_22351# vssd1 0.508f $ **FLOATING
C3040 a_23211_22351# vssd1 0.604f $ **FLOATING
C3041 _0863_ vssd1 19.4f $ **FLOATING
C3042 a_20671_22351# vssd1 0.609f $ **FLOATING
C3043 a_20839_22325# vssd1 0.817f $ **FLOATING
C3044 a_20246_22351# vssd1 0.626f $ **FLOATING
C3045 a_20414_22325# vssd1 0.581f $ **FLOATING
C3046 a_19973_22357# vssd1 1.43f $ **FLOATING
C3047 _0064_ vssd1 0.872f $ **FLOATING
C3048 a_19807_22357# vssd1 1.81f $ **FLOATING
C3049 net44 vssd1 14.6f $ **FLOATING
C3050 a_19531_22351# vssd1 0.524f $ **FLOATING
C3051 _0240_ vssd1 1.09f $ **FLOATING
C3052 cal_lut\[65\] vssd1 2.36f $ **FLOATING
C3053 a_18669_22325# vssd1 0.672f $ **FLOATING
C3054 a_16803_22689# vssd1 0.56f $ **FLOATING
C3055 a_15023_22464# vssd1 0.619f $ **FLOATING
C3056 _0483_ vssd1 13.5f $ **FLOATING
C3057 _0531_ vssd1 17.8f $ **FLOATING
C3058 a_13459_22359# vssd1 0.648f $ **FLOATING
C3059 _0838_ vssd1 16.4f $ **FLOATING
C3060 a_13144_22325# vssd1 0.648f $ **FLOATING
C3061 a_12723_22351# vssd1 0.524f $ **FLOATING
C3062 _0258_ vssd1 3.92f $ **FLOATING
C3063 _0671_ vssd1 2.69f $ **FLOATING
C3064 _0665_ vssd1 2.51f $ **FLOATING
C3065 _0631_ vssd1 2.84f $ **FLOATING
C3066 _0664_ vssd1 4.41f $ **FLOATING
C3067 _0709_ vssd1 0.833f $ **FLOATING
C3068 _0674_ vssd1 1.25f $ **FLOATING
C3069 _0672_ vssd1 2f $ **FLOATING
C3070 a_8383_22583# vssd1 0.743f $ **FLOATING
C3071 _0785_ vssd1 1.25f $ **FLOATING
C3072 a_7716_22325# vssd1 0.847f $ **FLOATING
C3073 _0787_ vssd1 1.71f $ **FLOATING
C3074 _0786_ vssd1 0.868f $ **FLOATING
C3075 _0432_ vssd1 7.55f $ **FLOATING
C3076 a_6611_22583# vssd1 0.972f $ **FLOATING
C3077 _0788_ vssd1 0.819f $ **FLOATING
C3078 ctr\[4\] vssd1 14.1f $ **FLOATING
C3079 a_5507_22325# vssd1 0.791f $ **FLOATING
C3080 clknet_0_net67 vssd1 8.39f $ **FLOATING
C3081 a_3685_22325# vssd1 4.03f $ **FLOATING
C3082 _0782_ vssd1 1.14f $ **FLOATING
C3083 a_2931_22325# vssd1 0.791f $ **FLOATING
C3084 _0783_ vssd1 0.643f $ **FLOATING
C3085 a_2287_22325# vssd1 0.796f $ **FLOATING
C3086 a_1773_22467# vssd1 0.601f $ **FLOATING
C3087 a_1673_22351# vssd1 0.488f $ **FLOATING
C3088 a_24761_22895# vssd1 0.23f $ **FLOATING
C3089 a_25271_23261# vssd1 0.609f $ **FLOATING
C3090 a_25439_23163# vssd1 0.817f $ **FLOATING
C3091 a_24846_23261# vssd1 0.626f $ **FLOATING
C3092 a_25014_23007# vssd1 0.581f $ **FLOATING
C3093 a_24573_22895# vssd1 1.43f $ **FLOATING
C3094 _0031_ vssd1 1.21f $ **FLOATING
C3095 a_24407_22895# vssd1 1.81f $ **FLOATING
C3096 a_23201_23145# vssd1 0.206f $ **FLOATING
C3097 _0686_ vssd1 3.47f $ **FLOATING
C3098 a_22457_23145# vssd1 0.214f $ **FLOATING
C3099 a_22373_23145# vssd1 0.167f $ **FLOATING
C3100 cal_lut\[60\] vssd1 3.41f $ **FLOATING
C3101 _0522_ vssd1 5.55f $ **FLOATING
C3102 _0619_ vssd1 1.19f $ **FLOATING
C3103 _0618_ vssd1 0.907f $ **FLOATING
C3104 _0452_ vssd1 17.1f $ **FLOATING
C3105 _0454_ vssd1 14.8f $ **FLOATING
C3106 _0465_ vssd1 11.5f $ **FLOATING
C3107 a_17129_23145# vssd1 0.206f $ **FLOATING
C3108 _0578_ vssd1 2.08f $ **FLOATING
C3109 _0647_ vssd1 5.64f $ **FLOATING
C3110 a_15208_23145# vssd1 0.259f $ **FLOATING
C3111 net81 vssd1 2.6f $ **FLOATING
C3112 a_12893_22895# vssd1 0.23f $ **FLOATING
C3113 cal_lut\[32\] vssd1 2.78f $ **FLOATING
C3114 a_23055_23047# vssd1 0.804f $ **FLOATING
C3115 a_22291_22895# vssd1 0.972f $ **FLOATING
C3116 a_21136_23145# vssd1 0.502f $ **FLOATING
C3117 a_19807_22895# vssd1 0.619f $ **FLOATING
C3118 a_19303_23047# vssd1 0.619f $ **FLOATING
C3119 a_18611_22895# vssd1 0.619f $ **FLOATING
C3120 a_17999_22923# vssd1 0.56f $ **FLOATING
C3121 _0500_ vssd1 9.7f $ **FLOATING
C3122 a_16983_23047# vssd1 0.804f $ **FLOATING
C3123 a_16069_22923# vssd1 0.713f $ **FLOATING
C3124 a_15378_22895# vssd1 0.672f $ **FLOATING
C3125 _0646_ vssd1 1.06f $ **FLOATING
C3126 _0644_ vssd1 0.903f $ **FLOATING
C3127 a_14287_22895# vssd1 0.619f $ **FLOATING
C3128 a_13403_23261# vssd1 0.609f $ **FLOATING
C3129 a_13571_23163# vssd1 0.817f $ **FLOATING
C3130 a_12978_23261# vssd1 0.626f $ **FLOATING
C3131 a_13146_23007# vssd1 0.581f $ **FLOATING
C3132 a_12705_22895# vssd1 1.43f $ **FLOATING
C3133 _0081_ vssd1 0.955f $ **FLOATING
C3134 a_12539_22895# vssd1 1.81f $ **FLOATING
C3135 a_9209_22895# vssd1 0.211f $ **FLOATING
C3136 _0710_ vssd1 1.26f $ **FLOATING
C3137 a_8485_23145# vssd1 0.238f $ **FLOATING
C3138 _0775_ vssd1 2.02f $ **FLOATING
C3139 _0774_ vssd1 0.966f $ **FLOATING
C3140 a_5813_22895# vssd1 0.18f $ **FLOATING
C3141 a_10915_22923# vssd1 0.56f $ **FLOATING
C3142 _0716_ vssd1 2.75f $ **FLOATING
C3143 a_9673_23047# vssd1 0.502f $ **FLOATING
C3144 a_8971_22895# vssd1 0.706f $ **FLOATING
C3145 _0704_ vssd1 2.7f $ **FLOATING
C3146 a_7939_22895# vssd1 0.619f $ **FLOATING
C3147 a_6182_22895# vssd1 4.03f $ **FLOATING
C3148 clknet_0_io_in[0] vssd1 6.84f $ **FLOATING
C3149 a_3882_22895# vssd1 4.03f $ **FLOATING
C3150 a_2939_23047# vssd1 0.56f $ **FLOATING
C3151 a_2327_22895# vssd1 0.988f $ **FLOATING
C3152 _0417_ vssd1 1.79f $ **FLOATING
C3153 cal_lut\[63\] vssd1 3.25f $ **FLOATING
C3154 a_23683_23439# vssd1 0.167f $ **FLOATING
C3155 a_23481_23439# vssd1 0.214f $ **FLOATING
C3156 a_25313_23439# vssd1 0.23f $ **FLOATING
C3157 _0471_ vssd1 3.34f $ **FLOATING
C3158 a_22185_23439# vssd1 0.23f $ **FLOATING
C3159 _0523_ vssd1 5.27f $ **FLOATING
C3160 _0620_ vssd1 1.16f $ **FLOATING
C3161 _0464_ vssd1 10.4f $ **FLOATING
C3162 cal_lut\[95\] vssd1 3.48f $ **FLOATING
C3163 a_15009_23439# vssd1 0.23f $ **FLOATING
C3164 cal_lut\[10\] vssd1 5.48f $ **FLOATING
C3165 a_13445_23439# vssd1 0.23f $ **FLOATING
C3166 a_10603_23439# vssd1 0.253f $ **FLOATING
C3167 a_7101_23439# vssd1 0.206f $ **FLOATING
C3168 a_6619_23439# vssd1 0.245f $ **FLOATING
C3169 _0717_ vssd1 1.61f $ **FLOATING
C3170 a_5545_23439# vssd1 0.203f $ **FLOATING
C3171 _0776_ vssd1 2.77f $ **FLOATING
C3172 _0753_ vssd1 2.56f $ **FLOATING
C3173 a_4997_23805# vssd1 0.186f $ **FLOATING
C3174 a_4040_23759# vssd1 0.118f $ **FLOATING
C3175 a_3850_23759# vssd1 0.215f $ **FLOATING
C3176 a_1867_23759# vssd1 0.279f $ **FLOATING
C3177 a_25823_23439# vssd1 0.609f $ **FLOATING
C3178 a_25991_23413# vssd1 0.817f $ **FLOATING
C3179 a_25398_23439# vssd1 0.626f $ **FLOATING
C3180 a_25566_23413# vssd1 0.581f $ **FLOATING
C3181 a_25125_23445# vssd1 1.43f $ **FLOATING
C3182 _0062_ vssd1 0.872f $ **FLOATING
C3183 a_24959_23445# vssd1 1.81f $ **FLOATING
C3184 a_24683_23439# vssd1 0.524f $ **FLOATING
C3185 _0470_ vssd1 1.18f $ **FLOATING
C3186 _0466_ vssd1 4.45f $ **FLOATING
C3187 _0463_ vssd1 1.95f $ **FLOATING
C3188 a_23355_23671# vssd1 0.972f $ **FLOATING
C3189 a_22695_23439# vssd1 0.609f $ **FLOATING
C3190 a_22863_23413# vssd1 0.817f $ **FLOATING
C3191 a_22270_23439# vssd1 0.626f $ **FLOATING
C3192 a_22438_23413# vssd1 0.581f $ **FLOATING
C3193 a_21997_23445# vssd1 1.43f $ **FLOATING
C3194 _0060_ vssd1 0.983f $ **FLOATING
C3195 a_21831_23445# vssd1 1.81f $ **FLOATING
C3196 a_21279_23439# vssd1 0.524f $ **FLOATING
C3197 _0235_ vssd1 0.986f $ **FLOATING
C3198 a_20451_23439# vssd1 1.2f $ **FLOATING
C3199 a_19623_23552# vssd1 0.619f $ **FLOATING
C3200 _0459_ vssd1 10f $ **FLOATING
C3201 a_18751_23671# vssd1 0.619f $ **FLOATING
C3202 a_17323_23439# vssd1 0.524f $ **FLOATING
C3203 _0259_ vssd1 0.647f $ **FLOATING
C3204 a_16951_23439# vssd1 0.508f $ **FLOATING
C3205 cal_lut\[82\] vssd1 2.9f $ **FLOATING
C3206 a_16771_23439# vssd1 0.604f $ **FLOATING
C3207 a_16187_23671# vssd1 0.56f $ **FLOATING
C3208 a_15519_23439# vssd1 0.609f $ **FLOATING
C3209 a_15687_23413# vssd1 0.817f $ **FLOATING
C3210 a_15094_23439# vssd1 0.626f $ **FLOATING
C3211 a_15262_23413# vssd1 0.581f $ **FLOATING
C3212 a_14821_23445# vssd1 1.43f $ **FLOATING
C3213 a_14655_23445# vssd1 1.81f $ **FLOATING
C3214 a_13955_23439# vssd1 0.609f $ **FLOATING
C3215 a_14123_23413# vssd1 0.817f $ **FLOATING
C3216 a_13530_23439# vssd1 0.626f $ **FLOATING
C3217 a_13698_23413# vssd1 0.581f $ **FLOATING
C3218 a_13257_23445# vssd1 1.43f $ **FLOATING
C3219 a_13091_23445# vssd1 1.81f $ **FLOATING
C3220 a_12723_23439# vssd1 0.698f $ **FLOATING
C3221 a_10943_23671# vssd1 0.56f $ **FLOATING
C3222 _0679_ vssd1 4.09f $ **FLOATING
C3223 _0675_ vssd1 3.38f $ **FLOATING
C3224 _0680_ vssd1 3.59f $ **FLOATING
C3225 a_10385_23413# vssd1 0.55f $ **FLOATING
C3226 a_8390_23439# vssd1 4.03f $ **FLOATING
C3227 clknet_0__0380_ vssd1 6.06f $ **FLOATING
C3228 a_6955_23671# vssd1 0.804f $ **FLOATING
C3229 _0434_ vssd1 10.2f $ **FLOATING
C3230 _0435_ vssd1 3.19f $ **FLOATING
C3231 _0755_ vssd1 10.8f $ **FLOATING
C3232 _0820_ vssd1 1.4f $ **FLOATING
C3233 _0818_ vssd1 0.877f $ **FLOATING
C3234 _0819_ vssd1 3.25f $ **FLOATING
C3235 a_5416_23413# vssd1 0.655f $ **FLOATING
C3236 a_4714_23483# vssd1 0.538f $ **FLOATING
C3237 _0821_ vssd1 0.918f $ **FLOATING
C3238 a_4584_23671# vssd1 0.645f $ **FLOATING
C3239 _0789_ vssd1 1.55f $ **FLOATING
C3240 _0790_ vssd1 3.21f $ **FLOATING
C3241 a_3695_23671# vssd1 0.869f $ **FLOATING
C3242 a_24761_23983# vssd1 0.23f $ **FLOATING
C3243 a_25271_24349# vssd1 0.609f $ **FLOATING
C3244 a_25439_24251# vssd1 0.817f $ **FLOATING
C3245 a_24846_24349# vssd1 0.626f $ **FLOATING
C3246 a_25014_24095# vssd1 0.581f $ **FLOATING
C3247 a_24573_23983# vssd1 1.43f $ **FLOATING
C3248 a_24407_23983# vssd1 1.81f $ **FLOATING
C3249 _0061_ vssd1 1.07f $ **FLOATING
C3250 a_22649_24233# vssd1 0.206f $ **FLOATING
C3251 _0685_ vssd1 1.08f $ **FLOATING
C3252 cal_lut\[83\] vssd1 1.69f $ **FLOATING
C3253 a_17677_23983# vssd1 0.23f $ **FLOATING
C3254 a_23671_23983# vssd1 0.524f $ **FLOATING
C3255 _0236_ vssd1 0.647f $ **FLOATING
C3256 a_23299_24349# vssd1 0.508f $ **FLOATING
C3257 a_23119_24349# vssd1 0.604f $ **FLOATING
C3258 cal_lut\[61\] vssd1 1.41f $ **FLOATING
C3259 _0469_ vssd1 4.16f $ **FLOATING
C3260 cal_lut\[31\] vssd1 2.24f $ **FLOATING
C3261 _0468_ vssd1 6.47f $ **FLOATING
C3262 a_22503_24135# vssd1 0.804f $ **FLOATING
C3263 a_19333_24135# vssd1 0.502f $ **FLOATING
C3264 a_18187_24349# vssd1 0.609f $ **FLOATING
C3265 a_18355_24251# vssd1 0.817f $ **FLOATING
C3266 a_17762_24349# vssd1 0.626f $ **FLOATING
C3267 a_17930_24095# vssd1 0.581f $ **FLOATING
C3268 a_17489_23983# vssd1 1.43f $ **FLOATING
C3269 _0082_ vssd1 0.954f $ **FLOATING
C3270 a_17323_23983# vssd1 1.81f $ **FLOATING
C3271 _0481_ vssd1 20.4f $ **FLOATING
C3272 _0645_ vssd1 1.06f $ **FLOATING
C3273 _0094_ vssd1 1.23f $ **FLOATING
C3274 _0009_ vssd1 1.08f $ **FLOATING
C3275 a_12097_23983# vssd1 0.441f $ **FLOATING
C3276 a_11142_23983# vssd1 0.285f $ **FLOATING
C3277 a_12265_24233# vssd1 0.386f $ **FLOATING
C3278 a_11142_24233# vssd1 0.507f $ **FLOATING
C3279 a_10699_24233# vssd1 0.323f $ **FLOATING
C3280 a_10229_24233# vssd1 0.206f $ **FLOATING
C3281 a_9678_24233# vssd1 0.218f $ **FLOATING
C3282 _0765_ vssd1 2.86f $ **FLOATING
C3283 a_7079_24233# vssd1 0.245f $ **FLOATING
C3284 a_6277_24233# vssd1 0.238f $ **FLOATING
C3285 a_5555_24233# vssd1 0.436f $ **FLOATING
C3286 a_5077_24233# vssd1 0.206f $ **FLOATING
C3287 a_3339_23983# vssd1 0.18f $ **FLOATING
C3288 a_4277_23957# vssd1 0.607f $ **FLOATING
C3289 _0822_ vssd1 1.16f $ **FLOATING
C3290 _0411_ vssd1 12.9f $ **FLOATING
C3291 a_1863_24233# vssd1 0.506f $ **FLOATING
C3292 a_15531_24135# vssd1 0.619f $ **FLOATING
C3293 a_14979_24148# vssd1 0.524f $ **FLOATING
C3294 _0849_ vssd1 0.725f $ **FLOATING
C3295 a_13783_24148# vssd1 0.524f $ **FLOATING
C3296 a_13363_24349# vssd1 0.508f $ **FLOATING
C3297 a_13183_24349# vssd1 0.604f $ **FLOATING
C3298 a_11896_24233# vssd1 0.634f $ **FLOATING
C3299 a_10784_23983# vssd1 1.17f $ **FLOATING
C3300 _0707_ vssd1 2.62f $ **FLOATING
C3301 a_10083_24135# vssd1 0.804f $ **FLOATING
C3302 _0712_ vssd1 3.4f $ **FLOATING
C3303 _0723_ vssd1 2.2f $ **FLOATING
C3304 a_9372_24135# vssd1 0.7f $ **FLOATING
C3305 _0752_ vssd1 1.55f $ **FLOATING
C3306 _0797_ vssd1 1.85f $ **FLOATING
C3307 ctr\[5\] vssd1 8.88f $ **FLOATING
C3308 _0429_ vssd1 9.4f $ **FLOATING
C3309 a_4931_24135# vssd1 0.804f $ **FLOATING
C3310 a_3848_24135# vssd1 0.59f $ **FLOATING
C3311 _0804_ vssd1 1.49f $ **FLOATING
C3312 clknet_1_0__leaf_temp1.i_precharge_n vssd1 3.96f $ **FLOATING
C3313 _0823_ vssd1 1f $ **FLOATING
C3314 a_2741_24135# vssd1 0.767f $ **FLOATING
C3315 a_2563_23957# vssd1 0.83f $ **FLOATING
C3316 net22 vssd1 5.34f $ **FLOATING
C3317 _0791_ vssd1 1.78f $ **FLOATING
C3318 a_1464_23957# vssd1 1.22f $ **FLOATING
C3319 _0238_ vssd1 1.08f $ **FLOATING
C3320 a_16761_24527# vssd1 0.206f $ **FLOATING
C3321 a_19609_24527# vssd1 0.23f $ **FLOATING
C3322 _0577_ vssd1 2.33f $ **FLOATING
C3323 _0273_ vssd1 1.01f $ **FLOATING
C3324 a_14365_24527# vssd1 0.23f $ **FLOATING
C3325 a_11547_24847# vssd1 0.279f $ **FLOATING
C3326 a_9223_24527# vssd1 0.253f $ **FLOATING
C3327 a_8397_24527# vssd1 0.203f $ **FLOATING
C3328 a_9967_24847# vssd1 0.211f $ **FLOATING
C3329 a_6565_24527# vssd1 0.191f $ **FLOATING
C3330 a_5645_24527# vssd1 0.191f $ **FLOATING
C3331 _0796_ vssd1 0.909f $ **FLOATING
C3332 a_25003_24833# vssd1 0.604f $ **FLOATING
C3333 cal_lut\[62\] vssd1 2.73f $ **FLOATING
C3334 a_24827_24501# vssd1 0.508f $ **FLOATING
C3335 a_23763_24527# vssd1 0.524f $ **FLOATING
C3336 a_22291_24527# vssd1 0.524f $ **FLOATING
C3337 _0263_ vssd1 0.68f $ **FLOATING
C3338 a_21872_24643# vssd1 0.502f $ **FLOATING
C3339 _0262_ vssd1 0.725f $ **FLOATING
C3340 a_21327_24746# vssd1 0.524f $ **FLOATING
C3341 a_20907_24527# vssd1 0.508f $ **FLOATING
C3342 cal_lut\[84\] vssd1 3.45f $ **FLOATING
C3343 a_20727_24527# vssd1 0.604f $ **FLOATING
C3344 a_20119_24527# vssd1 0.609f $ **FLOATING
C3345 a_20287_24501# vssd1 0.817f $ **FLOATING
C3346 a_19694_24527# vssd1 0.626f $ **FLOATING
C3347 a_19862_24501# vssd1 0.581f $ **FLOATING
C3348 a_19421_24533# vssd1 1.43f $ **FLOATING
C3349 _0083_ vssd1 0.906f $ **FLOATING
C3350 a_19255_24533# vssd1 1.81f $ **FLOATING
C3351 a_18979_24527# vssd1 0.524f $ **FLOATING
C3352 _0261_ vssd1 1.02f $ **FLOATING
C3353 a_17831_24746# vssd1 0.524f $ **FLOATING
C3354 cal_lut\[42\] vssd1 2.67f $ **FLOATING
C3355 a_17401_24759# vssd1 0.502f $ **FLOATING
C3356 a_16679_24527# vssd1 0.804f $ **FLOATING
C3357 a_15711_24833# vssd1 0.604f $ **FLOATING
C3358 cal_lut\[94\] vssd1 1.56f $ **FLOATING
C3359 a_15535_24501# vssd1 0.508f $ **FLOATING
C3360 a_14875_24527# vssd1 0.609f $ **FLOATING
C3361 a_15043_24501# vssd1 0.817f $ **FLOATING
C3362 a_14450_24527# vssd1 0.626f $ **FLOATING
C3363 a_14618_24501# vssd1 0.581f $ **FLOATING
C3364 a_14177_24533# vssd1 1.43f $ **FLOATING
C3365 a_14011_24533# vssd1 1.81f $ **FLOATING
C3366 _0711_ vssd1 2.56f $ **FLOATING
C3367 a_10607_24640# vssd1 0.619f $ **FLOATING
C3368 _0705_ vssd1 4.06f $ **FLOATING
C3369 _0682_ vssd1 2.35f $ **FLOATING
C3370 _0681_ vssd1 3.07f $ **FLOATING
C3371 _0726_ vssd1 1.53f $ **FLOATING
C3372 a_9831_24501# vssd1 0.791f $ **FLOATING
C3373 _0725_ vssd1 1.34f $ **FLOATING
C3374 _0727_ vssd1 0.868f $ **FLOATING
C3375 a_9005_24501# vssd1 0.55f $ **FLOATING
C3376 a_8268_24501# vssd1 0.655f $ **FLOATING
C3377 a_7523_24833# vssd1 0.604f $ **FLOATING
C3378 a_7347_24501# vssd1 0.508f $ **FLOATING
C3379 _0437_ vssd1 8.63f $ **FLOATING
C3380 a_6428_24501# vssd1 0.847f $ **FLOATING
C3381 _0431_ vssd1 7.24f $ **FLOATING
C3382 _0793_ vssd1 0.843f $ **FLOATING
C3383 _0794_ vssd1 3.07f $ **FLOATING
C3384 a_5508_24501# vssd1 0.847f $ **FLOATING
C3385 a_5013_24825# vssd1 0.607f $ **FLOATING
C3386 _0798_ vssd1 1.13f $ **FLOATING
C3387 a_4584_24759# vssd1 0.59f $ **FLOATING
C3388 a_2778_24527# vssd1 4.03f $ **FLOATING
C3389 _0412_ vssd1 7.83f $ **FLOATING
C3390 _0415_ vssd1 1.39f $ **FLOATING
C3391 temp1.i_precharge_n vssd1 1.54f $ **FLOATING
C3392 a_2010_24759# vssd1 0.759f $ **FLOATING
C3393 a_1683_24527# vssd1 0.524f $ **FLOATING
C3394 _0416_ vssd1 0.745f $ **FLOATING
C3395 a_24761_25071# vssd1 0.23f $ **FLOATING
C3396 a_25271_25437# vssd1 0.609f $ **FLOATING
C3397 a_25439_25339# vssd1 0.817f $ **FLOATING
C3398 a_24846_25437# vssd1 0.626f $ **FLOATING
C3399 a_25014_25183# vssd1 0.581f $ **FLOATING
C3400 a_24573_25071# vssd1 1.43f $ **FLOATING
C3401 _0086_ vssd1 1.22f $ **FLOATING
C3402 a_24407_25071# vssd1 1.81f $ **FLOATING
C3403 _0264_ vssd1 0.863f $ **FLOATING
C3404 a_22553_25071# vssd1 0.23f $ **FLOATING
C3405 _0237_ vssd1 24.6f $ **FLOATING
C3406 a_23899_25045# vssd1 0.604f $ **FLOATING
C3407 cal_lut\[86\] vssd1 1.87f $ **FLOATING
C3408 a_23723_25045# vssd1 0.508f $ **FLOATING
C3409 a_23063_25437# vssd1 0.609f $ **FLOATING
C3410 a_23231_25339# vssd1 0.817f $ **FLOATING
C3411 a_22638_25437# vssd1 0.626f $ **FLOATING
C3412 a_22806_25183# vssd1 0.581f $ **FLOATING
C3413 a_22365_25071# vssd1 1.43f $ **FLOATING
C3414 _0085_ vssd1 0.908f $ **FLOATING
C3415 a_22199_25071# vssd1 1.81f $ **FLOATING
C3416 cal_lut\[85\] vssd1 2.08f $ **FLOATING
C3417 a_21081_25071# vssd1 0.23f $ **FLOATING
C3418 a_21591_25437# vssd1 0.609f $ **FLOATING
C3419 a_21759_25339# vssd1 0.817f $ **FLOATING
C3420 a_21166_25437# vssd1 0.626f $ **FLOATING
C3421 a_21334_25183# vssd1 0.581f $ **FLOATING
C3422 a_20893_25071# vssd1 1.43f $ **FLOATING
C3423 _0084_ vssd1 1.03f $ **FLOATING
C3424 a_20727_25071# vssd1 1.81f $ **FLOATING
C3425 cal_lut\[47\] vssd1 2.01f $ **FLOATING
C3426 a_17677_25071# vssd1 0.23f $ **FLOATING
C3427 a_19333_25223# vssd1 0.502f $ **FLOATING
C3428 a_18187_25437# vssd1 0.609f $ **FLOATING
C3429 a_18355_25339# vssd1 0.817f $ **FLOATING
C3430 a_17762_25437# vssd1 0.626f $ **FLOATING
C3431 a_17930_25183# vssd1 0.581f $ **FLOATING
C3432 a_17489_25071# vssd1 1.43f $ **FLOATING
C3433 _0046_ vssd1 0.994f $ **FLOATING
C3434 a_17323_25071# vssd1 1.81f $ **FLOATING
C3435 _0220_ vssd1 1.21f $ **FLOATING
C3436 _0872_ vssd1 16f $ **FLOATING
C3437 cal_lut\[46\] vssd1 1.22f $ **FLOATING
C3438 a_15745_25071# vssd1 0.23f $ **FLOATING
C3439 a_16904_25321# vssd1 0.502f $ **FLOATING
C3440 a_16255_25437# vssd1 0.609f $ **FLOATING
C3441 a_16423_25339# vssd1 0.817f $ **FLOATING
C3442 a_15830_25437# vssd1 0.626f $ **FLOATING
C3443 a_15998_25183# vssd1 0.581f $ **FLOATING
C3444 a_15557_25071# vssd1 1.43f $ **FLOATING
C3445 a_15391_25071# vssd1 1.81f $ **FLOATING
C3446 _0093_ vssd1 1.07f $ **FLOATING
C3447 cal_lut\[9\] vssd1 2.33f $ **FLOATING
C3448 a_11797_25071# vssd1 0.171f $ **FLOATING
C3449 a_10883_25071# vssd1 0.291f $ **FLOATING
C3450 a_10347_25071# vssd1 0.33f $ **FLOATING
C3451 a_9431_25071# vssd1 0.19f $ **FLOATING
C3452 a_9235_25071# vssd1 0.165f $ **FLOATING
C3453 a_8419_25071# vssd1 0.253f $ **FLOATING
C3454 a_8229_25071# vssd1 0.162f $ **FLOATING
C3455 a_12893_25071# vssd1 0.23f $ **FLOATING
C3456 _0272_ vssd1 0.725f $ **FLOATING
C3457 a_14703_25236# vssd1 0.524f $ **FLOATING
C3458 a_14283_25437# vssd1 0.508f $ **FLOATING
C3459 a_14103_25437# vssd1 0.604f $ **FLOATING
C3460 a_13403_25437# vssd1 0.609f $ **FLOATING
C3461 a_13571_25339# vssd1 0.817f $ **FLOATING
C3462 a_12978_25437# vssd1 0.626f $ **FLOATING
C3463 a_13146_25183# vssd1 0.581f $ **FLOATING
C3464 a_12705_25071# vssd1 1.43f $ **FLOATING
C3465 a_12539_25071# vssd1 1.81f $ **FLOATING
C3466 a_8951_25321# vssd1 0.609f $ **FLOATING
C3467 a_8055_25321# vssd1 0.526f $ **FLOATING
C3468 a_7755_25321# vssd1 0.286f $ **FLOATING
C3469 a_7289_25321# vssd1 0.318f $ **FLOATING
C3470 _0735_ vssd1 2.45f $ **FLOATING
C3471 a_6381_25321# vssd1 0.191f $ **FLOATING
C3472 _0795_ vssd1 0.971f $ **FLOATING
C3473 a_4069_25071# vssd1 0.171f $ **FLOATING
C3474 a_2959_25071# vssd1 0.319f $ **FLOATING
C3475 a_5105_25045# vssd1 0.607f $ **FLOATING
C3476 _0827_ vssd1 2.33f $ **FLOATING
C3477 _0747_ vssd1 6.87f $ **FLOATING
C3478 _0706_ vssd1 3.2f $ **FLOATING
C3479 _0730_ vssd1 0.98f $ **FLOATING
C3480 _0708_ vssd1 2.33f $ **FLOATING
C3481 a_11579_25045# vssd1 0.546f $ **FLOATING
C3482 _0731_ vssd1 1.5f $ **FLOATING
C3483 _0729_ vssd1 2.03f $ **FLOATING
C3484 a_10197_25223# vssd1 0.722f $ **FLOATING
C3485 _0714_ vssd1 3.92f $ **FLOATING
C3486 _0713_ vssd1 2.9f $ **FLOATING
C3487 a_7071_25045# vssd1 0.526f $ **FLOATING
C3488 _0805_ vssd1 4.58f $ **FLOATING
C3489 _0751_ vssd1 2f $ **FLOATING
C3490 a_6244_25045# vssd1 0.847f $ **FLOATING
C3491 _0737_ vssd1 7.15f $ **FLOATING
C3492 a_4676_25223# vssd1 0.59f $ **FLOATING
C3493 net21 vssd1 6.66f $ **FLOATING
C3494 _0799_ vssd1 1.02f $ **FLOATING
C3495 a_3851_25045# vssd1 0.546f $ **FLOATING
C3496 _0806_ vssd1 1.24f $ **FLOATING
C3497 _0803_ vssd1 1.06f $ **FLOATING
C3498 _0807_ vssd1 2.1f $ **FLOATING
C3499 a_2564_25045# vssd1 1.33f $ **FLOATING
C3500 a_19149_25615# vssd1 0.23f $ **FLOATING
C3501 a_7853_25615# vssd1 0.191f $ **FLOATING
C3502 a_7291_25615# vssd1 0.253f $ **FLOATING
C3503 _0008_ vssd1 1.02f $ **FLOATING
C3504 _0732_ vssd1 1.35f $ **FLOATING
C3505 a_9773_25935# vssd1 0.171f $ **FLOATING
C3506 _0721_ vssd1 2.74f $ **FLOATING
C3507 _0750_ vssd1 4.48f $ **FLOATING
C3508 _0792_ vssd1 1.68f $ **FLOATING
C3509 _0802_ vssd1 1.35f $ **FLOATING
C3510 a_2887_25615# vssd1 0.436f $ **FLOATING
C3511 a_2366_25615# vssd1 0.333f $ **FLOATING
C3512 a_4811_25935# vssd1 0.171f $ **FLOATING
C3513 a_3656_25847# vssd1 0.525f $ **FLOATING
C3514 temp1.dcdel_capnode_notouch_ vssd1 8.33f $ **FLOATING
C3515 a_21872_25731# vssd1 0.502f $ **FLOATING
C3516 cal_lut\[87\] vssd1 4.88f $ **FLOATING
C3517 a_21279_25615# vssd1 0.524f $ **FLOATING
C3518 _0265_ vssd1 1.06f $ **FLOATING
C3519 a_19659_25615# vssd1 0.609f $ **FLOATING
C3520 a_19827_25589# vssd1 0.817f $ **FLOATING
C3521 a_19234_25615# vssd1 0.626f $ **FLOATING
C3522 a_19402_25589# vssd1 0.581f $ **FLOATING
C3523 a_18961_25621# vssd1 1.43f $ **FLOATING
C3524 _0047_ vssd1 0.872f $ **FLOATING
C3525 a_18795_25621# vssd1 1.81f $ **FLOATING
C3526 a_18519_25615# vssd1 0.524f $ **FLOATING
C3527 _0221_ vssd1 1.23f $ **FLOATING
C3528 a_18111_25589# vssd1 0.698f $ **FLOATING
C3529 a_17135_25615# vssd1 0.508f $ **FLOATING
C3530 a_16955_25615# vssd1 0.604f $ **FLOATING
C3531 a_16219_25623# vssd1 0.648f $ **FLOATING
C3532 a_15904_25589# vssd1 0.648f $ **FLOATING
C3533 a_15479_25615# vssd1 0.508f $ **FLOATING
C3534 a_15299_25615# vssd1 0.604f $ **FLOATING
C3535 a_12955_25834# vssd1 0.524f $ **FLOATING
C3536 _0718_ vssd1 3.55f $ **FLOATING
C3537 _0715_ vssd1 3.48f $ **FLOATING
C3538 _0719_ vssd1 0.739f $ **FLOATING
C3539 _0720_ vssd1 7.66f $ **FLOATING
C3540 a_9555_25847# vssd1 0.546f $ **FLOATING
C3541 _0734_ vssd1 1.9f $ **FLOATING
C3542 _0749_ vssd1 2.06f $ **FLOATING
C3543 _0748_ vssd1 4.46f $ **FLOATING
C3544 _0728_ vssd1 4.83f $ **FLOATING
C3545 a_7716_25589# vssd1 0.847f $ **FLOATING
C3546 _0724_ vssd1 6.53f $ **FLOATING
C3547 _0722_ vssd1 3f $ **FLOATING
C3548 _0733_ vssd1 2.71f $ **FLOATING
C3549 a_7073_25589# vssd1 0.55f $ **FLOATING
C3550 a_4984_25615# vssd1 0.546f $ **FLOATING
C3551 a_4461_25913# vssd1 0.607f $ **FLOATING
C3552 _0828_ vssd1 1.27f $ **FLOATING
C3553 _0759_ vssd1 9.32f $ **FLOATING
C3554 a_4032_25847# vssd1 0.59f $ **FLOATING
C3555 ctr\[3\] vssd1 10.4f $ **FLOATING
C3556 a_2209_25589# vssd1 0.723f $ **FLOATING
C3557 a_23395_26159# vssd1 0.524f $ **FLOATING
C3558 a_21709_26159# vssd1 0.23f $ **FLOATING
C3559 cal_lut\[88\] vssd1 4.02f $ **FLOATING
C3560 a_17861_26159# vssd1 0.23f $ **FLOATING
C3561 _0087_ vssd1 1.07f $ **FLOATING
C3562 a_21291_26159# vssd1 0.581f $ **FLOATING
C3563 a_21362_26133# vssd1 0.626f $ **FLOATING
C3564 a_21155_26133# vssd1 1.81f $ **FLOATING
C3565 a_21162_26433# vssd1 1.43f $ **FLOATING
C3566 a_20871_26133# vssd1 0.609f $ **FLOATING
C3567 a_20775_26311# vssd1 0.817f $ **FLOATING
C3568 a_19531_26159# vssd1 0.524f $ **FLOATING
C3569 a_18371_26525# vssd1 0.609f $ **FLOATING
C3570 a_18539_26427# vssd1 0.817f $ **FLOATING
C3571 a_17946_26525# vssd1 0.626f $ **FLOATING
C3572 a_18114_26271# vssd1 0.581f $ **FLOATING
C3573 a_17673_26159# vssd1 1.43f $ **FLOATING
C3574 a_17507_26159# vssd1 1.81f $ **FLOATING
C3575 _0088_ vssd1 0.906f $ **FLOATING
C3576 _0045_ vssd1 1.23f $ **FLOATING
C3577 _0848_ vssd1 0.902f $ **FLOATING
C3578 a_6377_26409# vssd1 0.253f $ **FLOATING
C3579 a_5801_26409# vssd1 0.329f $ **FLOATING
C3580 a_5547_26409# vssd1 0.381f $ **FLOATING
C3581 ctr\[1\] vssd1 13.6f $ **FLOATING
C3582 _0410_ vssd1 9.04f $ **FLOATING
C3583 a_17231_26159# vssd1 0.524f $ **FLOATING
C3584 _0267_ vssd1 0.895f $ **FLOATING
C3585 _0215_ vssd1 1.6f $ **FLOATING
C3586 a_16635_26324# vssd1 0.524f $ **FLOATING
C3587 _0219_ vssd1 0.81f $ **FLOATING
C3588 a_15623_26324# vssd1 0.524f $ **FLOATING
C3589 a_12995_26525# vssd1 0.508f $ **FLOATING
C3590 a_12815_26525# vssd1 0.604f $ **FLOATING
C3591 a_12443_26525# vssd1 0.508f $ **FLOATING
C3592 a_12263_26525# vssd1 0.604f $ **FLOATING
C3593 _0841_ vssd1 20f $ **FLOATING
C3594 _0846_ vssd1 3.97f $ **FLOATING
C3595 a_12035_26324# vssd1 0.524f $ **FLOATING
C3596 a_9559_26481# vssd1 0.83f $ **FLOATING
C3597 a_9319_26159# vssd1 0.767f $ **FLOATING
C3598 a_6546_26159# vssd1 0.55f $ **FLOATING
C3599 _0399_ vssd1 0.906f $ **FLOATING
C3600 a_3991_26409# vssd1 0.436f $ **FLOATING
C3601 clknet_1_1__leaf_temp1.i_precharge_n vssd1 3.27f $ **FLOATING
C3602 a_4678_26311# vssd1 0.759f $ **FLOATING
C3603 _0418_ vssd1 14.3f $ **FLOATING
C3604 clknet_0_temp1.i_precharge_n vssd1 5.63f $ **FLOATING
C3605 a_1753_26133# vssd1 4.03f $ **FLOATING
C3606 a_24101_27081# vssd1 0.23f $ **FLOATING
C3607 cal_lut\[57\] vssd1 3.62f $ **FLOATING
C3608 _0231_ vssd1 1.01f $ **FLOATING
C3609 a_16845_26703# vssd1 0.214f $ **FLOATING
C3610 a_16761_26703# vssd1 0.167f $ **FLOATING
C3611 a_19793_26703# vssd1 0.23f $ **FLOATING
C3612 _0227_ vssd1 1.15f $ **FLOATING
C3613 _0691_ vssd1 7.17f $ **FLOATING
C3614 cal_lut\[93\] vssd1 3.31f $ **FLOATING
C3615 a_13905_26703# vssd1 0.23f $ **FLOATING
C3616 a_10423_26703# vssd1 0.388f $ **FLOATING
C3617 a_12065_26703# vssd1 0.23f $ **FLOATING
C3618 _0592_ vssd1 4.04f $ **FLOATING
C3619 _0056_ vssd1 1.25f $ **FLOATING
C3620 a_23683_27081# vssd1 0.581f $ **FLOATING
C3621 a_23754_26980# vssd1 0.626f $ **FLOATING
C3622 a_23554_26825# vssd1 1.43f $ **FLOATING
C3623 a_23547_26921# vssd1 1.81f $ **FLOATING
C3624 a_23263_26935# vssd1 0.609f $ **FLOATING
C3625 a_23167_26935# vssd1 0.817f $ **FLOATING
C3626 a_22747_26703# vssd1 0.508f $ **FLOATING
C3627 a_22567_26703# vssd1 0.604f $ **FLOATING
C3628 a_20303_26703# vssd1 0.609f $ **FLOATING
C3629 a_20471_26677# vssd1 0.817f $ **FLOATING
C3630 a_19878_26703# vssd1 0.626f $ **FLOATING
C3631 a_20046_26677# vssd1 0.581f $ **FLOATING
C3632 a_19605_26709# vssd1 1.43f $ **FLOATING
C3633 _0052_ vssd1 0.961f $ **FLOATING
C3634 a_19439_26709# vssd1 1.81f $ **FLOATING
C3635 a_19057_26935# vssd1 0.502f $ **FLOATING
C3636 a_16679_26703# vssd1 0.972f $ **FLOATING
C3637 a_15469_26935# vssd1 0.502f $ **FLOATING
C3638 a_14415_26703# vssd1 0.609f $ **FLOATING
C3639 a_14583_26677# vssd1 0.817f $ **FLOATING
C3640 a_13990_26703# vssd1 0.626f $ **FLOATING
C3641 a_14158_26677# vssd1 0.581f $ **FLOATING
C3642 a_13717_26709# vssd1 1.43f $ **FLOATING
C3643 _0092_ vssd1 0.872f $ **FLOATING
C3644 a_13551_26709# vssd1 1.81f $ **FLOATING
C3645 net48 vssd1 13.7f $ **FLOATING
C3646 a_13275_26703# vssd1 0.524f $ **FLOATING
C3647 a_12575_26703# vssd1 0.609f $ **FLOATING
C3648 a_12743_26677# vssd1 0.817f $ **FLOATING
C3649 a_12150_26703# vssd1 0.626f $ **FLOATING
C3650 a_12318_26677# vssd1 0.581f $ **FLOATING
C3651 a_11877_26709# vssd1 1.43f $ **FLOATING
C3652 _0006_ vssd1 0.961f $ **FLOATING
C3653 a_11711_26709# vssd1 1.81f $ **FLOATING
C3654 _0385_ vssd1 0.907f $ **FLOATING
C3655 a_9835_26703# vssd1 0.83f $ **FLOATING
C3656 a_9595_26703# vssd1 0.767f $ **FLOATING
C3657 _0460_ vssd1 26.8f $ **FLOATING
C3658 ctr\[6\] vssd1 11.3f $ **FLOATING
C3659 clknet_1_1__leaf__0380_ vssd1 8f $ **FLOATING
C3660 _0409_ vssd1 1.63f $ **FLOATING
C3661 net76 vssd1 0.868f $ **FLOATING
C3662 _0400_ vssd1 0.935f $ **FLOATING
C3663 a_3171_26703# vssd1 0.388f $ **FLOATING
C3664 a_2327_26703# vssd1 0.525f $ **FLOATING
C3665 a_2000_26935# vssd1 0.525f $ **FLOATING
C3666 a_1407_26703# vssd1 0.525f $ **FLOATING
C3667 a_7618_26935# vssd1 0.702f $ **FLOATING
C3668 a_6739_26703# vssd1 0.553f $ **FLOATING
C3669 a_6633_26703# vssd1 0.794f $ **FLOATING
C3670 a_6397_26703# vssd1 0.788f $ **FLOATING
C3671 a_5864_26819# vssd1 0.502f $ **FLOATING
C3672 a_5227_26935# vssd1 0.619f $ **FLOATING
C3673 _0414_ vssd1 11.6f $ **FLOATING
C3674 _0746_ vssd1 4.42f $ **FLOATING
C3675 a_23811_27412# vssd1 0.524f $ **FLOATING
C3676 a_23273_27247# vssd1 0.23f $ **FLOATING
C3677 cal_lut\[56\] vssd1 3.08f $ **FLOATING
C3678 _0230_ vssd1 1.41f $ **FLOATING
C3679 cal_lut\[53\] vssd1 4.77f $ **FLOATING
C3680 cal_lut\[48\] vssd1 2.75f $ **FLOATING
C3681 _0222_ vssd1 11.5f $ **FLOATING
C3682 cal_lut\[89\] vssd1 3.25f $ **FLOATING
C3683 a_16481_27247# vssd1 0.23f $ **FLOATING
C3684 _0055_ vssd1 0.872f $ **FLOATING
C3685 a_22855_27247# vssd1 0.581f $ **FLOATING
C3686 a_22926_27221# vssd1 0.626f $ **FLOATING
C3687 a_22719_27221# vssd1 1.81f $ **FLOATING
C3688 a_22726_27521# vssd1 1.43f $ **FLOATING
C3689 a_22435_27221# vssd1 0.609f $ **FLOATING
C3690 a_22339_27399# vssd1 0.817f $ **FLOATING
C3691 a_21919_27613# vssd1 0.508f $ **FLOATING
C3692 a_21739_27613# vssd1 0.604f $ **FLOATING
C3693 a_21136_27497# vssd1 0.502f $ **FLOATING
C3694 _0228_ vssd1 0.758f $ **FLOATING
C3695 a_20775_27412# vssd1 0.524f $ **FLOATING
C3696 a_20308_27497# vssd1 0.502f $ **FLOATING
C3697 a_19664_27497# vssd1 0.502f $ **FLOATING
C3698 a_18560_27497# vssd1 0.502f $ **FLOATING
C3699 a_17871_27613# vssd1 0.508f $ **FLOATING
C3700 a_17691_27613# vssd1 0.604f $ **FLOATING
C3701 _0266_ vssd1 18.3f $ **FLOATING
C3702 a_16991_27613# vssd1 0.609f $ **FLOATING
C3703 a_17159_27515# vssd1 0.817f $ **FLOATING
C3704 a_16566_27613# vssd1 0.626f $ **FLOATING
C3705 a_16734_27359# vssd1 0.581f $ **FLOATING
C3706 a_16293_27247# vssd1 1.43f $ **FLOATING
C3707 _0042_ vssd1 1.21f $ **FLOATING
C3708 a_16127_27247# vssd1 1.81f $ **FLOATING
C3709 _0489_ vssd1 7.06f $ **FLOATING
C3710 a_15557_27497# vssd1 0.214f $ **FLOATING
C3711 a_15473_27497# vssd1 0.167f $ **FLOATING
C3712 _0690_ vssd1 1.36f $ **FLOATING
C3713 a_14829_27497# vssd1 0.206f $ **FLOATING
C3714 a_14185_27497# vssd1 0.206f $ **FLOATING
C3715 a_12709_27247# vssd1 0.23f $ **FLOATING
C3716 a_15391_27247# vssd1 0.972f $ **FLOATING
C3717 _0482_ vssd1 3.76f $ **FLOATING
C3718 _0484_ vssd1 7.36f $ **FLOATING
C3719 _0488_ vssd1 0.896f $ **FLOATING
C3720 a_14747_27497# vssd1 0.804f $ **FLOATING
C3721 cal_lut\[7\] vssd1 2.46f $ **FLOATING
C3722 a_14103_27497# vssd1 0.804f $ **FLOATING
C3723 _0486_ vssd1 6.61f $ **FLOATING
C3724 _0487_ vssd1 10.6f $ **FLOATING
C3725 cal_lut\[8\] vssd1 1.83f $ **FLOATING
C3726 a_13219_27613# vssd1 0.609f $ **FLOATING
C3727 a_13387_27515# vssd1 0.817f $ **FLOATING
C3728 a_12794_27613# vssd1 0.626f $ **FLOATING
C3729 a_12962_27359# vssd1 0.581f $ **FLOATING
C3730 a_12521_27247# vssd1 1.43f $ **FLOATING
C3731 a_12355_27247# vssd1 1.81f $ **FLOATING
C3732 a_10777_27247# vssd1 0.216f $ **FLOATING
C3733 a_11287_27613# vssd1 0.599f $ **FLOATING
C3734 a_11458_27500# vssd1 1.41f $ **FLOATING
C3735 a_10871_27613# vssd1 0.627f $ **FLOATING
C3736 a_11030_27383# vssd1 0.587f $ **FLOATING
C3737 a_10589_27247# vssd1 1.39f $ **FLOATING
C3738 _0196_ vssd1 1.06f $ **FLOATING
C3739 a_10423_27247# vssd1 1.77f $ **FLOATING
C3740 a_7281_27247# vssd1 0.23f $ **FLOATING
C3741 a_4897_27247# vssd1 0.21f $ **FLOATING
C3742 a_9096_27221# vssd1 0.648f $ **FLOATING
C3743 a_7791_27613# vssd1 0.609f $ **FLOATING
C3744 a_7959_27515# vssd1 0.97f $ **FLOATING
C3745 a_7366_27613# vssd1 0.626f $ **FLOATING
C3746 a_7534_27359# vssd1 0.581f $ **FLOATING
C3747 a_7093_27247# vssd1 1.43f $ **FLOATING
C3748 a_6927_27247# vssd1 1.81f $ **FLOATING
C3749 a_6437_27247# vssd1 0.23f $ **FLOATING
C3750 _0206_ vssd1 1.23f $ **FLOATING
C3751 a_6019_27247# vssd1 0.581f $ **FLOATING
C3752 a_6090_27221# vssd1 0.626f $ **FLOATING
C3753 a_5883_27221# vssd1 1.81f $ **FLOATING
C3754 a_5890_27521# vssd1 1.43f $ **FLOATING
C3755 a_5599_27221# vssd1 0.609f $ **FLOATING
C3756 a_5503_27399# vssd1 0.817f $ **FLOATING
C3757 a_4705_27552# vssd1 0.446f $ **FLOATING
C3758 a_4277_27221# vssd1 0.607f $ **FLOATING
C3759 _0829_ vssd1 1.59f $ **FLOATING
C3760 _0424_ vssd1 9.02f $ **FLOATING
C3761 a_3848_27399# vssd1 0.59f $ **FLOATING
C3762 _0830_ vssd1 0.883f $ **FLOATING
C3763 a_3017_27399# vssd1 0.767f $ **FLOATING
C3764 a_2839_27221# vssd1 0.83f $ **FLOATING
C3765 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 2.42f $ **FLOATING
C3766 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd vssd1 1.9f $ **FLOATING
C3767 a_1775_27247# vssd1 0.525f $ **FLOATING
C3768 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 2.08f $ **FLOATING
C3769 cal_lut\[55\] vssd1 3.78f $ **FLOATING
C3770 a_22185_27791# vssd1 0.23f $ **FLOATING
C3771 cal_lut\[54\] vssd1 4.22f $ **FLOATING
C3772 a_20621_27791# vssd1 0.23f $ **FLOATING
C3773 a_18489_28169# vssd1 0.23f $ **FLOATING
C3774 cal_lut\[91\] vssd1 2.15f $ **FLOATING
C3775 a_15009_27791# vssd1 0.23f $ **FLOATING
C3776 a_9779_27791# vssd1 0.388f $ **FLOATING
C3777 _0271_ vssd1 1.37f $ **FLOATING
C3778 _0007_ vssd1 0.975f $ **FLOATING
C3779 a_6745_27791# vssd1 0.253f $ **FLOATING
C3780 _0816_ vssd1 0.916f $ **FLOATING
C3781 a_5639_27791# vssd1 0.238f $ **FLOATING
C3782 _0212_ vssd1 0.994f $ **FLOATING
C3783 _0401_ vssd1 1.3f $ **FLOATING
C3784 a_4521_27791# vssd1 0.23f $ **FLOATING
C3785 net70 vssd1 1.01f $ **FLOATING
C3786 a_2879_27791# vssd1 0.525f $ **FLOATING
C3787 a_22695_27791# vssd1 0.609f $ **FLOATING
C3788 a_22863_27765# vssd1 0.817f $ **FLOATING
C3789 a_22270_27791# vssd1 0.626f $ **FLOATING
C3790 a_22438_27765# vssd1 0.581f $ **FLOATING
C3791 a_21997_27797# vssd1 1.43f $ **FLOATING
C3792 a_21831_27797# vssd1 1.81f $ **FLOATING
C3793 net47 vssd1 11.8f $ **FLOATING
C3794 a_21131_27791# vssd1 0.609f $ **FLOATING
C3795 a_21299_27765# vssd1 0.817f $ **FLOATING
C3796 a_20706_27791# vssd1 0.626f $ **FLOATING
C3797 a_20874_27765# vssd1 0.581f $ **FLOATING
C3798 a_20433_27797# vssd1 1.43f $ **FLOATING
C3799 _0053_ vssd1 1.07f $ **FLOATING
C3800 a_20267_27797# vssd1 1.81f $ **FLOATING
C3801 _0223_ vssd1 0.947f $ **FLOATING
C3802 a_19763_28010# vssd1 0.524f $ **FLOATING
C3803 a_18979_27791# vssd1 0.524f $ **FLOATING
C3804 _0268_ vssd1 0.947f $ **FLOATING
C3805 a_18071_28169# vssd1 0.581f $ **FLOATING
C3806 a_18142_28068# vssd1 0.626f $ **FLOATING
C3807 a_17942_27913# vssd1 1.43f $ **FLOATING
C3808 a_17935_28009# vssd1 1.81f $ **FLOATING
C3809 a_17651_28023# vssd1 0.609f $ **FLOATING
C3810 a_17555_28023# vssd1 0.817f $ **FLOATING
C3811 a_15519_27791# vssd1 0.609f $ **FLOATING
C3812 a_15687_27765# vssd1 0.817f $ **FLOATING
C3813 a_15094_27791# vssd1 0.626f $ **FLOATING
C3814 a_15262_27765# vssd1 0.581f $ **FLOATING
C3815 a_14821_27797# vssd1 1.43f $ **FLOATING
C3816 a_14655_27797# vssd1 1.81f $ **FLOATING
C3817 net41 vssd1 14.9f $ **FLOATING
C3818 _0260_ vssd1 20.6f $ **FLOATING
C3819 cal_lut\[92\] vssd1 2f $ **FLOATING
C3820 a_13997_28023# vssd1 0.502f $ **FLOATING
C3821 _0847_ vssd1 1.31f $ **FLOATING
C3822 a_12679_28010# vssd1 0.524f $ **FLOATING
C3823 _0386_ vssd1 1.37f $ **FLOATING
C3824 a_9275_28023# vssd1 0.619f $ **FLOATING
C3825 dec1.i_ones vssd1 8.76f $ **FLOATING
C3826 a_8845_28023# vssd1 0.502f $ **FLOATING
C3827 a_6914_28111# vssd1 0.55f $ **FLOATING
C3828 _0826_ vssd1 2.91f $ **FLOATING
C3829 _0408_ vssd1 1.66f $ **FLOATING
C3830 ctr\[7\] vssd1 7.67f $ **FLOATING
C3831 _0811_ vssd1 9.22f $ **FLOATING
C3832 a_5031_27791# vssd1 0.609f $ **FLOATING
C3833 a_5199_27765# vssd1 0.817f $ **FLOATING
C3834 a_4606_27791# vssd1 0.626f $ **FLOATING
C3835 a_4774_27765# vssd1 0.581f $ **FLOATING
C3836 a_4333_27797# vssd1 1.43f $ **FLOATING
C3837 _0207_ vssd1 1.23f $ **FLOATING
C3838 a_4167_27797# vssd1 1.81f $ **FLOATING
C3839 clknet_1_1__leaf_net67 vssd1 7.77f $ **FLOATING
C3840 _0744_ vssd1 11.5f $ **FLOATING
C3841 _0824_ vssd1 2.41f $ **FLOATING
C3842 a_1913_28023# vssd1 0.767f $ **FLOATING
C3843 a_1735_27765# vssd1 0.83f $ **FLOATING
C3844 _0054_ vssd1 1.09f $ **FLOATING
C3845 cal_lut\[90\] vssd1 4.58f $ **FLOATING
C3846 a_19609_28335# vssd1 0.23f $ **FLOATING
C3847 a_21463_28335# vssd1 0.524f $ **FLOATING
C3848 _0229_ vssd1 1.09f $ **FLOATING
C3849 a_20119_28701# vssd1 0.609f $ **FLOATING
C3850 a_20287_28603# vssd1 0.817f $ **FLOATING
C3851 a_19694_28701# vssd1 0.626f $ **FLOATING
C3852 a_19862_28447# vssd1 0.581f $ **FLOATING
C3853 a_19421_28335# vssd1 1.43f $ **FLOATING
C3854 _0089_ vssd1 1.06f $ **FLOATING
C3855 a_19255_28335# vssd1 1.81f $ **FLOATING
C3856 _0090_ vssd1 1.16f $ **FLOATING
C3857 _0091_ vssd1 1.04f $ **FLOATING
C3858 a_10685_28335# vssd1 0.216f $ **FLOATING
C3859 a_17875_28335# vssd1 0.524f $ **FLOATING
C3860 _0269_ vssd1 1.15f $ **FLOATING
C3861 a_17415_28335# vssd1 0.524f $ **FLOATING
C3862 a_17047_28335# vssd1 0.524f $ **FLOATING
C3863 _0270_ vssd1 1.3f $ **FLOATING
C3864 a_15255_28500# vssd1 0.524f $ **FLOATING
C3865 a_14747_28335# vssd1 0.524f $ **FLOATING
C3866 _0225_ vssd1 0.647f $ **FLOATING
C3867 a_14375_28701# vssd1 0.508f $ **FLOATING
C3868 a_14195_28701# vssd1 0.604f $ **FLOATING
C3869 a_13691_28500# vssd1 0.524f $ **FLOATING
C3870 a_11195_28701# vssd1 0.599f $ **FLOATING
C3871 a_11366_28588# vssd1 1.41f $ **FLOATING
C3872 a_10779_28701# vssd1 0.627f $ **FLOATING
C3873 a_10938_28471# vssd1 0.587f $ **FLOATING
C3874 a_10497_28335# vssd1 1.39f $ **FLOATING
C3875 _0197_ vssd1 1.31f $ **FLOATING
C3876 a_10331_28335# vssd1 1.77f $ **FLOATING
C3877 a_8951_28335# vssd1 0.21f $ **FLOATING
C3878 a_7749_28335# vssd1 0.21f $ **FLOATING
C3879 a_9563_28487# vssd1 0.56f $ **FLOATING
C3880 a_9179_28309# vssd1 0.446f $ **FLOATING
C3881 _0407_ vssd1 0.788f $ **FLOATING
C3882 _0406_ vssd1 1.54f $ **FLOATING
C3883 a_7557_28640# vssd1 0.446f $ **FLOATING
C3884 _0839_ vssd1 14.9f $ **FLOATING
C3885 _0405_ vssd1 0.768f $ **FLOATING
C3886 a_7111_28585# vssd1 0.238f $ **FLOATING
C3887 a_6647_28585# vssd1 0.253f $ **FLOATING
C3888 net74 vssd1 0.957f $ **FLOATING
C3889 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd vssd1 0.968f $ **FLOATING
C3890 a_3081_28309# vssd1 0.607f $ **FLOATING
C3891 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 1.39f $ **FLOATING
C3892 _0403_ vssd1 1.1f $ **FLOATING
C3893 a_6429_28309# vssd1 0.55f $ **FLOATING
C3894 a_6003_28335# vssd1 0.553f $ **FLOATING
C3895 a_5897_28335# vssd1 0.794f $ **FLOATING
C3896 a_5661_28335# vssd1 0.788f $ **FLOATING
C3897 ctr\[8\] vssd1 6.11f $ **FLOATING
C3898 _0419_ vssd1 6.41f $ **FLOATING
C3899 a_2652_28487# vssd1 0.59f $ **FLOATING
C3900 _0832_ vssd1 0.692f $ **FLOATING
C3901 a_2377_28500# vssd1 0.524f $ **FLOATING
C3902 _0825_ vssd1 0.839f $ **FLOATING
C3903 a_1641_28500# vssd1 0.524f $ **FLOATING
C3904 a_19793_28879# vssd1 0.23f $ **FLOATING
C3905 cal_lut\[52\] vssd1 4.6f $ **FLOATING
C3906 a_18137_28879# vssd1 0.23f $ **FLOATING
C3907 _0217_ vssd1 0.922f $ **FLOATING
C3908 _0226_ vssd1 0.973f $ **FLOATING
C3909 cal_lut\[45\] vssd1 3.4f $ **FLOATING
C3910 a_15285_28879# vssd1 0.23f $ **FLOATING
C3911 cal_lut\[50\] vssd1 1.9f $ **FLOATING
C3912 a_13629_28879# vssd1 0.23f $ **FLOATING
C3913 a_10025_29257# vssd1 0.23f $ **FLOATING
C3914 net78 vssd1 0.916f $ **FLOATING
C3915 _0815_ vssd1 2.94f $ **FLOATING
C3916 net73 vssd1 1.13f $ **FLOATING
C3917 net79 vssd1 1.29f $ **FLOATING
C3918 _0812_ vssd1 2.6f $ **FLOATING
C3919 a_5173_29199# vssd1 0.21f $ **FLOATING
C3920 a_20303_28879# vssd1 0.609f $ **FLOATING
C3921 a_20471_28853# vssd1 0.817f $ **FLOATING
C3922 a_19878_28879# vssd1 0.626f $ **FLOATING
C3923 a_20046_28853# vssd1 0.581f $ **FLOATING
C3924 a_19605_28885# vssd1 1.43f $ **FLOATING
C3925 _0048_ vssd1 1.17f $ **FLOATING
C3926 a_19439_28885# vssd1 1.81f $ **FLOATING
C3927 a_18647_28879# vssd1 0.609f $ **FLOATING
C3928 a_18815_28853# vssd1 0.817f $ **FLOATING
C3929 a_18222_28879# vssd1 0.626f $ **FLOATING
C3930 a_18390_28853# vssd1 0.581f $ **FLOATING
C3931 a_17949_28885# vssd1 1.43f $ **FLOATING
C3932 _0051_ vssd1 1.16f $ **FLOATING
C3933 a_17783_28885# vssd1 1.81f $ **FLOATING
C3934 net46 vssd1 7.03f $ **FLOATING
C3935 a_17459_29185# vssd1 0.604f $ **FLOATING
C3936 cal_lut\[43\] vssd1 2.12f $ **FLOATING
C3937 a_17283_28853# vssd1 0.508f $ **FLOATING
C3938 a_16859_28879# vssd1 0.508f $ **FLOATING
C3939 a_16679_28879# vssd1 0.604f $ **FLOATING
C3940 a_15795_28879# vssd1 0.609f $ **FLOATING
C3941 a_15963_28853# vssd1 0.817f $ **FLOATING
C3942 a_15370_28879# vssd1 0.626f $ **FLOATING
C3943 a_15538_28853# vssd1 0.581f $ **FLOATING
C3944 a_15097_28885# vssd1 1.43f $ **FLOATING
C3945 a_14931_28885# vssd1 1.81f $ **FLOATING
C3946 a_14139_28879# vssd1 0.609f $ **FLOATING
C3947 a_14307_28853# vssd1 0.817f $ **FLOATING
C3948 a_13714_28879# vssd1 0.626f $ **FLOATING
C3949 a_13882_28853# vssd1 0.581f $ **FLOATING
C3950 a_13441_28885# vssd1 1.43f $ **FLOATING
C3951 _0049_ vssd1 1.01f $ **FLOATING
C3952 a_13275_28885# vssd1 1.81f $ **FLOATING
C3953 a_11120_28853# vssd1 0.648f $ **FLOATING
C3954 _0211_ vssd1 1.43f $ **FLOATING
C3955 a_9607_29257# vssd1 0.581f $ **FLOATING
C3956 a_9678_29156# vssd1 0.626f $ **FLOATING
C3957 a_9478_29001# vssd1 1.43f $ **FLOATING
C3958 a_9471_29097# vssd1 1.81f $ **FLOATING
C3959 a_9187_29111# vssd1 0.609f $ **FLOATING
C3960 a_9091_29111# vssd1 0.817f $ **FLOATING
C3961 a_8671_28879# vssd1 0.553f $ **FLOATING
C3962 a_8565_28879# vssd1 0.794f $ **FLOATING
C3963 a_8329_28879# vssd1 0.788f $ **FLOATING
C3964 ctr\[12\] vssd1 6.94f $ **FLOATING
C3965 a_7847_28992# vssd1 0.619f $ **FLOATING
C3966 a_7475_28879# vssd1 0.553f $ **FLOATING
C3967 a_7369_28879# vssd1 0.794f $ **FLOATING
C3968 a_7133_28879# vssd1 0.788f $ **FLOATING
C3969 a_6799_28853# vssd1 0.788f $ **FLOATING
C3970 a_6541_28853# vssd1 0.794f $ **FLOATING
C3971 a_6445_29111# vssd1 0.553f $ **FLOATING
C3972 a_5915_28879# vssd1 0.524f $ **FLOATING
C3973 _0813_ vssd1 0.666f $ **FLOATING
C3974 a_5487_29217# vssd1 0.56f $ **FLOATING
C3975 _0402_ vssd1 0.868f $ **FLOATING
C3976 a_4981_28940# vssd1 0.446f $ **FLOATING
C3977 _0390_ vssd1 17.2f $ **FLOATING
C3978 a_2879_28879# vssd1 0.525f $ **FLOATING
C3979 a_2000_29111# vssd1 0.525f $ **FLOATING
C3980 a_4187_28918# vssd1 0.59f $ **FLOATING
C3981 a_3933_28918# vssd1 0.607f $ **FLOATING
C3982 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 1.66f $ **FLOATING
C3983 net45 vssd1 13.3f $ **FLOATING
C3984 a_17845_29423# vssd1 0.23f $ **FLOATING
C3985 cal_lut\[51\] vssd1 4.67f $ **FLOATING
C3986 a_15009_29423# vssd1 0.23f $ **FLOATING
C3987 _0043_ vssd1 1.47f $ **FLOATING
C3988 a_17427_29423# vssd1 0.581f $ **FLOATING
C3989 a_17498_29397# vssd1 0.626f $ **FLOATING
C3990 a_17291_29397# vssd1 1.81f $ **FLOATING
C3991 a_17298_29697# vssd1 1.43f $ **FLOATING
C3992 a_17007_29397# vssd1 0.609f $ **FLOATING
C3993 a_16911_29575# vssd1 0.817f $ **FLOATING
C3994 a_16355_29397# vssd1 0.604f $ **FLOATING
C3995 cal_lut\[44\] vssd1 2.47f $ **FLOATING
C3996 a_16179_29397# vssd1 0.508f $ **FLOATING
C3997 a_15519_29789# vssd1 0.609f $ **FLOATING
C3998 a_15687_29691# vssd1 0.817f $ **FLOATING
C3999 a_15094_29789# vssd1 0.626f $ **FLOATING
C4000 a_15262_29535# vssd1 0.581f $ **FLOATING
C4001 a_14821_29423# vssd1 1.43f $ **FLOATING
C4002 _0050_ vssd1 1.27f $ **FLOATING
C4003 a_14655_29423# vssd1 1.81f $ **FLOATING
C4004 net40 vssd1 10.6f $ **FLOATING
C4005 _0224_ vssd1 1.17f $ **FLOATING
C4006 net71 vssd1 1.78f $ **FLOATING
C4007 a_7741_29423# vssd1 0.23f $ **FLOATING
C4008 _0216_ vssd1 17.7f $ **FLOATING
C4009 a_14331_29397# vssd1 0.604f $ **FLOATING
C4010 cal_lut\[49\] vssd1 5.26f $ **FLOATING
C4011 a_14155_29397# vssd1 0.508f $ **FLOATING
C4012 a_11527_29423# vssd1 0.525f $ **FLOATING
C4013 a_11200_29575# vssd1 0.525f $ **FLOATING
C4014 a_10740_29575# vssd1 0.525f $ **FLOATING
C4015 _0784_ vssd1 8.67f $ **FLOATING
C4016 a_9687_29423# vssd1 0.698f $ **FLOATING
C4017 ctr\[11\] vssd1 6.91f $ **FLOATING
C4018 a_9375_29397# vssd1 0.788f $ **FLOATING
C4019 a_9117_29397# vssd1 0.794f $ **FLOATING
C4020 a_9021_29575# vssd1 0.553f $ **FLOATING
C4021 a_8251_29789# vssd1 0.609f $ **FLOATING
C4022 a_8419_29691# vssd1 0.817f $ **FLOATING
C4023 a_7826_29789# vssd1 0.626f $ **FLOATING
C4024 a_7994_29535# vssd1 0.581f $ **FLOATING
C4025 a_7553_29423# vssd1 1.43f $ **FLOATING
C4026 _0210_ vssd1 1.2f $ **FLOATING
C4027 a_7387_29423# vssd1 1.81f $ **FLOATING
C4028 a_6269_29423# vssd1 0.23f $ **FLOATING
C4029 a_6779_29789# vssd1 0.609f $ **FLOATING
C4030 a_6947_29691# vssd1 0.817f $ **FLOATING
C4031 a_6354_29789# vssd1 0.626f $ **FLOATING
C4032 a_6522_29535# vssd1 0.581f $ **FLOATING
C4033 a_6081_29423# vssd1 1.43f $ **FLOATING
C4034 _0209_ vssd1 1.2f $ **FLOATING
C4035 a_5915_29423# vssd1 1.81f $ **FLOATING
C4036 ctr\[9\] vssd1 5.74f $ **FLOATING
C4037 a_4797_29423# vssd1 0.23f $ **FLOATING
C4038 a_5307_29789# vssd1 0.609f $ **FLOATING
C4039 a_5475_29691# vssd1 0.817f $ **FLOATING
C4040 a_4882_29789# vssd1 0.626f $ **FLOATING
C4041 a_5050_29535# vssd1 0.581f $ **FLOATING
C4042 a_4609_29423# vssd1 1.43f $ **FLOATING
C4043 _0208_ vssd1 1.11f $ **FLOATING
C4044 a_4443_29423# vssd1 1.81f $ **FLOATING
C4045 clknet_1_1__leaf_io_in[0] vssd1 17.9f $ **FLOATING
C4046 a_2327_29423# vssd1 0.525f $ **FLOATING
C4047 a_1867_29423# vssd1 0.525f $ **FLOATING
C4048 a_1407_29423# vssd1 0.525f $ **FLOATING
C4049 _0044_ vssd1 1.33f $ **FLOATING
C4050 a_12672_30199# vssd1 0.525f $ **FLOATING
C4051 a_12212_30199# vssd1 0.525f $ **FLOATING
C4052 a_11619_29967# vssd1 0.525f $ **FLOATING
C4053 a_10975_29967# vssd1 0.525f $ **FLOATING
C4054 a_10515_29967# vssd1 0.525f $ **FLOATING
C4055 a_10055_29967# vssd1 0.525f $ **FLOATING
C4056 a_9595_29967# vssd1 0.525f $ **FLOATING
C4057 a_9135_29967# vssd1 0.525f $ **FLOATING
C4058 temp1.dac.vdac_single.einvp_batch\[0\].pupd_66.LO vssd1 0.479f $ **FLOATING
C4059 _0404_ vssd1 1.36f $ **FLOATING
C4060 _0218_ vssd1 0.961f $ **FLOATING
C4061 a_15715_30186# vssd1 0.524f $ **FLOATING
C4062 _0814_ vssd1 4.34f $ **FLOATING
C4063 ctr\[10\] vssd1 7.3f $ **FLOATING
C4064 a_6729_30199# vssd1 0.502f $ **FLOATING
C4065 a_3247_29967# vssd1 0.525f $ **FLOATING
C4066 a_1407_29967# vssd1 0.227f $ **FLOATING
C4067 a_4003_30006# vssd1 0.59f $ **FLOATING
C4068 a_3749_30006# vssd1 0.607f $ **FLOATING
C4069 net66 vssd1 1.2f $ **FLOATING
C4070 temp1.dac.vdac_single.en_pupd vssd1 1.12f $ **FLOATING
C4071 a_2805_30265# vssd1 0.607f $ **FLOATING
C4072 _0800_ vssd1 7.3f $ **FLOATING
C4073 _0801_ vssd1 8.78f $ **FLOATING
C4074 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 7.94f $ **FLOATING
C4075 a_2376_30199# vssd1 0.59f $ **FLOATING
C4076 _0833_ vssd1 0.77f $ **FLOATING
C4077 a_2060_30199# vssd1 0.535f $ **FLOATING
C4078 a_1741_30199# vssd1 0.5f $ **FLOATING
C4079 a_1554_29941# vssd1 0.578f $ **FLOATING
C4080 a_1458_30199# vssd1 0.498f $ **FLOATING
C4081 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vssd1 1.44f $ **FLOATING
C4082 a_11619_30511# vssd1 0.525f $ **FLOATING
C4083 a_11292_30663# vssd1 0.525f $ **FLOATING
C4084 a_10832_30663# vssd1 0.525f $ **FLOATING
C4085 net13 vssd1 5.67f $ **FLOATING
C4086 a_10239_30511# vssd1 0.525f $ **FLOATING
C4087 a_9687_30511# vssd1 0.525f $ **FLOATING
C4088 a_9360_30663# vssd1 0.525f $ **FLOATING
C4089 a_8543_30485# vssd1 0.698f $ **FLOATING
C4090 a_6835_30511# vssd1 0.524f $ **FLOATING
C4091 _0835_ vssd1 2.36f $ **FLOATING
C4092 a_4811_30511# vssd1 0.648f $ **FLOATING
C4093 _0834_ vssd1 1.01f $ **FLOATING
C4094 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 3.64f $ **FLOATING
C4095 a_4484_30663# vssd1 0.525f $ **FLOATING
C4096 _0773_ vssd1 7f $ **FLOATING
C4097 a_2419_30511# vssd1 0.525f $ **FLOATING
C4098 _0831_ vssd1 2.23f $ **FLOATING
C4099 a_2009_30676# vssd1 0.524f $ **FLOATING
C4100 net8 vssd1 8.45f $ **FLOATING
C4101 net14 vssd1 5.54f $ **FLOATING
C4102 a_9779_31055# vssd1 0.525f $ **FLOATING
C4103 a_9319_31055# vssd1 0.525f $ **FLOATING
C4104 a_8123_31055# vssd1 0.525f $ **FLOATING
C4105 a_7663_31055# vssd1 0.525f $ **FLOATING
C4106 a_7203_31055# vssd1 0.525f $ **FLOATING
C4107 a_6375_31055# vssd1 0.525f $ **FLOATING
C4108 a_4351_31055# vssd1 0.388f $ **FLOATING
C4109 a_5823_31055# vssd1 0.525f $ **FLOATING
C4110 a_4811_31055# vssd1 0.525f $ **FLOATING
C4111 a_3891_31055# vssd1 0.525f $ **FLOATING
C4112 a_2879_31055# vssd1 0.525f $ **FLOATING
C4113 a_2552_31287# vssd1 0.525f $ **FLOATING
C4114 a_2092_31287# vssd1 0.525f $ **FLOATING
C4115 net9 vssd1 7.38f $ **FLOATING
C4116 a_10844_31029# vssd1 0.648f $ **FLOATING
C4117 a_10239_31055# vssd1 0.698f $ **FLOATING
C4118 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd vssd1 1.36f $ **FLOATING
C4119 _0817_ vssd1 12.2f $ **FLOATING
C4120 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 4.28f $ **FLOATING
C4121 a_10924_31751# vssd1 0.525f $ **FLOATING
C4122 a_10239_31599# vssd1 0.525f $ **FLOATING
C4123 a_9779_31599# vssd1 0.525f $ **FLOATING
C4124 a_9319_31599# vssd1 0.525f $ **FLOATING
C4125 a_8951_31599# vssd1 0.648f $ **FLOATING
C4126 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref vssd1 2.33f $ **FLOATING
C4127 a_8532_31751# vssd1 0.525f $ **FLOATING
C4128 a_7847_31599# vssd1 0.525f $ **FLOATING
C4129 a_7387_31599# vssd1 0.525f $ **FLOATING
C4130 a_7060_31751# vssd1 0.525f $ **FLOATING
C4131 a_6467_31599# vssd1 0.525f $ **FLOATING
C4132 a_6007_31599# vssd1 0.525f $ **FLOATING
C4133 a_5547_31599# vssd1 0.525f $ **FLOATING
C4134 a_5087_31599# vssd1 0.525f $ **FLOATING
C4135 a_4351_31599# vssd1 0.525f $ **FLOATING
C4136 a_3891_31599# vssd1 0.525f $ **FLOATING
C4137 net65 vssd1 1.33f $ **FLOATING
C4138 temp1.dac.vdac_single.einvp_batch\[0\].vref_65.HI vssd1 0.415f $ **FLOATING
C4139 a_9452_32375# vssd1 0.525f $ **FLOATING
C4140 a_8348_32375# vssd1 0.525f $ **FLOATING
C4141 a_7888_32375# vssd1 0.525f $ **FLOATING
C4142 a_6835_32143# vssd1 0.525f $ **FLOATING
C4143 a_6508_32375# vssd1 0.525f $ **FLOATING
C4144 a_4811_32143# vssd1 0.525f $ **FLOATING
C4145 a_4484_32375# vssd1 0.525f $ **FLOATING
C4146 a_3891_32143# vssd1 0.525f $ **FLOATING
C4147 net11 vssd1 5.66f $ **FLOATING
C4148 net10 vssd1 8.75f $ **FLOATING
C4149 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 7.27f $ **FLOATING
C4150 temp1.dac_vout_notouch_ vssd1 52.3f $ **FLOATING
C4151 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vssd1 4.74f $ **FLOATING
C4152 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 6.84f $ **FLOATING
.ends

* PEX produced on Wed Apr 19 01:52:19 PM CEST 2023 using /foss/tools/iic-osic/iic-pex.sh with m=1 and s=1
* NGSPICE file created from hpretl_tt03_temperature_sensor.ext - technology: sky130A

.subckt hpretl_tt03_temperature_sensor io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_in[0] vccd1 vssd1
X0 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 vccd1 a_7389_25335# _0825_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 vssd1 a_7226_16885# _0518_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 _0594_.C a_15759_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 vssd1 a_28015_5755# a_27973_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5 a_10356_10089# _0475_.X a_9895_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X6 a_16573_26159# _1052_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 _0544_.C a_13551_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X10 vccd1 _0679_.A1 a_8478_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X11 _1019_.Q a_21759_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_10309_9673# a_9319_9301# a_10183_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14 vccd1 _0523_.B1 a_16853_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X15 vccd1 a_2114_1653# _0860_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X17 vccd1 _0893_.CLK a_24775_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X18 vssd1 _0660_.X a_20635_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_19099_4943# a_18317_4949# a_19015_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 a_3394_26677# a_3226_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X22 _1057_.Q a_15503_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_24209_20175# _0965_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 _0845_.Y _0845_.C1 a_3993_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X28 a_14913_14013# _0511_.D a_14813_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X29 vssd1 _0927_.D a_22940_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X30 a_9942_11471# a_9503_11477# a_9857_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X32 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15916_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X33 vccd1 a_23891_17999# a_24059_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X34 vccd1 _0582_.A a_20083_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_11782_18909# a_11343_18543# a_11697_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X36 a_14372_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X37 vssd1 _0844_.B a_3154_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X38 vssd1 a_10811_2741# a_10769_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X39 a_9865_11249# _0466_.A a_9284_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X40 vccd1 a_4040_10901# _0745_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X42 a_9765_4399# _0959_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X43 vssd1 a_24335_6005# a_24293_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X44 vccd1 _0521_.A a_13183_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X45 a_12441_17705# _0797_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X46 vssd1 a_8545_14709# _0546_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X47 _0798_.A2 _0722_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X48 vssd1 fanout23.X a_25235_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X50 _0607_.B a_21575_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X51 a_4847_2589# a_4149_2223# a_4590_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X52 vccd1 clkbuf_1_0__f_io_in[0].X a_1591_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X54 _0845_.C1 a_4811_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_7939_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 vssd1 a_5383_2741# a_5341_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X58 vccd1 _0566_.A1 a_10613_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X60 a_26099_25615# a_25401_25621# a_25842_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X62 vccd1 a_9926_9269# a_9853_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X64 a_25306_6941# a_24867_6575# a_25221_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X65 vccd1 a_2658_25183# a_2585_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X66 a_10459_13647# a_9761_13653# a_10202_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X68 a_19697_2773# a_19531_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 a_2823_27613# a_1959_27247# a_2566_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X70 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X71 a_10034_13647# a_9595_13653# a_9949_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X73 a_21499_21085# a_20635_20719# a_21242_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X74 a_12245_6031# a_11711_6037# a_12150_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X75 vccd1 _0809_.B2 a_4863_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X76 a_9230_16143# _0842_.A0 a_9003_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X77 vccd1 a_17725_15073# _0487_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X78 a_4221_8725# _0711_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X79 a_22905_17455# _0994_.Q a_22833_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X80 vssd1 a_3559_4943# a_3727_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X81 a_27337_3311# _1069_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X82 a_25225_14441# _0966_.Q a_25143_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X83 vccd1 _0527_.X a_16127_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X85 vccd1 _0807_.B a_11885_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X86 a_15427_3855# a_14729_3861# a_15170_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X88 a_10126_22351# a_9687_22357# a_10041_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X89 a_22637_16367# _1019_.Q a_22291_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X92 a_2493_27613# a_1959_27247# a_2398_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X93 a_20709_5853# a_20175_5487# a_20614_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X94 vccd1 a_21426_19743# a_21353_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X95 vccd1 _0805_.A a_4386_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X96 a_8473_7125# a_8307_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X97 a_21169_21085# a_20635_20719# a_21074_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X98 vccd1 a_21115_21237# a_21031_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X99 vssd1 a_21039_5853# a_21207_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X100 a_22181_16917# a_22015_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 vssd1 _0722_.A _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X102 a_14637_18005# a_14471_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X103 _0650_.X a_25511_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X104 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X107 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X109 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X110 vssd1 _0829_.A1 _0864_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X112 a_14139_4943# a_13275_4949# a_13882_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X113 vssd1 a_16897_12897# _0533_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X114 a_13265_7485# _0521_.A a_13183_7232# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X115 _0807_.B a_9043_12567# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X118 vssd1 _0679_.A2 a_8033_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X119 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X120 a_5483_4765# a_4701_4399# a_5399_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 a_6553_17705# _0717_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X124 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X125 vccd1 a_25658_8863# a_25585_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X127 vccd1 a_23047_22325# a_22963_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X129 vccd1 _0471_.X a_12763_12879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X130 a_26413_18543# a_26247_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X131 vssd1 _0844_.B a_4902_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X132 vccd1 a_16515_20987# a_16431_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X133 a_19793_15279# _0962_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X134 vccd1 _0619_.B1 a_23201_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X136 a_22269_2223# a_21279_2223# a_22143_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X137 a_22963_1679# a_22181_1685# a_22879_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 a_3057_18319# _0872_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X139 vccd1 clkbuf_1_1__f__0390_.A a_2686_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X140 a_17773_15529# _0522_.X a_17691_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X142 _0814_.B1 _0798_.A2 a_5909_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 _1050_.Q a_19183_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X146 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 temp1.capload\[10\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X147 a_10084_9839# _0545_.B1 a_9993_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X148 a_19107_21263# a_18409_21269# a_18850_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X149 a_6449_2589# a_5915_2223# a_6354_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X150 _1050_.Q a_19183_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 a_1674_32143# clkbuf_1_1__f_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X153 a_20755_14735# a_19973_14741# a_20671_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 a_20985_19631# a_20819_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X156 _0472_.X a_8859_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X158 a_22169_6397# _0575_.B a_22097_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 vssd1 a_17435_22075# a_17393_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X162 vccd1 _0922_.CLK a_2787_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X164 a_17420_18319# _0522_.B1 a_16929_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X165 a_8763_14735# _0546_.B1 a_8545_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X166 vssd1 a_15963_1653# a_15921_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X168 a_24941_23445# a_24775_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X169 vccd1 _0740_.X a_4769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X170 _1042_.Q a_18447_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X171 vssd1 _0662_.A3 a_16097_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X172 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X173 vccd1 a_15963_27765# a_15879_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X174 vssd1 _0872_.A1 a_4705_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X175 vccd1 a_20195_6005# a_20111_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X176 a_2455_9117# a_1757_8751# a_2198_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X177 _0920_.Q a_16515_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X178 a_14269_20181# a_14103_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X179 _0588_.A1 a_15319_12283# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X180 a_11908_20719# a_11509_20719# a_11782_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X181 vccd1 a_15078_17973# a_15005_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X182 a_4769_23145# _0788_.C a_4403_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X183 a_12893_21807# a_12716_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X185 a_9999_1501# a_9301_1135# a_9742_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X187 a_23837_9295# a_23303_9301# a_23742_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X188 vccd1 a_7902_6005# a_7829_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X189 vssd1 a_12743_8181# a_12701_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X190 a_9853_9295# a_9319_9301# a_9758_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X191 vccd1 fanout23.X a_26983_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X192 vssd1 _0734_.A2 _0696_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X193 a_27847_10205# a_26983_9839# a_27590_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X196 a_20387_15645# a_19605_15279# a_20303_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X200 a_12428_1135# a_11895_1385# _0854_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X202 a_12207_18909# a_11343_18543# a_11950_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X203 a_25401_7125# a_25235_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X206 a_25497_12015# _0893_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X207 a_15611_3677# a_14913_3311# a_15354_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X208 vccd1 a_2626_9269# _0835_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X210 _1012_.Q a_28015_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X211 vccd1 _0670_.A2 a_15005_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X212 a_8803_4943# a_8105_4949# a_8546_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X213 a_22653_9295# _0620_.X a_22547_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X214 a_6682_27907# _0825_.A0 a_6600_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X215 a_9333_16143# _0838_.A0 a_9230_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X216 a_15929_4399# _0497_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X217 vssd1 _0888_.CLK a_4627_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X218 _0843_.Y _0843_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X219 a_2953_26709# a_2787_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X220 a_16826_26271# a_16658_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X222 vssd1 _0717_.A2 a_10585_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X223 a_7829_6031# a_7295_6037# a_7734_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X224 vssd1 a_12316_24135# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X225 vccd1 a_16090_20831# a_16017_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X226 a_25432_6575# a_25033_6575# a_25306_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X227 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X229 a_2585_25621# a_2419_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 vssd1 a_22990_14303# a_22948_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X231 _0860_.A a_2114_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X232 a_5888_31055# a_5639_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X233 vccd1 a_22879_20175# a_23047_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X234 _0987_.D a_9983_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X235 a_2673_4233# a_1683_3861# a_2547_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X238 vssd1 _1053_.CLK a_14563_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X239 vccd1 a_2566_27359# a_2493_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X240 a_25401_25621# a_25235_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X241 vccd1 a_10627_13621# a_10543_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X242 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X243 vccd1 _0438_.A a_9043_12567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X244 a_12736_21641# a_12337_21269# a_12610_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X245 a_16090_20831# a_15922_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X246 vssd1 a_22879_20175# a_23047_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X248 vccd1 _0824_.Y a_13183_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X249 a_2686_10383# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X250 a_21994_22173# a_21555_21807# a_21909_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X253 a_12981_9301# a_12815_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X254 vssd1 _0874_.X a_2684_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X256 a_23650_21263# a_23211_21269# a_23565_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X258 vccd1 _1077_.Q a_9963_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X259 vccd1 a_18355_6005# a_18271_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X260 a_25585_9117# a_25051_8751# a_25490_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X261 _0776_.A2 a_7623_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X262 a_13771_22351# a_13073_22357# a_13514_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X263 _0684_.A1 _0644_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 a_19099_20175# a_18317_20181# a_19015_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X266 vccd1 a_19770_3829# a_19697_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X267 vssd1 _0745_.A1 a_6563_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X269 vssd1 a_20303_15645# a_20471_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X270 vccd1 _0873_.Y a_2599_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X271 a_22461_2767# _0497_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X272 vccd1 _0685_.B a_6498_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X274 _0673_.A1 a_12927_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X276 a_4248_29673# _0845_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X277 a_21718_2589# a_21445_2223# a_21633_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X278 vccd1 a_15170_23413# a_15097_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X279 vccd1 a_7775_3829# a_7691_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X280 _0506_.X a_22659_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X281 a_15105_11471# _0588_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X282 vccd1 temp1.capload\[14\].cap_44.LO temp1.capload\[14\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X283 a_27422_10205# a_27149_9839# a_27337_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X284 vccd1 _0827_.A a_7479_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X286 _0471_.X a_9503_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X288 a_4337_1135# _0849_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X289 a_2381_16885# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X290 vssd1 a_23139_2741# a_23097_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X291 a_8746_7119# a_8307_7125# a_8661_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X292 a_22373_12559# _0563_.B1 a_22457_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X293 a_10948_21813# _0441_.B a_10876_21813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X294 a_2136_9673# a_1757_9301# a_2039_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X295 a_5445_24527# _0809_.B2 _0788_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X296 a_2566_1247# a_2398_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X297 a_21357_13103# _0890_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X299 a_23634_26677# a_23466_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X301 a_13360_25935# _0824_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X302 a_6559_19087# _0440_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X303 vssd1 _0675_.C a_15391_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
R1 vccd1 temp1.capload\[6\].cap_51.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X304 a_25217_7663# a_25051_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X305 vssd1 fanout10.A a_10791_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X307 a_21775_18909# a_20911_18543# a_21518_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X309 vccd1 _0917_.CLK a_14287_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X310 vccd1 a_17895_10357# a_17811_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X311 vssd1 fanout9.A a_12999_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X312 a_26225_5321# a_25235_4949# a_26099_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X313 a_10126_6031# a_9853_6037# a_10041_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X314 a_14089_19087# _0936_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X315 _0919_.D a_12375_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X316 _0545_.B2 a_14011_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X317 vccd1 temp1.inv1_1.Y a_1766_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X319 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X320 a_5361_30287# _0809_.B2 a_5141_30199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X322 a_27337_7663# _1064_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X323 a_23466_26703# a_23193_26709# a_23381_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X325 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 a_8305_19087# _0761_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X329 a_13616_28879# a_13367_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X330 a_12725_19087# _0864_.Y _0865_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 a_25401_1135# a_25235_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X333 vccd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_2686_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X334 a_21445_18909# a_20911_18543# a_21350_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X335 a_9301_1135# a_9135_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X337 _0616_.B1 a_16771_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X338 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X339 vssd1 _0893_.CLK a_26983_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X341 a_11831_3677# a_11049_3311# a_11747_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X342 a_15446_2335# a_15278_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X343 temp1.capload\[5\].cap.Y temp1.capload\[5\].cap_50.LO a_10509_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X345 a_16009_9001# _0587_.X a_15937_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X346 a_7479_29673# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R2 vssd1 temp1.capload\[9\].cap_54.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X347 a_7097_3855# _0622_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 vssd1 a_25715_13371# a_25673_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X350 a_15446_2335# a_15278_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X351 vssd1 a_25807_23413# a_25765_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X352 vccd1 a_27590_21919# a_27517_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X354 a_27149_9839# a_26983_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X355 vccd1 _0444_.A _0444_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X356 a_8937_3855# _0902_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X357 vssd1 a_25623_5755# a_25581_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X359 a_11437_16617# _0827_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X360 vssd1 _0679_.A2 a_8393_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X361 vssd1 _0471_.X a_10183_12061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X363 vssd1 a_15135_20149# a_15093_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X364 a_25971_13647# _0648_.B1 a_26053_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X365 a_25769_16911# a_25235_16917# a_25674_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X366 a_17470_3829# a_17302_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X367 a_22454_1679# a_22015_1685# a_22369_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X368 vccd1 _1015_.CLK a_23671_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X370 _0814_.A1 clkbuf_1_1__f_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X371 a_9436_16143# _0508_.Y a_9333_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X373 a_27590_21919# a_27422_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X374 a_11950_18655# a_11782_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X375 vccd1 _0602_.A a_18887_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X377 vssd1 a_9615_3829# a_9573_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X380 a_27422_8029# a_26983_7663# a_27337_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X381 a_20161_14735# _1024_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 _0969_.D a_23415_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X384 _0666_.D a_25143_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X386 a_5813_10383# _0745_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X387 vssd1 _0922_.CLK a_11711_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X389 a_15365_5059# _0556_.B a_15293_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X391 vccd1 a_4403_25589# _0840_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X392 a_7829_15529# _0760_.B2 a_7745_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X393 a_2949_2223# a_1959_2223# a_2823_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X394 vccd1 a_24535_11471# a_24703_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X395 a_21169_13103# a_21003_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X396 vccd1 _0535_.X a_11333_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X397 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X398 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X399 a_12801_15823# _0920_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X401 vccd1 _0456_.B _0722_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X402 vssd1 a_25474_6687# a_25432_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X403 vssd1 a_24535_11471# a_24703_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X404 vssd1 a_4864_11445# _0745_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X405 a_4337_26159# _0843_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X406 fanout23.X a_27202_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X407 a_14093_7235# _0544_.D a_14011_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X408 a_27422_25437# a_26983_25071# a_27337_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X410 a_1674_26159# clkbuf_1_1__f_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X411 a_25125_22173# a_24591_21807# a_25030_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X412 vccd1 _0572_.X a_19689_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X413 a_5177_27023# _0835_.A1 _0835_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X415 a_20345_20175# _1061_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X416 vssd1 _0908_.CLK a_6743_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X417 a_22273_2773# a_22107_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X418 a_25842_21237# a_25674_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X419 a_25674_7119# a_25235_7125# a_25589_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X420 vccd1 _0696_.A1 _0698_.A2_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X421 a_20385_12043# _0842_.A0 a_20299_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X422 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15023_28887# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X423 vccd1 _1075_.Q a_14729_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X424 a_17995_17821# a_17213_17455# a_17911_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X426 a_19969_11791# _1057_.Q a_19531_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X427 vssd1 _0474_.X _0630_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X428 _0494_.X a_14637_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X429 _1078_.D _0840_.X a_1591_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 vccd1 _1078_.Q a_14287_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X432 a_12521_4399# a_12355_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X433 a_18455_11293# a_17673_10927# a_18371_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X434 vccd1 _0795_.A2_N a_6646_18865# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X437 vssd1 _1077_.Q a_9963_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X438 a_26099_15823# a_25401_15829# a_25842_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X439 a_4429_16672# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X441 vssd1 a_17251_26427# a_17209_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X442 a_27590_17567# a_27422_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X443 vccd1 _1028_.CLK a_10423_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X444 _1006_.D a_27739_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X445 a_6653_10933# _0746_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 a_25674_21263# a_25401_21269# a_25589_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X447 a_17231_19200# _1061_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X448 a_21502_15529# _0998_.D a_21345_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X449 a_17819_1679# a_16955_1685# a_17562_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X450 a_7599_5853# a_6817_5487# a_7515_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X452 vssd1 a_27847_17821# a_28015_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X454 a_17470_3829# a_17302_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X456 a_5913_25335# _0445_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X457 vccd1 _0888_.CLK a_7295_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X458 vccd1 a_14307_4917# a_14223_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X460 a_18969_17277# _0602_.A a_18887_17024# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X462 a_15759_1385# _0645_.B1 a_15841_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X464 vssd1 a_7902_6005# a_7860_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X465 a_25030_2589# a_24591_2223# a_24945_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X467 _1045_.D a_19827_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X468 a_8872_7497# a_8473_7125# a_8746_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X469 temp1.capload\[4\].cap.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X470 vssd1 a_18758_4917# a_18716_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X471 vssd1 _0523_.B1 a_22637_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X472 a_5724_19881# _0722_.C a_5642_19637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X474 a_21518_18655# a_21350_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X475 vssd1 a_17562_1653# a_17520_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X476 _0760_.B2 _0717_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X477 a_21591_27613# a_20893_27247# a_21334_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X479 vssd1 _0643_.B1 a_24212_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X480 a_13906_12925# _0840_.A0 a_13817_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X481 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13616_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X483 _0797_.A1 a_5549_17719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X484 a_12355_8751# _0472_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X485 _0845_.C1 a_4811_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X486 a_15377_16367# _0990_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X487 vssd1 a_16897_16395# _0522_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X488 vccd1 _0579_.C a_17231_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X489 vccd1 a_21518_18655# a_21445_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X490 a_23331_3677# a_22549_3311# a_23247_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X491 vccd1 _0479_.Y a_13551_8215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X492 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X493 a_26007_3677# a_25309_3311# a_25750_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X494 vccd1 a_20839_7931# a_20755_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X495 _0708_.A2 a_4447_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X496 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A _0825_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X497 a_26962_13469# a_26523_13103# a_26877_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X498 a_8749_3861# a_8583_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X499 a_13422_9269# a_13254_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X500 a_24535_11471# a_23671_11477# a_24278_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X501 vssd1 _0512_.X a_19693_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X502 vssd1 a_25842_21237# a_25800_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X503 a_5115_1679# a_4333_1685# a_5031_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X504 a_27517_15645# a_26983_15279# a_27422_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X505 a_25489_14191# _0996_.Q a_25143_14441# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X506 a_25539_2589# a_24757_2223# a_25455_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X507 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_13984_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X508 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X509 a_7801_11079# _0438_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X511 vssd1 a_15078_17973# a_15036_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X512 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X513 a_16014_14557# a_15741_14191# a_15929_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X514 a_16863_7119# _0487_.X a_17041_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X515 vssd1 a_26267_19899# a_26225_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X516 vccd1 _0535_.X a_12797_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X519 a_27931_14557# a_27149_14191# a_27847_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X520 _0545_.B1 a_19439_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X521 a_12276_14025# a_11877_13653# a_12150_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X522 a_24757_21807# a_24591_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X523 vssd1 _0877_.A2 a_4621_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X524 vssd1 _1028_.CLK a_9687_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X525 a_21499_21085# a_20801_20719# a_21242_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X527 a_10567_19061# _0771_.C1 a_10998_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X528 _0893_.CLK a_23487_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X529 a_21074_21085# a_20635_20719# a_20989_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X530 _0962_.D a_15319_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X531 a_13073_22357# a_12907_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X532 vssd1 _0964_.CLK a_26983_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X533 vssd1 _0621_.X _0624_.D_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X534 a_2999_28701# a_2217_28335# a_2915_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X536 vssd1 _0438_.A a_8122_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X537 a_4769_22895# _0742_.A2 a_4959_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X538 a_24297_13653# a_24131_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 a_25674_21263# a_25235_21269# a_25589_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X540 a_22580_2057# a_22181_1685# a_22454_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X541 a_6559_10383# _0655_.X _0656_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X542 vccd1 a_19199_25615# a_19367_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X543 vccd1 _0574_.C a_17725_15073# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X544 a_24209_1679# _0976_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X545 vccd1 _0850_.A a_7389_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X546 a_9942_11471# a_9669_11477# a_9857_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X547 a_5537_15529# _0758_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X548 vccd1 _1075_.Q a_15115_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X549 vccd1 _1062_.CLK a_19991_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X550 vssd1 a_6062_3423# a_6020_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X551 _1055_.Q a_13939_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X552 vccd1 a_19045_15797# _0658_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X553 a_26597_4399# a_26431_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X554 a_27548_7663# a_27149_7663# a_27422_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X556 vssd1 a_19199_25615# a_19367_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X557 vssd1 _0964_.CLK a_25235_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X558 vccd1 a_15812_6005# _0675_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X559 vssd1 _0479_.Y a_11435_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X560 vccd1 a_25198_21919# a_25125_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X561 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X562 vssd1 a_23247_3677# a_23415_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X563 vssd1 a_23431_7119# a_23599_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X564 _1055_.Q a_13939_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X565 vccd1 _0656_.Y a_6815_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X570 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X571 vssd1 a_8307_17455# _1053_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X572 vssd1 _0863_.A2 a_15777_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X573 a_21997_26159# a_21831_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X574 vccd1 _0735_.A2 a_9301_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.1525 ps=1.305 w=1 l=0.15
X575 vccd1 _0840_.A0 a_12355_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X576 _0789_.B1 a_5913_25335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X577 vssd1 a_21426_19743# a_21384_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X579 a_11287_11293# a_10423_10927# a_11030_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X582 a_25800_7497# a_25401_7125# a_25674_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X583 a_23469_9301# a_23303_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X584 vccd1 a_25915_17821# a_26083_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X585 a_5069_4765# a_4535_4399# a_4974_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X587 vssd1 a_28015_22075# a_27973_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X588 a_24945_16367# _0938_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X589 a_17378_19743# a_17210_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X590 vssd1 _0579_.C a_17995_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X591 a_9485_9301# a_9319_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X592 _0745_.A2 a_4040_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X594 vccd1 a_18095_23261# a_18263_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X595 a_5612_8207# _0694_.A2 a_5510_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X596 a_24110_11471# a_23837_11477# a_24025_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X597 _0861_.A1 _0860_.A a_16581_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X598 a_3141_19148# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X600 a_4959_22895# _0809_.B2 a_4403_22869# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X601 vssd1 _0797_.A1 a_14644_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X602 vssd1 _0574_.C a_22905_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X603 a_15151_10205# a_14287_9839# a_14894_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X605 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X606 a_19969_16367# _0963_.D a_19531_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X607 a_15565_11177# _0614_.D a_15483_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X608 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12065_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X609 a_22549_1679# a_22015_1685# a_22454_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X610 a_19770_26677# a_19602_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X611 vccd1 a_26267_15797# a_26183_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X612 a_5445_9295# _0710_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X613 vccd1 _0825_.A0 _0815_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X616 vssd1 a_11435_22895# _0847_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X617 a_20414_14709# a_20246_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X618 _0694_.A2 _0681_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.12675 ps=1.04 w=0.65 l=0.15
X619 vssd1 a_22311_2491# a_22269_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X621 a_18095_23261# a_17397_22895# a_17838_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X623 a_4590_26271# a_4422_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X624 vccd1 a_21886_2335# a_21813_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X625 a_16025_14013# _0583_.A a_15943_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X627 a_24845_2057# a_23855_1685# a_24719_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X628 vssd1 a_19015_4943# a_19183_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X629 vssd1 a_3394_26677# a_3352_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X630 a_20690_21237# a_20522_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X631 a_23661_14735# _0648_.A2 a_23745_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 a_25156_2223# a_24757_2223# a_25030_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X633 _0529_.Y _0836_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X635 vccd1 _0512_.A a_18611_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X636 a_20897_4399# _0649_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X637 a_23013_4399# _0548_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X638 vssd1 a_3026_25589# a_2984_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X639 a_7829_21269# a_7663_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X640 a_14341_17429# _0798_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X641 a_25129_8207# _0621_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X642 a_11238_17705# _0833_.A a_11041_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X643 a_5629_17027# _0807_.B a_5547_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X645 a_24397_10749# _0602_.A a_24315_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X646 a_23741_8585# a_22751_8213# a_23615_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X647 a_11938_25071# _0847_.A3 a_11848_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X648 a_20598_20149# a_20430_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X650 vccd1 _0713_.A1 _0758_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X652 vccd1 _0908_.CLK a_4167_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X655 a_19199_25615# a_18335_25621# a_18942_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X656 vccd1 a_10294_6005# a_10221_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X657 _0563_.C1 a_24591_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X659 vssd1 a_26007_10205# a_26175_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X660 a_3651_26703# a_2953_26709# a_3394_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X661 vccd1 a_10055_23983# _0847_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X662 _0936_.Q a_8695_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X664 _0746_.A2 _0679_.A2 a_8116_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X665 a_22622_22325# a_22454_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X666 vccd1 _0583_.A a_17139_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X667 a_3512_16911# _0722_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X668 vssd1 a_13479_15797# a_13437_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X669 vssd1 _0959_.CLK a_9779_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X670 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X671 _0443_.A a_10789_22071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X672 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X673 _0582_.A a_13551_8215# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X674 vssd1 a_10294_22325# a_10252_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X675 _0624_.D_N _0623_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X676 vccd1 a_27847_5853# a_28015_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X677 a_15277_12015# a_14287_12015# a_15151_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X678 a_15235_12381# a_14453_12015# a_15151_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X680 vssd1 a_18942_25589# a_18900_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X681 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10488_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X682 a_5617_5321# a_4627_4949# a_5491_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X683 _1006_.D a_27739_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X684 vccd1 _0523_.B1 a_20257_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X685 vssd1 a_8971_1653# a_8929_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X686 a_22454_22351# a_22181_22357# a_22369_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X687 vssd1 _0648_.A2 a_23649_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X688 a_9184_25223# _0825_.A1 a_9326_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X689 temp1.capload\[15\].cap.Y temp1.capload\[15\].cap_45.LO a_15017_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 vssd1 _0807_.C a_8241_16161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 a_26099_7119# a_25401_7125# a_25842_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X692 vccd1 a_17928_8181# _0587_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X693 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_14287_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X694 _0825_.A1 a_7389_25335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X695 vssd1 a_10814_15797# _0529_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X696 _0518_.Y a_7226_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X697 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X698 a_21334_27359# a_21166_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X699 vssd1 _0920_.D a_17420_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X700 a_27571_6941# a_26873_6575# a_27314_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X701 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X703 a_10735_2589# a_9871_2223# a_10478_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X704 vssd1 a_2382_4511# a_2340_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X706 a_24757_21807# a_24591_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X707 a_8101_15279# _0439_.A a_7663_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X709 vccd1 a_27130_13215# a_27057_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X710 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_14372_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X711 a_17260_12265# _0565_.B1 a_17158_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X713 a_9687_23439# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X714 _0935_.CLK a_10791_16919# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X715 a_17086_17999# _0577_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X718 vccd1 _0583_.A a_19439_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X721 vssd1 _0445_.A a_7544_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
X722 a_19973_14741# a_19807_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X723 vssd1 a_20690_21237# a_20648_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X724 vssd1 a_27590_7775# a_27548_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X725 a_20847_9633# _0582_.A a_20761_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X728 a_10386_2741# a_10218_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X729 _0664_.X a_25971_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X731 a_10769_2057# a_9779_1685# a_10643_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X732 vccd1 a_10167_5755# a_10083_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X733 a_13679_9295# a_12981_9301# a_13422_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X734 a_23201_10089# _1069_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X735 a_26210_26271# a_26042_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X737 a_23193_18005# a_23027_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X738 a_11705_6575# _0921_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X739 a_17727_3855# a_16863_3861# a_17470_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X740 a_23649_4399# a_22659_4399# a_23523_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X741 vccd1 _0764_.A1 a_6682_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X742 vccd1 _0783_.A1 a_5819_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X744 a_4958_2741# a_4790_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X745 _0837_.A1 a_2991_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X746 vccd1 _1028_.CLK a_12539_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X747 _0908_.CLK a_1959_4951# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X749 a_20947_21263# a_20249_21269# a_20690_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X750 a_10133_1679# _0639_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X751 a_26827_23261# a_26045_22895# a_26743_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X752 vccd1 a_3523_13655# _0768_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X753 vssd1 a_22622_22325# a_22580_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X754 _0768_.A2 _0684_.A2 a_7745_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X755 a_1757_9301# a_1591_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X756 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X757 vssd1 _0505_.X a_22659_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X758 a_25382_12533# a_25214_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X759 a_6423_8903# _0681_.X a_6892_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X760 vssd1 _1015_.CLK a_25051_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X761 a_21813_2589# a_21279_2223# a_21718_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X763 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X764 vccd1 a_11895_1385# _0854_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X765 a_8887_4943# a_8105_4949# a_8803_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X767 a_20165_16189# _0582_.A a_20083_15936# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X770 a_2566_27359# a_2398_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X772 _0666_.B a_20635_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X773 vssd1 a_16495_5487# fanout24.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X774 vssd1 a_17470_3829# a_17428_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X775 _0634_.B1 a_18519_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X776 vccd1 a_11764_20149# _0858_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X777 vccd1 a_5600_14165# _0736_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X778 vccd1 a_17987_1653# a_17903_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X779 _1067_.D a_27555_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X781 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X782 vssd1 _0456_.B a_3435_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X784 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X785 a_10221_6031# a_9687_6037# a_10126_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X787 a_15538_1653# a_15370_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X789 vssd1 _0679_.A1 a_8033_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X790 a_16771_9001# _0630_.A2 a_16853_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X791 a_21213_12043# _0512_.A a_21127_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X792 a_4989_12879# _0791_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X794 vccd1 a_1585_24135# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X795 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9769_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X796 vssd1 _0964_.CLK a_22015_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X797 vssd1 a_25198_2335# a_25156_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X798 vccd1 _0823_.A a_11746_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X799 vccd1 _0532_.A2 a_14661_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X803 _0717_.B1 _0714_.B1 a_9312_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.069875 ps=0.865 w=0.65 l=0.15
X804 a_25401_1135# a_25235_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 a_4701_4399# a_4535_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X806 vssd1 _0812_.A2 a_9492_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X807 a_9301_1135# a_9135_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X808 a_7663_12879# _0684_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X809 a_9993_9839# _0466_.A a_9895_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X810 a_4422_2589# a_3983_2223# a_4337_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X812 vssd1 _0630_.X a_15671_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X813 _0737_.X a_8256_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X814 vccd1 clkbuf_1_1__f__0390_.A a_2686_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X815 vssd1 _0999_.CLK a_23855_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X816 _1064_.Q a_27003_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X817 vssd1 _1062_.CLK a_26247_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X818 vssd1 _0572_.A2 a_22085_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X819 _0798_.X a_4036_30663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X820 _0722_.B _0456_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X821 a_7649_6031# _0611_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X822 vssd1 a_18355_6005# a_18313_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X823 _0666_.X a_21831_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X824 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X825 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14563_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X826 vssd1 a_5015_26427# a_4973_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X827 vssd1 a_11929_9633# _0491_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X828 a_20993_1385# _1034_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X829 a_27130_13215# a_26962_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X831 a_27149_2223# a_26983_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X832 _0651_.X a_22199_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X833 _0662_.A3 a_14453_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X834 a_18505_4943# _0543_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X835 _0684_.A1 _0651_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X836 vssd1 a_5642_19637# _0761_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X839 a_17309_1679# _0515_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X840 a_5909_26159# _0827_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X841 a_20939_20175# a_20157_20181# a_20855_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X842 a_22817_18517# _0662_.B1 a_22974_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X843 vccd1 a_23047_16885# a_22963_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X844 a_24757_15279# a_24591_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X847 vssd1 fanout23.X a_26983_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X848 vssd1 a_20027_6031# a_20195_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X849 a_26505_11293# a_25971_10927# a_26410_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X850 vccd1 a_4259_6031# _0922_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X852 vccd1 a_5015_2491# _0829_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X853 a_20025_10955# _0602_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X854 vccd1 a_15905_25589# _0861_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X856 a_2584_9673# a_1591_9301# a_2455_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X857 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_12355_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X858 vccd1 a_24462_20149# a_24389_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X859 vssd1 _0472_.X _0574_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X861 vccd1 _0994_.CLK a_24775_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X862 a_4769_23145# _0740_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X863 _0969_.D a_23415_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X864 a_25639_12559# a_24941_12565# a_25382_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X865 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12355_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X866 vccd1 _0579_.C a_17539_16161# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X867 vccd1 a_26175_6005# a_26091_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X868 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X869 a_16968_21807# a_16569_21807# a_16842_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X870 vccd1 _0466_.A _0679_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X871 a_25214_12559# a_24775_12565# a_25129_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X872 vssd1 _0931_.CLK a_15483_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X873 a_4403_22869# _0788_.C a_4769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.585 ps=2.17 w=1 l=0.15
X874 a_14740_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X877 a_25589_19631# _1047_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X878 _0917_.CLK a_9411_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X879 a_5829_8527# _0710_.A1 a_5510_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X882 vccd1 _0994_.CLK a_25603_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X884 a_3326_2057# a_2752_1897# a_2956_1956# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X885 vssd1 fanout27.A a_16863_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X887 a_27517_5853# a_26983_5487# a_27422_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X889 _0987_.D a_9983_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X890 a_17562_1653# a_17394_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X891 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X892 _0713_.A1 _0745_.A3 a_5813_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X893 vssd1 a_23634_26677# a_23592_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X894 vccd1 _0582_.C a_21495_14219# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
R3 vccd1 temp1.capload\[2\].cap_47.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X895 _0602_.X a_18887_17024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X896 _0959_.CLK a_10423_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X897 vssd1 a_27847_5853# a_28015_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X899 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_15667_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X900 a_3321_26703# a_2787_26709# a_3226_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X901 vssd1 _0444_.A a_2787_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X902 a_8243_6031# a_7461_6037# a_8159_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X904 a_14917_23439# _1053_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X906 vssd1 a_25198_21919# a_25156_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X907 vccd1 _0502_.X a_20393_8545# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X908 a_25800_15113# a_25401_14741# a_25674_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X909 vssd1 a_25750_12127# a_25708_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X911 a_23975_17999# a_23193_18005# a_23891_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X916 vccd1 a_6427_11989# _0768_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X917 vssd1 _0994_.CLK a_25235_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X918 a_6821_6575# _0596_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X919 vccd1 a_4035_9813# _0698_.A1_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X921 a_23891_26703# a_23193_26709# a_23634_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X922 a_9436_16143# _0840_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 a_19973_17821# a_19439_17455# a_19878_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X924 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X925 a_7477_18319# _0737_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X926 a_15115_13103# _0471_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X930 vccd1 a_19689_9269# _0590_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X931 a_15128_23817# a_14729_23445# a_15002_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X932 a_4769_23145# _0847_.A3 a_4403_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X933 a_2823_3677# a_1959_3311# a_2566_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X934 a_25129_12559# _1000_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X935 vccd1 a_12467_10107# a_12383_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X937 a_5210_9001# _0734_.A2 a_5128_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X938 vccd1 _1022_.Q a_20214_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X939 a_10048_28111# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X940 a_17819_1679# a_17121_1685# a_17562_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X941 a_2030_9117# a_1591_8751# a_1945_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X942 _0696_.A1 _0734_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X944 a_2616_25071# a_2217_25071# a_2490_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X946 a_17861_1135# _0631_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X947 a_8746_7119# a_8473_7125# a_8661_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X948 a_25631_13469# a_24849_13103# a_25547_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X950 a_27337_15279# _0893_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X951 a_7164_14191# a_6938_14237# a_6795_14343# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X954 a_12502_3829# a_12334_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X956 _0670_.A2 a_16895_5281# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X957 vccd1 a_3819_26677# a_3735_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X958 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13360_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X959 fanout27.A a_16863_11479# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X960 a_27421_4399# a_26431_4399# a_27295_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X961 vssd1 a_2991_27515# a_2949_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X964 temp1.capload\[14\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X965 vccd1 _0821_.B a_10239_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X967 vssd1 _0572_.A2 a_24937_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X968 vssd1 a_17289_13249# _0605_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X969 a_9398_20175# _0761_.B a_9095_20407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X971 a_13437_16201# a_12447_15829# a_13311_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X972 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X973 a_22457_12559# _0891_.D a_22373_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X974 a_14725_19465# a_13735_19093# a_14599_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X976 a_9190_3829# a_9022_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X977 a_4548_2223# a_4149_2223# a_4422_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X978 a_8378_4943# a_7939_4949# a_8293_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X979 a_5796_19881# _0456_.B a_5724_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X980 a_6815_7913# _0657_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X981 vssd1 _0807_.B a_4537_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X983 vccd1 a_19275_21237# a_19191_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X984 a_2869_17501# _0722_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X985 a_22325_6603# _0504_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X986 a_16209_13103# _0521_.A a_16127_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X987 vssd1 _0549_.C1 a_16127_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X988 vssd1 _0863_.A1 a_15777_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X989 _0589_.X a_19439_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X991 vssd1 a_16182_4511# a_16140_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X992 vccd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_2686_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X994 a_2455_9295# a_1757_9301# a_2198_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X995 a_2313_1135# _0863_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X996 a_21230_10927# _1046_.D a_21140_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X997 vccd1 a_26578_11039# a_26505_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X998 a_5173_12265# a_4985_12061# a_5091_12021# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X999 vssd1 _0935_.CLK a_11343_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1001 vssd1 _0845_.A2 _0836_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 vssd1 a_10294_6005# a_10252_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1004 vssd1 _0689_.X _0694_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1007 vccd1 a_14341_15797# _0763_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1009 _0865_.Y _0864_.Y a_12725_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1010 a_4213_25223# _0844_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1011 a_11287_11293# a_10589_10927# a_11030_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1012 a_19878_15645# a_19439_15279# a_19793_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1013 vccd1 a_25455_5853# a_25623_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1014 a_5510_8527# _0734_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X1015 a_15170_23413# a_15002_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1018 vssd1 io_in[7] a_1591_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1019 a_3099_2767# a_2235_2773# a_2842_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1020 a_5215_2767# a_4351_2773# a_4958_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1021 vccd1 a_10903_2491# a_10819_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1022 a_7457_6575# a_6467_6575# a_7331_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1023 _0657_.X a_6416_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X1024 a_11509_20719# a_11343_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1025 a_10509_28335# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1026 a_4213_25223# _0844_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X1028 a_21598_15279# _1021_.Q a_21508_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1029 a_12502_3829# a_12334_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1031 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1032 a_21997_26159# a_21831_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1033 a_14563_16911# _1078_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1034 a_10478_2335# a_10310_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1035 a_4774_1653# a_4606_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1036 _0756_.A2 _0776_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1037 vccd1 _0444_.B a_11251_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1038 a_7625_14709# _0461_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1040 vccd1 a_16829_12161# _0565_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1041 a_24941_12565# a_24775_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1043 vccd1 _0827_.A a_11437_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1046 _0543_.B2 a_17895_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1047 vccd1 a_25750_12127# a_25677_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1049 vccd1 _0583_.C a_19195_18337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1052 a_5087_11791# _0708_.A2 a_4993_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1053 vccd1 a_3394_26677# a_3321_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1054 a_9190_3829# a_9022_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1055 vssd1 a_23599_7093# a_23557_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1057 vccd1 _0931_.CLK a_15483_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1058 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1059 a_6416_10089# _0778_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1060 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1062 a_9942_21263# a_9503_21269# a_9857_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1064 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1065 vccd1 _0456_.B _0722_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1067 a_12527_17455# _0472_.X _0751_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1068 vccd1 a_17895_3829# a_17811_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1071 a_25214_8207# a_24775_8213# a_25129_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1072 a_25674_7119# a_25401_7125# a_25589_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1073 a_20981_20553# a_19991_20181# a_20855_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1074 a_16548_10901# _0565_.B1 a_16940_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1075 vccd1 a_27590_16479# a_27517_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1076 vccd1 _0444_.B _0444_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 a_27337_7663# _1064_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1078 a_13897_10761# a_12907_10389# a_13771_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1079 a_3228_3145# a_2235_2773# a_3099_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X1080 vccd1 _0694_.A1 a_4934_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1081 _0622_.B2 a_10167_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1082 vccd1 _0935_.CLK a_12171_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1083 a_25999_17821# a_25217_17455# a_25915_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1084 a_7663_8527# _0475_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1085 a_1735_29941# _0845_.C1 a_2291_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1086 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1088 a_17404_12015# _0565_.A1 a_16829_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X1089 _1011_.D a_26267_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1090 a_11697_15279# _0988_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1091 a_3324_14441# _0722_.B a_3240_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1092 _0698_.A2_N _0699_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1093 _0816_.S _0444_.B a_9687_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 a_2030_6941# a_1757_6575# a_1945_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1096 vccd1 a_13035_21263# a_13203_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1097 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1098 vssd1 _0931_.CLK a_20911_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1099 _0630_.A2 _0474_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1100 a_21407_4765# a_20709_4399# a_21150_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1101 a_11251_24233# _0825_.A1 _0825_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1102 vssd1 fanout27.A a_22659_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1104 a_17323_2223# _0516_.B1 a_17501_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1105 a_5361_30287# _0809_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1106 vssd1 a_13035_21263# a_13203_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1107 vssd1 clkbuf_1_0__f_io_in[0].X a_1775_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1108 a_10325_10703# _0466_.A a_10107_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1109 a_18288_18543# _0577_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X1110 a_6817_5487# a_6651_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1111 a_2156_8751# a_1757_8751# a_2030_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1112 _0890_.D a_12467_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1114 a_8305_19087# _0813_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1115 vssd1 _0768_.B1 a_7111_13655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1116 a_22963_20175# a_22181_20181# a_22879_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1117 a_25125_16733# a_24591_16367# a_25030_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1118 vccd1 a_23855_15831# _0964_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1119 _0695_.A1 _0686_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1120 _0835_.A1 a_2626_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1121 vccd1 _0972_.CLK a_19163_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1123 a_16784_26159# a_16385_26159# a_16658_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1124 a_25842_15797# a_25674_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1125 vssd1 a_22879_1679# a_23047_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1127 a_17217_3855# _0671_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1128 vssd1 a_17657_13621# _0609_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X1129 a_23381_17999# _0963_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1131 a_4973_28335# a_3983_28335# a_4847_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1132 _0869_.Y _0869_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1133 a_23465_9839# _1069_.Q a_23119_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1135 a_2686_15823# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1136 a_15671_7235# a_15565_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1137 _0439_.A a_2623_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1138 _0707_.A1 _0655_.X a_5357_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1140 a_16048_20719# a_15649_20719# a_15922_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1141 vssd1 _0774_.A2 a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X1142 vssd1 a_4590_2335# a_4548_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1143 a_8504_5321# a_8105_4949# a_8378_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1144 vccd1 _0582_.A a_19439_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1146 a_25674_15823# a_25401_15829# a_25589_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1147 a_21729_7913# _0516_.B1 a_21813_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 a_14373_32463# temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1150 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1151 a_24469_10749# _0573_.B a_24397_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1154 a_9558_16885# a_9390_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1155 vccd1 ANTENNA_7.DIODE a_25789_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X1156 vccd1 a_20303_15645# a_20471_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1157 a_21533_3311# a_20543_3311# a_21407_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1158 a_4790_2767# a_4351_2773# a_4705_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1159 vccd1 _0842_.A0 a_14195_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1160 vccd1 a_12610_21807# a_12716_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1161 vccd1 a_16929_17973# _0522_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1162 a_22580_16201# a_22181_15829# a_22454_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1163 vssd1 a_4035_9813# _0698_.A1_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1164 a_12318_11445# a_12150_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1165 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8767_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1167 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1168 a_27590_15391# a_27422_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1169 vssd1 _0527_.X a_21213_11809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1170 _0787_.X a_6600_27907# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1171 _0591_.X a_14655_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1172 a_21442_13469# a_21003_13103# a_21357_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1174 a_27337_12015# _1013_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1175 _1022_.Q a_22587_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1177 a_9390_16911# a_9117_16917# a_9305_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1179 a_6559_27023# _0814_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 a_19773_18689# _0583_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X1181 a_27973_2223# a_26983_2223# a_27847_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1182 a_2823_3677# a_2125_3311# a_2566_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1183 a_24757_2223# a_24591_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1185 _0847_.A3 a_10055_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1186 a_9999_5853# a_9301_5487# a_9742_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1187 vccd1 _0438_.A a_8135_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1188 a_23607_9117# a_22825_8751# a_23523_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1189 a_27847_14557# a_26983_14191# a_27590_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1190 a_27038_4511# a_26870_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1191 vccd1 a_6608_29111# _0825_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_2113_23983# _0444_.A a_1585_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.10725 ps=0.98 w=0.65 l=0.15
X1193 vccd1 _1015_.CLK a_26983_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1196 _0527_.X a_14603_15325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X1197 vssd1 a_23691_4667# a_23649_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1198 vssd1 a_3891_21263# _0814_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1200 a_25800_19631# a_25401_19631# a_25674_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1201 vccd1 a_9447_3855# a_9615_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1202 vssd1 _0975_.CLK a_24591_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1203 a_13035_21263# a_12171_21269# a_12778_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1204 a_11509_20719# a_11343_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1206 vssd1 _0931_.CLK a_16771_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1207 a_24535_11471# a_23837_11477# a_24278_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1208 a_14813_14013# _1076_.Q a_14741_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X1209 a_3099_2767# a_2401_2773# a_2842_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X1210 vssd1 _0764_.A1 a_6600_27907# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1211 _0563_.B1 a_20299_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1213 a_14557_14191# a_14287_14557# a_14453_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1214 _0491_.X a_11929_9633# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X1215 vccd1 _0684_.A1 a_8478_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1216 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1218 vssd1 a_15427_3855# a_15595_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1219 _0902_.Q a_10719_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1220 vssd1 a_9095_10615# _0597_.A2_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1221 a_21867_24349# a_21169_23983# a_21610_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1222 _0584_.C1 a_22015_18112# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1223 vccd1 a_13771_22351# a_13939_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1224 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_6191_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1225 a_13901_19093# a_13735_19093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1226 vssd1 _0860_.B _0856_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1227 a_25340_8585# a_24941_8213# a_25214_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1229 a_20349_6825# _0548_.B2 a_20267_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1230 vssd1 _0776_.A2 a_4340_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1231 vccd1 _0444_.Y a_5273_29687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X1233 _0605_.C1 a_17783_12672# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1235 _0667_.B1 a_18001_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1236 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1237 a_5727_7119# _0686_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1238 a_17727_3855# a_17029_3861# a_17470_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1239 a_11877_11477# a_11711_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1240 vssd1 _0529_.Y a_22169_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1241 a_10968_31375# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1242 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13183_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1243 vssd1 a_1735_29941# _0847_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 a_25582_3677# a_25143_3311# a_25497_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1245 vccd1 _0505_.A2 a_20993_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1247 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1249 a_26417_20719# _0966_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1250 _0576_.B1 a_24315_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1251 a_20525_22351# a_19991_22357# a_20430_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1252 vssd1 a_25455_5853# a_25623_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1253 vssd1 clkbuf_1_0__f_io_in[0].X a_1591_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1254 a_7623_10901# _0546_.X a_7850_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X1255 a_22948_19465# a_22549_19093# a_22822_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1256 a_22546_2767# a_22273_2773# a_22461_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1257 vccd1 _0685_.B a_7653_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1260 vccd1 a_25198_16479# a_25125_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1261 _0677_.A1 a_6487_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1262 _0649_.B2 a_20563_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1263 _0679_.A2 _0475_.X a_7745_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1265 a_27548_21807# a_27149_21807# a_27422_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1266 a_20237_16189# _0930_.Q a_20165_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1267 vssd1 a_15595_23413# a_15553_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1268 a_4403_22869# _0809_.B2 a_4959_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 vccd1 _0456_.A a_5243_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1271 vccd1 _0794_.A2 a_6741_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1272 vssd1 a_11435_22895# _0847_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1273 vssd1 _0999_.CLK a_26063_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1274 vccd1 a_2991_3579# a_2907_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1275 a_16258_18793# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1276 vssd1 a_10386_4917# a_10344_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1279 a_9945_1685# a_9779_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1280 a_20782_5599# a_20614_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1281 vssd1 a_2198_8863# a_2156_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1283 a_27422_14557# a_27149_14191# a_27337_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1284 vccd1 a_5015_2491# a_4931_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1285 vssd1 a_25842_1247# a_25800_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1286 vccd1 a_8914_7093# a_8841_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1287 vccd1 a_22015_8215# _1033_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1288 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1289 a_1585_24135# _0765_.B1 a_1916_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
X1291 a_20046_17567# a_19878_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1292 a_19878_15645# a_19605_15279# a_19793_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1293 a_15001_3087# _0959_.D a_14655_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1294 vssd1 a_9742_1247# a_9700_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1295 _0815_.Y _0825_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1296 a_27330_9117# a_27057_8751# a_27245_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1297 a_18505_20175# _1049_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1298 a_21831_10089# _0666_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1299 _0512_.A a_19439_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1300 a_4931_1501# a_4149_1135# a_4847_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1301 vccd1 _0908_.CLK a_3799_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1302 vccd1 clkbuf_1_0__f_io_in[0].X a_1683_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1303 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1304 vccd1 fanout10.A a_10147_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1306 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1308 a_24941_8213# a_24775_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1311 a_20982_3677# a_20709_3311# a_20897_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1313 a_7636_29967# a_7387_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1315 a_4251_11249# _0698_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.335 w=0.64 l=0.15
X1316 a_12935_12879# a_12643_12559# a_12849_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1317 a_2693_15543# _0722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1318 a_14726_10205# a_14287_9839# a_14641_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1322 vccd1 a_17727_2767# a_17895_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1323 a_25658_8863# a_25490_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1324 vssd1 a_26670_20831# a_26628_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1325 vccd1 a_10055_23983# _0847_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1326 a_2962_14735# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1327 a_20083_19200# _1019_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1328 a_24757_15279# a_24591_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1330 a_16983_12897# _0583_.A a_16897_12897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1331 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1332 a_27931_8029# a_27149_7663# a_27847_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1333 a_26877_13103# _1066_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1334 a_6369_22057# _0797_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1335 a_26854_18655# a_26686_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1336 vccd1 a_27847_17821# a_28015_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1338 a_4916_3145# a_4517_2773# a_4790_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1339 vccd1 a_2198_6687# a_2125_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1340 a_21279_6825# _0630_.A2 a_21361_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1341 a_22227_2589# a_21445_2223# a_22143_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1342 _0662_.A1 a_18611_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1343 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A _0816_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1344 vccd1 a_27571_6941# a_27739_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1345 a_23385_10703# _0621_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1347 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1348 vccd1 a_26210_26271# a_26137_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1349 a_5047_21781# _0727_.A1 a_5329_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X1351 vccd1 _0768_.A1 a_10693_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X1352 a_3154_24893# _0860_.A a_2655_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X1355 a_14913_14741# a_14747_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1358 _0538_.C1 a_11251_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1359 vssd1 _0994_.CLK a_25603_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1360 a_27931_25437# a_27149_25071# a_27847_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1361 a_27590_14303# a_27422_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1363 a_5128_9001# _0734_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1364 a_3141_26703# _0835_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1365 vssd1 _0807_.A a_5547_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1366 a_15462_16733# a_15023_16367# a_15377_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1367 vccd1 a_5383_2741# a_5299_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1368 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1369 _0475_.X a_11815_12265# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X1370 vccd1 _0583_.C a_20083_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1371 vssd1 _0658_.B1 a_16565_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1373 vssd1 fanout24.A a_22015_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1374 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1376 vssd1 a_26578_11039# a_26536_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1381 a_27590_9951# a_27422_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1382 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1384 vssd1 _0994_.CLK a_26983_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1386 a_22622_16885# a_22454_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1387 a_11233_14441# _0860_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1388 a_21476_18543# a_21077_18543# a_21350_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1389 _0516_.B1 a_18645_7457# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1390 a_12659_11471# a_11877_11477# a_12575_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1392 a_10041_6031# _0901_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1393 a_7435_26324# _0817_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1394 a_15016_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1395 a_15197_5059# _0556_.D a_15115_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1396 _0608_.X a_20083_15936# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1397 vssd1 a_28015_15547# a_27973_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1400 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1402 vssd1 _0584_.A2 a_20348_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1403 _0439_.A a_2623_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1404 a_12123_27069# _0825_.A1 a_11760_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1405 vccd1 a_24719_1679# a_24887_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1406 _0861_.B1 a_3799_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1407 vssd1 _0812_.A2 a_10147_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1408 a_4165_14455# _0456_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1410 a_22879_16911# a_22181_16917# a_22622_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1411 a_10413_17999# _0797_.A1 a_10331_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1414 a_9769_19631# _0751_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1415 vccd1 _1075_.Q a_13257_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X1417 _0444_.B a_11803_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1418 vssd1 _0440_.A _0872_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1419 a_22454_16911# a_22015_16917# a_22369_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1420 a_22454_16911# a_22181_16917# a_22369_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1421 a_11333_5487# _0986_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1422 a_14910_17999# a_14471_18005# a_14825_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1423 vssd1 fanout27.A a_19807_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1425 a_22545_21807# a_21555_21807# a_22419_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1428 vccd1 a_25842_7093# a_25769_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1429 vccd1 _0508_.Y a_12355_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X1430 vssd1 _0778_.A2 _0680_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1431 _0489_.X a_19531_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1432 vccd1 a_20598_22325# a_20525_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1433 vssd1 a_14767_19061# a_14725_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1435 vccd1 _0964_.CLK a_23027_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1436 _1069_.Q a_26175_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1437 _0512_.A a_19439_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1438 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1439 a_25708_3311# a_25309_3311# a_25582_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1440 a_27590_2335# a_27422_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1441 a_14603_15325# _1075_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1442 vssd1 a_10443_4667# a_10401_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1444 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1446 a_17865_9845# _0624_.D_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1447 vssd1 _0972_.CLK a_15575_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1448 a_23657_6031# _0607_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1449 vssd1 a_12743_11445# a_12701_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1450 vssd1 a_12631_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1452 a_8841_7119# a_8307_7125# a_8746_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1455 a_25915_8029# a_25051_7663# a_25658_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1457 a_15088_29673# a_14839_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1458 vssd1 _0515_.B1 a_21073_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1459 vssd1 a_26175_6005# a_26133_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1460 a_10107_10615# _0466_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X1462 a_18371_1501# a_17673_1135# a_18114_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1467 vssd1 a_10643_4943# a_10811_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1468 vssd1 a_22438_26271# a_22396_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1469 a_23385_16617# _0929_.Q a_23303_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1470 a_10037_2223# a_9871_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1471 a_15565_7235# _0642_.D_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1472 _0941_.Q a_21851_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1473 vssd1 a_12242_27791# a_12348_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1474 vssd1 _0513_.X a_13395_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1475 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1476 a_5525_4399# a_4535_4399# a_5399_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1477 _0613_.A1 a_10351_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 vccd1 io_in[0] a_2962_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1479 a_22737_1135# _0967_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1483 a_4902_25981# _0840_.A1 a_4403_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X1484 _0596_.A1 a_5659_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1485 a_15151_8029# a_14453_7663# a_14894_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1486 a_12356_19203# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1487 a_15841_9001# _0595_.D a_15759_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1488 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_7636_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1490 vssd1 a_2381_16885# _0875_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1491 a_27146_6941# a_26707_6575# a_27061_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1494 a_20341_5487# a_20175_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1495 vccd1 _0695_.A1 a_4439_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1496 a_2455_9295# a_1591_9301# a_2198_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1497 _0891_.D a_22035_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1498 vccd1 _0999_.CLK a_26063_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1499 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1500 a_21683_9117# a_20985_8751# a_21426_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1501 vssd1 _0893_.CLK a_26523_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1502 a_2125_6941# a_1591_6575# a_2030_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1503 vccd1 _0533_.X a_13717_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X1505 a_19402_1653# a_19234_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1506 a_23910_6005# a_23742_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1507 a_23565_21263# _1048_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1508 _0803_.X a_6283_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1509 vccd1 _0532_.A2 a_11693_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X1510 vssd1 _1019_.CLK a_19163_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1513 a_4451_7913# a_4259_7669# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1514 a_10120_27791# a_9871_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1515 _0552_.B2 a_28015_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1516 vssd1 _1030_.CLK a_15667_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1517 vssd1 _0778_.A2 a_6087_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X1518 vssd1 a_27590_24095# a_27548_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1519 a_14852_9839# a_14453_9839# a_14726_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1521 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1522 vssd1 clkbuf_1_0__f_io_in[0].X a_2235_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1523 a_17336_19631# a_16937_19631# a_17210_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1524 a_22990_19061# a_22822_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1525 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_12316_24135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1528 vccd1 _1053_.CLK a_10791_16919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1530 a_22120_21807# a_21721_21807# a_21994_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1531 vccd1 a_1867_15831# _0722_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1532 a_17854_3677# a_17581_3311# a_17769_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1533 vccd1 a_21345_15253# _0542_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1535 a_11874_10205# a_11601_9839# a_11789_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1537 a_22659_10927# _0648_.B1 a_22837_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1538 a_16385_26159# a_16219_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1539 vssd1 a_7499_6843# a_7457_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1540 a_9945_4765# a_9411_4399# a_9850_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1542 a_22990_14303# a_22822_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1543 a_9497_13353# _0746_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1544 _0890_.D a_12467_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1545 vssd1 a_9095_20407# _0459_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1546 vssd1 a_19770_26677# a_19728_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1547 a_15005_17999# a_14471_18005# a_14910_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1548 a_18850_21237# a_18682_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1549 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1550 vssd1 a_22143_2589# a_22311_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R4 temp1.capload\[0\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1551 a_4337_2223# _0865_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1552 _0894_.Q a_26175_12283# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1553 vccd1 a_27498_8863# a_27425_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1554 vccd1 _0931_.CLK a_19439_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1555 a_10643_2767# a_9945_2773# a_10386_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1556 vssd1 io_in[4] a_1591_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1557 a_5245_12265# _0711_.B a_5173_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X1558 a_4548_26159# a_4149_26159# a_4422_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1559 a_2858_25615# a_2419_25621# a_2773_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1560 a_11936_17027# _0813_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1561 vssd1 a_21575_3579# a_21533_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1562 a_2398_2589# a_1959_2223# a_2313_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1566 a_19770_3829# a_19602_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1567 _0850_.A a_3270_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X1568 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1569 a_3333_19407# _0872_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1570 a_6440_29673# a_6191_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1571 vccd1 _0583_.C a_18887_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1572 a_25674_25615# a_25235_25621# a_25589_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1573 vssd1 clkbuf_1_1__f__0390_.A a_2686_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1574 a_23423_21085# a_22641_20719# a_23339_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 a_12801_2767# _0946_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1576 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12355_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1578 a_18682_21263# a_18409_21269# a_18597_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1579 a_7288_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1580 a_22695_26525# a_21831_26159# a_22438_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1582 a_24803_1679# a_24021_1685# a_24719_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1583 _0576_.D1 a_22015_6144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1585 a_22929_7663# _0618_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X1586 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1587 a_5215_2767# a_4517_2773# a_4958_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1588 a_13735_12925# _0602_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X1589 vccd1 a_4035_13077# _0780_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1590 vssd1 a_22622_15797# a_22580_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1591 a_23331_19087# a_22549_19093# a_23247_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1592 vssd1 a_4774_1653# a_4732_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1593 vccd1 a_20671_8029# a_20839_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1594 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1597 a_19202_15823# _0582_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X1600 a_22365_26525# a_21831_26159# a_22270_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1601 vccd1 a_20027_26703# a_20195_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1602 vssd1 a_28015_14459# a_27973_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1603 a_17489_2473# _0956_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1604 _0740_.X a_6600_26409# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X1606 a_11776_28585# a_11527_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1610 temp1.capload\[0\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1611 a_2907_2589# a_2125_2223# a_2823_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1612 vssd1 _0808_.A a_8123_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1613 vssd1 a_2991_1403# a_2949_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1615 vssd1 _0861_.A2 a_16208_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1617 _0639_.X a_13735_3968# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1619 a_11983_22351# _0858_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1620 vssd1 a_25750_3423# a_25708_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1621 a_19531_11471# _0648_.A2 a_19709_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1622 a_26225_17289# a_25235_16917# a_26099_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1623 a_15563_9295# _0652_.C a_15369_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1625 a_17302_2767# a_16863_2773# a_17217_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1626 vssd1 a_13459_8751# _0521_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1629 vccd1 _0643_.B1 a_25309_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X1630 vccd1 a_10643_1679# a_10811_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1633 _0745_.A3 _0776_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1634 a_10396_30761# a_10147_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1635 a_25382_23413# a_25214_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1636 _1060_.D a_18079_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1637 a_10110_11445# a_9942_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1638 _0558_.A2 a_21127_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1639 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1640 a_9643_25398# _0825_.A1 a_9184_25223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1641 vssd1 a_16548_10901# _0616_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1642 vssd1 a_18850_21237# a_18808_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1643 a_19770_3829# a_19602_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1644 vccd1 a_22714_2741# a_22641_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1645 a_22449_15253# _0648_.B1 a_22606_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1646 a_25030_4765# a_24757_4399# a_24945_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1647 a_15833_12559# _0990_.D a_15749_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1648 a_15538_1653# a_15370_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1649 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1650 vccd1 a_15576_21379# _0863_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1652 _0584_.A2 a_15607_15307# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1653 a_2217_3855# a_1683_3861# a_2122_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1654 vssd1 _0702_.B1_N a_4259_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X1655 vssd1 _0935_.Q a_9436_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X1658 fanout37.A a_3523_6039# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1659 a_4262_13103# _0758_.A1 a_4035_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X1660 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14011_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1661 _0933_.Q a_18263_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1662 a_13729_6351# _0538_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X1663 a_27272_6575# a_26873_6575# a_27146_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1666 vssd1 _0959_.CLK a_14747_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1668 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10120_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1669 a_26168_26159# a_25769_26159# a_26042_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1670 a_10551_6031# a_9853_6037# a_10294_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1672 a_19298_16143# _1023_.Q a_19208_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1673 vccd1 clkbuf_1_0__f_io_in[0].X a_3983_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1674 vccd1 _1015_.CLK a_25143_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1675 a_18045_11471# _0897_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1676 a_18225_17999# _1018_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1677 vssd1 _0628_.X a_17473_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X1678 a_10727_1679# a_9945_1685# a_10643_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1679 a_25723_8207# a_24941_8213# a_25639_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1680 a_23381_26703# _0994_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1681 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1684 vccd1 a_28015_12283# a_27931_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1685 a_25547_13469# a_24683_13103# a_25290_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1686 vssd1 _0847_.A3 a_13080_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1687 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1689 vssd1 a_14894_9951# a_14852_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1690 a_10133_4943# _0952_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1691 a_1945_5487# _0880_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1692 vccd1 a_18025_7809# _0634_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1693 vssd1 a_5601_18517# _0784_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1694 a_4621_11249# _0807_.B a_4040_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X1695 _0665_.B2 a_25623_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1697 a_21065_16189# _0995_.Q a_20993_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1698 a_25589_1135# _0552_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1699 vccd1 a_20690_21237# a_20617_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1700 vccd1 _0518_.Y a_15607_15307# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1701 a_27425_9117# a_26891_8751# a_27330_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1702 a_9489_1135# _0646_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1704 a_11987_4943# _0535_.X a_12069_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1705 _0711_.B _0710_.B1 a_5445_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1707 vssd1 _0523_.X a_14011_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1708 a_15795_1679# a_15097_1685# a_15538_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1709 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10876_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1711 a_12613_2773# a_12447_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1713 a_18409_9001# _0897_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1714 _0824_.Y temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1716 a_25143_14441# _0648_.A2 a_25225_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1717 a_24845_22729# a_23855_22357# a_24719_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1718 a_24301_2767# _1034_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1719 vccd1 temp1.capload\[10\].cap.A temp1.capload\[10\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1720 _0995_.CLK a_9227_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1721 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1722 a_5142_4511# a_4974_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1723 a_16105_12879# _0918_.D a_15667_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1725 a_19899_1385# _0516_.B1 a_19981_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1727 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_6440_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1728 vssd1 _0444_.B _0819_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X1729 a_12575_8207# a_11877_8213# a_12318_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1730 vccd1 _0975_.CLK a_23855_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1731 a_5066_4943# a_4793_4949# a_4981_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1732 vssd1 _0487_.X a_18681_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1733 vccd1 a_14433_24501# _0852_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1734 vssd1 a_10110_11445# a_10068_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1735 a_12643_12559# _0836_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X1736 a_2125_3311# a_1959_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1737 vccd1 _0861_.B1 a_4981_21024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X1738 _0966_.D a_24887_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1739 a_2524_2223# a_2125_2223# a_2398_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1740 vccd1 a_25807_12533# a_25723_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1741 a_27973_17455# a_26983_17455# a_27847_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1743 a_1674_32143# clkbuf_1_1__f_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1744 _0643_.X a_22291_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1745 temp1.capload\[6\].cap.Y temp1.capload\[6\].cap_51.LO a_14373_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1746 vssd1 _1079_.Q _0479_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1747 a_11877_18909# a_11343_18543# a_11782_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1748 a_19605_4649# _0497_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1749 vssd1 _0844_.B a_4534_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X1750 _0966_.D a_24887_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1751 vssd1 clkbuf_1_0__f_io_in[0].X a_1591_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1753 _0739_.A2 a_6559_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1754 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1755 _1080_.Q a_3083_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1756 vccd1 a_22438_26271# a_22365_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1757 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10140_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1758 _0866_.Y _0866_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1759 a_20345_22351# _0932_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1760 a_17719_19997# a_16937_19631# a_17635_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1762 _0572_.D1 a_23303_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1763 a_25639_23439# a_24941_23445# a_25382_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1764 a_13449_6575# _0521_.A a_13367_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1765 a_16569_21807# a_16403_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1766 a_13257_17821# a_13091_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X1767 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1769 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11776_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1770 vccd1 _0844_.B a_4547_25393# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1771 a_25214_23439# a_24775_23445# a_25129_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1772 vssd1 a_25198_15391# a_25156_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1773 a_27167_10383# _0619_.B1 a_27249_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1774 vssd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_1766_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1775 vccd1 a_26175_3579# a_26091_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1776 vccd1 a_17657_13621# _0609_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1778 a_7348_17973# _0813_.A2 a_7571_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1779 a_2710_1679# a_2114_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.1218 ps=1.42 w=0.42 l=0.15
X1780 a_15841_1385# _0946_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1783 vccd1 _0722_.C a_3983_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1784 a_27088_13103# a_26689_13103# a_26962_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1785 a_25122_13469# a_24849_13103# a_25037_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1786 vssd1 _0893_.CLK a_24775_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1789 a_22641_2767# a_22107_2773# a_22546_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1791 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10396_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1792 a_13897_22729# a_12907_22357# a_13771_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1794 _0835_.Y _0833_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1796 vssd1 a_10202_18517# _0577_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1797 a_8105_4949# a_7939_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1798 vccd1 a_2655_24501# _0839_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X1800 a_17428_3145# a_17029_2773# a_17302_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1801 a_20543_9839# _1025_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1802 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12539_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1803 _0646_.A1 a_6947_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1804 _0672_.C1 a_14747_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1807 _0627_.X a_20911_15936# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1809 a_24420_22729# a_24021_22357# a_24294_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1812 a_24294_1679# a_23855_1685# a_24209_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1813 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1814 a_19531_16367# _0522_.B1 a_19709_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1815 a_6427_11989# _0745_.A2 a_6645_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X1816 _0444_.Y _0444_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1817 a_13889_4221# _0639_.B a_13817_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1818 a_4365_13103# _0791_.A3 a_4262_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X1819 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1820 a_4729_26703# _0845_.C1 _0835_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1823 _0908_.Q a_8235_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1825 a_25842_4917# a_25674_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1826 vccd1 _1019_.CLK a_21003_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1828 vccd1 a_22325_6603# _0619_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X1829 a_2686_10383# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1830 vccd1 _1033_.CLK a_24775_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1833 a_6905_2223# a_5915_2223# a_6779_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1834 vccd1 a_25382_12533# a_25309_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1836 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1837 _0582_.C a_14729_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X1838 a_16293_7913# _0549_.B2 a_16209_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1839 a_25129_23439# _0995_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1841 vssd1 _0722_.A _0456_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1842 vssd1 a_27314_6687# a_27272_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
R5 vccd1 temp1.capload\[10\].cap_40.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1846 a_24068_12559# _0643_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1847 a_2217_25071# a_2051_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1848 a_25198_16479# a_25030_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1849 vssd1 _1062_.CLK a_18611_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1850 a_27337_3311# _1069_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1851 vccd1 _0959_.CLK a_9779_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1852 vccd1 _0582_.C a_20543_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1853 a_4581_25847# _0844_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X1854 a_5245_21807# _0723_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1855 vssd1 a_14341_17429# _0773_.A2_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1856 a_23361_13249# _0569_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1857 _0471_.X a_9503_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1858 a_9497_14735# _0735_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1859 a_5445_9295# _0710_.B2 _0711_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1860 a_24113_2773# a_23947_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1861 a_17497_5737# _0622_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1862 a_9301_5487# a_9135_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1864 a_26041_7663# a_25051_7663# a_25915_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1865 vccd1 a_7896_11703# _0734_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1866 a_22879_20175# a_22015_20181# a_22622_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1867 a_2686_15823# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1868 vccd1 _0521_.A a_16863_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1871 a_17029_2773# a_16863_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1872 vssd1 _0774_.A2 a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1874 a_25455_15645# a_24591_15279# a_25198_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1875 vccd1 clkbuf_1_0__f_io_in[0].X a_3983_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1876 a_24570_13647# a_24131_13653# a_24485_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1877 a_13984_31055# a_13735_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1879 vssd1 a_26486_23007# a_26444_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1880 a_18421_8751# _0987_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X1881 a_9495_11249# _0597_.A2_N a_9494_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X1883 vssd1 _1078_.Q a_14287_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X1884 a_14661_6825# _0901_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1887 a_22921_7119# _1045_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1888 a_5357_10927# _0685_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1889 a_22549_20175# a_22015_20181# a_22454_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1890 vccd1 a_25198_4511# a_25125_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1893 a_19439_10496# _0607_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1894 a_12759_3855# a_12061_3861# a_12502_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1895 _0975_.CLK a_22015_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1896 vccd1 a_20138_2741# a_20065_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1897 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1898 a_4612_25981# a_4581_25847# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X1899 a_26099_1501# a_25235_1135# a_25842_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1900 a_8122_10927# _0546_.X a_7623_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X1902 a_20303_15645# a_19605_15279# a_20046_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1903 _0916_.D a_10167_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1904 _0606_.X a_16863_14848# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1905 a_19521_4649# _0496_.X a_19439_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1906 a_25842_4917# a_25674_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1907 a_3049_4943# _0673_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1908 _0941_.Q a_21851_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1909 vssd1 a_21683_19997# a_21851_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1910 a_14917_3855# _0954_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1911 vssd1 a_15335_17999# a_15503_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1912 _0579_.C a_13257_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1914 a_23610_13353# _0572_.D1 a_23361_13249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X1916 vccd1 _0657_.X a_6815_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X1917 a_23649_16367# _0966_.D a_23303_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1918 a_6741_14735# _0794_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1919 vssd1 a_2566_2335# a_2524_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1920 a_9447_3855# a_8749_3861# a_9190_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1921 vccd1 _0935_.CLK a_15023_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1922 vccd1 a_23523_4765# a_23691_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1923 vssd1 _0508_.Y a_14012_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X1924 vccd1 a_22419_22173# a_22587_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1925 vssd1 a_1639_7338# input2.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1927 a_7641_5487# a_6651_5487# a_7515_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1928 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE a_9871_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1929 a_25589_3855# _1072_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1930 a_23098_4765# a_22659_4399# a_23013_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1932 vccd1 a_23415_14459# a_23331_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1933 vccd1 _0504_.A a_20911_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1934 a_14737_3087# _0952_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1938 a_6641_19631# _0807_.A a_6559_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1939 _0533_.X a_16897_12897# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1941 a_20027_3855# a_19163_3861# a_19770_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1942 _0665_.B2 a_25623_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1945 a_24849_13103# a_24683_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1947 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1948 a_4149_26159# a_3983_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1949 a_24941_23445# a_24775_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1950 a_16569_21807# a_16403_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1951 a_18129_15279# _0932_.D a_17691_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1953 vccd1 _0681_.X a_5902_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1954 _0546_.A2 _0466_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1955 vccd1 a_3083_28603# a_2999_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1956 a_14269_20181# a_14103_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1957 a_25674_15823# a_25235_15829# a_25589_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1958 vccd1 _0585_.X a_16009_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1959 vccd1 _0845_.A1 a_7197_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X1962 a_12805_3561# _0910_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1963 a_10294_6005# a_10126_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1964 a_11874_10205# a_11435_9839# a_11789_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1965 vccd1 _0596_.A1 a_9398_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1966 vccd1 temp1.capload\[3\].cap.A temp1.capload\[3\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1967 vssd1 a_14307_4917# a_14265_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1968 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13183_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1969 _0966_.Q a_27095_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1970 _0708_.A3 a_4451_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X1971 a_19429_8207# _1016_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1972 a_8116_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1975 vccd1 a_4772_13621# _0794_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1976 vssd1 a_5567_4667# a_5525_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1977 a_4468_13103# _0791_.A2 a_4365_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X1978 a_13514_22325# a_13346_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1979 vssd1 a_16515_20987# a_16473_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1980 a_6906_6941# a_6633_6575# a_6821_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1981 vccd1 a_6613_22325# _0868_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1982 vccd1 _0807_.C a_8155_16161# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
D0 vssd1 _0863_.Y sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1983 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1984 vccd1 _0935_.CLK a_13735_19093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1985 a_25800_19465# a_25401_19093# a_25674_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1986 _0856_.Y _0860_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1988 vccd1 _0696_.A1 a_4530_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X1989 a_9496_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1990 vssd1 a_19770_3829# a_19728_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1991 a_23247_1501# a_22549_1135# a_22990_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1993 a_4300_17027# _0872_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1994 vssd1 a_17895_10357# a_17853_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1995 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1996 a_24420_2057# a_24021_1685# a_24294_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1997 a_11895_1385# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1998 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1999 a_6498_24233# _0764_.A1 a_6416_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2000 a_19970_2767# a_19697_2773# a_19885_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2001 vssd1 _0662_.A1 a_11815_12265# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X2002 vssd1 a_22817_18517# _0662_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X2003 vccd1 _0695_.A2 a_4015_5515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2005 a_17946_1501# a_17673_1135# a_17861_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2006 a_12604_28585# a_12355_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2007 a_25497_3311# _0505_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
R6 temp1.capload\[7\].cap_52.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2008 vssd1 a_21279_22895# _0994_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 a_9781_10927# _0840_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2010 vssd1 a_9171_7119# a_9339_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2011 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2013 vssd1 _0589_.X a_15759_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2015 a_21717_27247# a_20727_27247# a_21591_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2016 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2017 io_out[1] a_4403_22869# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2018 a_20073_5309# _0582_.A a_19991_5056# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2021 a_13633_14013# _0521_.A a_13551_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2022 a_3435_17231# _0456_.A a_3298_17143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2023 vccd1 _0964_.CLK a_24591_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2024 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2025 _0552_.B2 a_28015_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2026 vssd1 fanout24.A a_16035_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2027 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2028 a_5724_31599# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2029 vccd1 a_3283_25615# a_3451_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2032 a_11224_30761# a_10975_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2033 a_16385_26159# a_16219_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2034 a_25125_4765# a_24591_4399# a_25030_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2035 _0837_.Y _0845_.C1 a_6937_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2036 a_25957_26159# _0994_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2038 a_11782_15645# a_11343_15279# a_11697_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2039 a_20065_2767# a_19531_2773# a_19970_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2040 a_13337_7485# _0611_.B a_13265_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2041 a_15661_11177# _0609_.X a_15565_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2042 vccd1 a_1591_16367# _0722_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2043 vssd1 a_2956_1956# a_2885_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0989 ps=0.995 w=0.64 l=0.15
X2044 vssd1 a_3283_25615# a_3451_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2045 vssd1 _0784_.A2 a_7376_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2048 a_14729_3861# a_14563_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2049 a_12763_12879# a_12447_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2050 _0610_.X a_13551_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2052 a_10091_8029# a_9227_7663# a_9834_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2053 _0686_.X a_6653_10933# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X2054 vssd1 _0931_.CLK a_19439_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2055 a_26091_12381# a_25309_12015# a_26007_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2056 a_10714_20541# _0773_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2057 a_2398_1501# a_2125_1135# a_2313_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2058 a_24021_1685# a_23855_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2059 a_24389_1679# a_23855_1685# a_24294_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2060 vssd1 a_26854_18655# a_26812_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2061 vssd1 _0722_.B _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2063 vccd1 _0791_.A2 a_5821_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2064 a_2885_2057# a_2762_1801# a_2464_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0657 ps=0.725 w=0.36 l=0.15
X2066 a_10310_2589# a_10037_2223# a_10225_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2067 vssd1 _0680_.Y a_5817_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X2068 a_9255_7119# a_8473_7125# a_9171_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2069 _0662_.A1 a_18611_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2071 a_14726_8029# a_14453_7663# a_14641_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2073 vssd1 a_9189_18517# _0782_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2074 a_6522_2335# a_6354_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2075 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2076 vssd1 a_26267_16885# a_26225_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2078 _0570_.X a_23303_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2079 a_5725_17027# _0807_.A a_5629_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2080 a_14641_9839# _0961_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2081 a_21357_13103# _0890_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2082 vssd1 _1078_.Q a_14729_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X2083 vccd1 a_5234_4917# a_5161_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2085 a_5165_19087# a_4988_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2086 vccd1 _0533_.X a_23385_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2088 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_11527_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2089 a_13441_4949# a_13275_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2090 a_5720_20495# _0845_.A1 a_5417_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2091 vssd1 clkbuf_0__0390_.A a_4802_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2092 vssd1 _1030_.CLK a_18151_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2093 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2095 a_25593_11471# _1013_.Q a_25511_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2096 a_5635_20175# _0812_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2097 a_17971_10089# _0616_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2098 vssd1 _0972_.CLK a_16955_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2099 vssd1 _0959_.CLK a_9411_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2100 vssd1 a_4170_20291# _0764_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2101 vccd1 _0722_.B a_2693_15543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X2102 a_21108_4399# a_20709_4399# a_20982_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2105 a_23224_4399# a_22825_4399# a_23098_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2106 a_17773_15529# _0523_.B1 a_17857_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2107 vccd1 _0935_.CLK a_14747_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2108 a_25589_14735# _0966_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2109 a_23910_6005# a_23742_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2110 a_27847_25437# a_26983_25071# a_27590_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2111 vssd1 a_12375_18811# a_12333_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2112 vccd1 a_2114_1653# _0860_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2113 a_25401_19631# a_25235_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2116 vssd1 a_25842_14709# a_25800_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2117 _0673_.B2 a_4831_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2118 _0438_.A a_2715_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2119 vssd1 a_5325_8181# _0711_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X2120 vssd1 _0845_.C1 _0843_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 a_19770_26677# a_19602_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2122 a_20635_10383# _0563_.B1 a_20717_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2123 _0626_.B1 a_17971_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2124 vccd1 a_6611_25589# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2126 a_27422_12381# a_26983_12015# a_27337_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2127 _0798_.A2 _0722_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 a_20046_15391# a_19878_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2129 vssd1 a_8175_9527# _0689_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2130 a_10957_11293# a_10423_10927# a_10862_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2131 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2132 a_11049_3311# a_10883_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2133 a_13544_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2134 a_17986_13647# _0609_.C1 a_17906_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2135 vccd1 _0439_.A a_5639_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2136 _0849_.X a_12114_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2138 _0673_.A1 a_12927_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2139 vccd1 fanout23.X a_25143_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2140 a_12000_9839# a_11601_9839# a_11874_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2142 _0928_.Q a_28015_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2143 a_17928_8181# _0587_.C1 a_18320_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2144 vccd1 a_4065_14237# a_4165_14455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X2145 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2146 a_16258_18793# _0988_.D a_16101_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2147 a_3283_25615# a_2419_25621# a_3026_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2148 vssd1 _0630_.A2 a_18048_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X2149 vccd1 a_10275_4765# a_10443_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2152 a_27548_15279# a_27149_15279# a_27422_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2153 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2154 vssd1 _1015_.CLK a_23671_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2155 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2156 _0872_.A2 _0803_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2157 vccd1 _1052_.D a_17086_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2158 _0916_.D a_10167_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2159 vccd1 a_15793_6603# _0645_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2160 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15016_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2161 a_27590_5599# a_27422_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2162 a_11251_5737# _0667_.B1 a_11333_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2163 _0572_.A2 a_13735_12925# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X2164 a_11902_26742# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2165 vccd1 fanout37.A a_16495_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2166 vccd1 a_12999_31055# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2168 a_12015_9633# _0479_.Y a_11929_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2171 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_12604_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2172 a_25309_8207# a_24775_8213# a_25214_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2173 vssd1 a_24887_22325# a_24845_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2174 vccd1 a_15151_8029# a_15319_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2175 vccd1 a_26670_20831# a_26597_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2177 vssd1 a_23523_4765# a_23691_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2178 a_7258_5599# a_7090_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2181 _0863_.A2 _0840_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2182 vccd1 a_9983_16885# a_9899_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2183 a_21165_5487# a_20175_5487# a_21039_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2184 a_20153_6409# a_19163_6037# a_20027_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2185 a_8546_1653# a_8378_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2186 a_20635_10383# _0563_.B1 a_20717_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2189 a_17853_10761# a_16863_10389# a_17727_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2190 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2191 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13735_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2192 a_11842_25321# _0825_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2193 vssd1 _0551_.C1 a_17323_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2194 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12631_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2195 a_26670_20831# a_26502_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2197 a_8477_13967# _1080_.Q a_8123_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2198 a_12065_8207# _0916_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2199 a_15496_28169# a_15097_27797# a_15370_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2200 vssd1 a_17010_21919# a_16968_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2201 vssd1 _1076_.Q a_8031_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2203 vccd1 a_5273_29687# _0445_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2204 a_27149_21807# a_26983_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2205 a_23634_17973# a_23466_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2206 vccd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_2686_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2207 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11224_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2208 a_10497_17999# _0749_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2210 a_26183_7119# a_25401_7125# a_26099_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2211 a_13855_22351# a_13073_22357# a_13771_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2212 vccd1 a_18645_7457# _0516_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2215 vccd1 a_23247_19087# a_23415_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2216 a_2455_5853# a_1757_5487# a_2198_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2220 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2221 a_7932_28111# _0821_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2222 a_3777_27081# a_2787_26709# a_3651_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2223 vccd1 a_10551_6031# a_10719_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2224 a_12526_8751# _0840_.A0 a_12437_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X2225 a_27422_25437# a_27149_25071# a_27337_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2226 vccd1 _0440_.A a_6559_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
R7 temp1.capload\[4\].cap_49.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2227 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2228 a_22549_3311# a_22383_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2229 a_18869_25615# a_18335_25621# a_18774_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2230 a_9135_9839# _0475_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2231 a_2464_1653# a_2752_1897# a_2687_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.066 ps=0.745 w=0.36 l=0.15
X2233 vssd1 a_21943_18811# a_21901_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2234 a_5256_15823# _0456_.B a_5001_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2236 a_17861_10927# _0565_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2237 a_21729_7913# _0515_.X a_21647_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2238 a_15105_11791# _0988_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2239 vssd1 fanout27.A a_21003_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2240 a_5141_30199# _0827_.A a_5361_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2242 a_19743_13647# a_18961_13653# a_19659_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2243 a_5161_4943# a_4627_4949# a_5066_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2244 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2245 vccd1 _0443_.A a_11803_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2246 vccd1 _0778_.B1 _0778_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2247 vccd1 _0515_.B1 a_15841_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2248 a_27061_6575# _0562_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2249 a_8803_1679# a_8105_1685# a_8546_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2250 vssd1 _0508_.Y a_12632_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2251 a_21913_10089# _0666_.D a_21831_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2252 vccd1 _0662_.A1 a_14559_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2253 vssd1 _0574_.C a_21065_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2254 a_21173_8751# _0940_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2255 vssd1 _0572_.A2 a_25857_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2256 vssd1 a_13939_22325# a_13897_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2258 vssd1 _0812_.A2 a_6559_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2259 vccd1 a_26267_1403# a_26183_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2260 _0619_.B1 a_22325_6603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X2261 a_13146_1653# a_12978_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2262 a_12299_10205# a_11601_9839# a_12042_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2265 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_7479_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2266 vssd1 a_12777_16885# _0739_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2267 a_27337_16367# _1012_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2268 vccd1 a_2956_1956# a_2885_2057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X2270 a_25857_6575# a_24867_6575# a_25731_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2273 vccd1 a_12299_10205# a_12467_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2274 a_2030_6031# a_1757_6037# a_1945_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2275 vssd1 a_2787_7119# _0888_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2276 a_25750_12127# a_25582_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2277 vccd1 a_12575_13647# a_12743_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2278 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2279 a_6559_19087# _0869_.B1 a_6813_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2280 vssd1 _0444_.B _0825_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2281 vssd1 clkbuf_1_1__f__0390_.A a_2686_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2282 _0583_.A a_20635_13655# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2283 a_14812_31055# a_14563_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2284 a_10689_21853# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2286 vssd1 _0663_.X a_21831_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2287 a_15879_1679# a_15097_1685# a_15795_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2288 a_6817_10703# _0685_.B _0656_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X2289 vssd1 a_26007_12381# a_26175_12283# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2291 vssd1 a_12575_13647# a_12743_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2292 a_17677_6031# _0615_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2293 a_27590_25183# a_27422_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2294 vssd1 a_21150_4511# a_21108_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2296 vssd1 a_23266_4511# a_23224_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2297 a_14747_6031# _0516_.B1 a_14829_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2298 vssd1 _0717_.A2 a_11067_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2300 a_21077_18543# a_20911_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2301 _0840_.X a_4403_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2302 vccd1 a_21023_20149# a_20939_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2303 a_7745_15529# _0812_.A2 a_7663_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2305 vccd1 a_6651_28335# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2306 vssd1 _0845_.C1 a_12547_23145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2307 a_5600_14165# _0734_.C1 a_5992_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2309 a_21258_9117# a_20819_8751# a_21173_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2310 _0531_.X a_20635_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2311 vssd1 a_20027_26703# a_20195_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2312 a_2313_2223# _0858_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2313 a_25309_9839# a_25143_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2314 vssd1 _0837_.A1 a_11764_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2315 a_12532_26159# _0824_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2317 a_11760_26935# _0825_.A1 a_11902_26742# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2318 a_23247_19087# a_22383_19093# a_22990_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2319 vccd1 _0840_.A1 a_9407_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2323 a_13073_22357# a_12907_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2324 a_11040_31055# a_10791_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2325 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2326 a_12604_29967# a_12355_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2327 _1067_.Q a_26267_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 vssd1 _0582_.C a_22169_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2329 a_22291_16617# _0643_.B1 a_22373_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2330 vccd1 a_7111_13655# _0735_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2331 vssd1 a_7775_3829# a_7733_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2333 a_19517_26703# _1018_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2335 vccd1 a_3026_25589# a_2953_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2336 a_17930_6005# a_17762_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2337 vccd1 _0861_.A1 a_16123_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2338 vssd1 a_17909_16395# _0648_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X2339 vssd1 a_6947_2491# a_6905_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2340 vssd1 a_17803_19899# a_17761_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2341 a_27655_6941# a_26873_6575# a_27571_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2342 vssd1 _1062_.CLK a_19991_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2343 a_12079_7119# _0487_.X a_12257_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2345 a_27548_14191# a_27149_14191# a_27422_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2347 vssd1 _0685_.X a_6653_10933# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2348 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2349 _0927_.D a_26083_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2350 vccd1 a_3983_31849# io_out[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2351 vccd1 a_24167_6031# a_24335_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2353 _0574_.C _0471_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2355 _1049_.Q a_21667_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2356 a_18237_18319# _0933_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2358 a_17654_17567# a_17486_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2359 a_9857_21263# _0988_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2362 _0708_.B1 _0807_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2363 vccd1 _0664_.A2 a_22917_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2365 a_10218_2767# a_9779_2773# a_10133_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2366 a_22369_15823# _0925_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2368 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14011_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2369 vssd1 a_8176_19061# _0765_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2371 vssd1 clkbuf_1_0__f_io_in[0].X a_3983_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2372 a_19402_1653# a_19234_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2373 vssd1 a_9742_5599# a_9700_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2374 _0798_.X a_4036_30663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2376 _0940_.Q a_23415_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2377 a_19517_3855# _0969_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2378 vssd1 a_25290_13215# a_25248_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2379 a_15749_12559# _0643_.X a_15667_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2380 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2381 a_27149_21807# a_26983_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2383 _0562_.A1 a_25899_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2384 vssd1 _0722_.C a_4170_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2385 a_12575_13647# a_11711_13653# a_12318_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2386 a_18681_11849# a_17691_11477# a_18555_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2387 _1021_.Q a_22035_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2388 vccd1 a_28015_24251# a_27931_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2391 a_11950_15391# a_11782_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2392 vssd1 _0681_.X _0694_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X2393 a_12995_16911# _0798_.A2 a_12777_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2394 a_23055_2767# a_22273_2773# a_22971_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2395 vssd1 a_10275_4765# a_10443_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2398 vssd1 a_27095_20987# a_27053_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2400 a_24945_21807# _0929_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2401 a_8393_16617# _0717_.A2 _0735_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2402 a_12245_13647# a_11711_13653# a_12150_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2405 _0619_.X a_27167_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2407 vccd1 a_2566_1247# a_2493_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2409 vccd1 _0535_.X a_12805_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2410 vccd1 a_9411_8751# _0917_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2411 a_1757_8751# a_1591_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2412 a_10948_31849# a_10699_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2413 a_2686_28879# clkbuf_1_1__f__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2414 _0577_.X a_17139_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2415 vssd1 _0935_.CLK a_15023_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2416 a_10968_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2417 vssd1 _0778_.B1 a_7164_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2418 a_2683_2767# a_2235_2773# a_2589_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2419 _0654_.Y _0546_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2420 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2421 vssd1 _0533_.X a_17404_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X2422 vccd1 a_14894_7775# a_14821_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2423 _1014_.Q a_28015_12283# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2424 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2425 a_7829_21269# a_7663_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2426 a_19659_1679# a_18961_1685# a_19402_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2427 a_18590_4943# a_18317_4949# a_18505_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2430 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_14812_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2432 a_22980_18543# _0662_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2433 a_21491_3677# a_20709_3311# a_21407_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2436 _0574_.X a_22751_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2438 a_6473_15529# _0758_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2439 vccd1 _0456_.A a_5796_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2441 a_6909_3861# a_6743_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2442 a_4149_26159# a_3983_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2443 vssd1 _0780_.A1 a_5731_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2444 _0902_.Q a_10719_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2445 a_1674_32143# clkbuf_1_1__f_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X2447 a_18072_1135# a_17673_1135# a_17946_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2449 _0460_.C a_1626_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2451 vccd1 fanout23.X a_27521_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2452 a_10551_6031# a_9687_6037# a_10294_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2453 a_4259_7669# _0710_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X2455 _0502_.X a_12763_12879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X2456 vccd1 a_24719_20175# a_24887_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2458 a_25589_16911# _0999_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2460 vccd1 _0825_.X a_6651_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2462 vccd1 _0888_.CLK a_2695_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2463 a_24485_13647# _1046_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2464 a_7001_6941# a_6467_6575# a_6906_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2465 vssd1 _0634_.C1 a_18025_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2466 _0686_.A _0778_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2467 vssd1 a_24719_20175# a_24887_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2468 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11040_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2469 temp1.capload\[2\].cap.Y temp1.capload\[2\].cap_47.LO a_8117_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2470 a_21384_8751# a_20985_8751# a_21258_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2471 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_12604_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2472 a_16768_10927# _0667_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2473 a_14655_4399# _0954_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2474 a_10126_6031# a_9687_6037# a_10041_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2475 a_25800_10761# a_25401_10389# a_25674_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2476 vssd1 a_26635_26427# a_26593_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2477 a_15777_21583# a_15576_21379# _0863_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2478 vssd1 a_7331_6941# a_7499_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2479 vssd1 a_24738_13621# a_24696_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2480 a_16902_6825# _0645_.B2 a_16745_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2484 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2485 a_24017_27081# a_23027_26709# a_23891_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2486 a_12622_24233# _0444_.B a_12316_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2488 a_12069_5263# _0673_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2489 vssd1 a_28015_25339# a_27973_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2490 _0835_.Y _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2491 _0664_.A2 a_21127_11809# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2492 vssd1 _0684_.A2 a_8393_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X2493 _0836_.Y _0836_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2495 a_22199_10499# _0650_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2496 _0556_.D a_12999_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X2497 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2498 a_11873_3311# a_10883_3311# a_11747_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2499 vccd1 a_2198_6005# a_2125_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2500 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15844_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2502 vccd1 _0837_.A1 a_10055_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2503 a_4037_11989# _0745_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2504 vssd1 a_21407_3677# a_21575_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2506 a_11902_27069# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2507 a_15370_1679# a_14931_1685# a_15285_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2509 a_5078_30511# temp1.dcdc.Z vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2510 vccd1 _1081_.Q a_10515_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X2511 vssd1 _0444_.B _0825_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2512 vssd1 _0964_.CLK a_24591_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2513 a_4864_11445# _0807_.B a_5087_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2514 vssd1 a_5417_20149# _0813_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2515 vssd1 _0518_.Y a_16983_12897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2518 vccd1 _0715_.X a_1775_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2519 _1030_.CLK a_16035_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2520 _0523_.B1 a_20393_8545# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X2521 a_6445_3311# a_5455_3311# a_6319_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2522 a_23190_8207# a_22917_8213# a_23105_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2523 a_12150_8207# a_11711_8213# a_12065_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2524 _0535_.X a_12355_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X2525 a_2686_10383# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X2527 a_2490_28701# a_2217_28335# a_2405_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2528 vccd1 _0504_.A a_18519_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2530 a_27149_15279# a_26983_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2531 a_10344_3145# a_9945_2773# a_10218_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2532 a_2655_24501# _0860_.A a_2882_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X2534 a_23745_14735# _0963_.Q a_23661_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2535 vssd1 a_9339_7093# a_9297_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2539 vccd1 a_26083_17723# a_25999_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2540 vssd1 a_12355_8751# _0535_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X2542 vccd1 a_18263_23163# a_18179_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2543 vccd1 _1053_.CLK a_7663_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2544 a_15354_14709# a_15186_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2545 a_2493_1501# a_1959_1135# a_2398_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2546 _0556_.B a_17323_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2547 a_13735_12925# _0472_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2548 a_17083_26525# a_16219_26159# a_16826_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2549 a_2999_25437# a_2217_25071# a_2915_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2551 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2552 a_12815_25071# _0850_.A _0850_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2553 _0471_.X a_9503_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2555 a_4811_27791# _0844_.B _0845_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2556 vccd1 _1028_.CLK a_12355_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2557 vccd1 a_12318_13621# a_12245_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2558 vssd1 a_2823_1501# a_2991_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2560 a_4468_13103# _0745_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2562 _0456_.A _0722_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2563 vccd1 _0935_.CLK a_11343_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2564 a_14821_8029# a_14287_7663# a_14726_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2566 a_19141_5321# a_18151_4949# a_19015_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2568 a_23649_8751# a_22659_8751# a_23523_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2569 vccd1 a_8527_21263# a_8695_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2570 a_27881_8751# a_26891_8751# a_27755_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2572 a_27149_5487# a_26983_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2574 vssd1 _0814_.A2 a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2575 vssd1 a_10147_15529# _0474_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X2576 a_9301_14441# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X2577 vccd1 _0524_.X a_12479_5515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2578 _0798_.A2 _0722_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2579 _1060_.D a_18079_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2580 a_27847_5853# a_26983_5487# a_27590_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2581 a_23174_7093# a_23006_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2583 _1057_.Q a_15503_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2584 _0564_.C a_19531_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2586 a_23005_2057# a_22015_1685# a_22879_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2587 vssd1 a_8527_21263# a_8695_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2588 a_14829_6031# _0671_.B2 a_14747_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2589 a_15134_10383# _0613_.C1 a_15054_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2590 a_15733_11177# _0605_.X a_15661_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2591 vccd1 a_6151_21781# _0809_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2593 a_2689_9839# _0699_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2594 a_4439_9001# _0695_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2595 a_8176_19061# _0763_.B1 a_8305_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2597 a_21767_19997# a_20985_19631# a_21683_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2599 a_17289_13249# _0605_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X2600 vssd1 a_27555_13371# a_27513_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2601 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2604 a_21502_15529# _0582_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2606 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2607 a_8760_28111# _0821_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2608 a_8241_16161# _0807_.A a_8155_16161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2609 a_19617_4399# _0497_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2611 vccd1 _1062_.Q a_17720_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X2613 a_22729_12879# _0938_.Q a_22291_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2614 _0529_.Y a_10814_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2616 a_2114_1653# a_2464_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X2617 a_23469_6037# a_23303_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2618 a_8464_31849# a_8215_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2619 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2621 a_12886_2767# a_12613_2773# a_12801_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2622 vssd1 a_24719_1679# a_24887_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2623 _0630_.A1 a_17895_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2624 a_25382_12533# a_25214_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2626 a_13551_13760# _0936_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2627 a_11238_17705# a_11458_17429# _0574_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2628 a_5797_17027# _0873_.A a_5725_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2631 vssd1 a_23047_1653# a_23005_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2632 vccd1 _0670_.A2 a_15949_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2634 _0863_.A1 a_15575_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2635 vssd1 a_15703_2589# a_15871_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2636 vssd1 a_18114_1247# a_18072_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2638 vccd1 _0835_.A1 a_9687_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2639 a_13012_16201# a_12613_15829# a_12886_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2641 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2642 vccd1 a_25807_23413# a_25723_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2643 _0512_.X a_19195_18337# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2644 a_3241_16617# _0439_.A _0877_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2645 vssd1 _0491_.X a_15001_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2646 _0562_.A1 a_25899_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2647 a_23431_7119# a_22733_7125# a_23174_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2648 vccd1 a_10535_11445# a_10451_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2649 vssd1 a_5323_29111# _0764_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2650 a_18363_3677# a_17581_3311# a_18279_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2651 _0651_.C a_20175_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2652 vssd1 a_4035_25045# _0843_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2655 a_23303_13760# _1012_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2656 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2659 vssd1 _0825_.X a_6651_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2660 a_4403_25589# _0840_.A1 a_4630_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X2661 a_2125_6031# a_1591_6037# a_2030_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2662 a_23373_3311# a_22383_3311# a_23247_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2663 fanout24.A a_16495_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2664 vssd1 a_21426_8863# a_21384_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2665 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2667 a_10252_6409# a_9853_6037# a_10126_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2668 vccd1 _0893_.CLK a_26983_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2669 _0553_.X a_18243_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2671 a_10212_29673# a_9963_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2673 vccd1 io_in[1] a_3983_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2674 vssd1 a_26267_7093# a_26225_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2675 vccd1 _0518_.Y a_13551_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2677 a_26743_23261# a_25879_22895# a_26486_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2681 vssd1 a_21207_5755# a_21165_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2682 vssd1 _0994_.CLK a_24775_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2683 a_5894_3677# a_5621_3311# a_5809_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2684 a_6641_23805# _0847_.A2 a_6559_23552# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2685 vccd1 _0643_.B1 a_23569_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2686 a_5821_13353# _0713_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2689 a_11527_6575# _0522_.B1 a_11705_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2690 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2691 a_22081_10089# _0666_.B a_22009_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2692 vssd1 a_9135_6575# _1028_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2693 a_5078_30511# temp1.dcdc.Z vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2695 _1054_.Q a_15595_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2696 a_15496_2057# a_15097_1685# a_15370_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2697 _0784_.A1 a_11936_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2698 vssd1 a_26083_9019# a_26041_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2699 vccd1 _0527_.X a_23303_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2700 a_15419_17999# a_14637_18005# a_15335_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2701 a_4632_13353# _0776_.A2 a_4035_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X2705 a_25589_19631# _1047_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2706 vccd1 a_14483_15279# a_14603_15325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2707 a_23385_10383# _0621_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2710 a_20993_16189# _0504_.A a_20911_15936# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2711 a_19793_15279# _0962_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2712 a_20761_9633# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2713 vccd1 _0994_.CLK a_23855_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2714 a_8478_9295# _0679_.A2 a_8175_9527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X2715 vccd1 _0778_.A2 a_6559_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X2716 a_13360_26159# _0824_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2717 a_9945_2773# a_9779_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2718 a_12276_8585# a_11877_8213# a_12150_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2719 vssd1 a_13847_9269# a_13805_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2720 a_20083_15936# _0930_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2721 a_17722_14441# _0629_.X a_17473_14337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X2722 vssd1 a_18279_3677# a_18447_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2724 vccd1 _0840_.A0 a_9865_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2726 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2728 a_4973_1135# a_3983_1135# a_4847_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2729 a_9022_3855# a_8583_3861# a_8937_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2731 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2733 vssd1 _0722_.A _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2734 vssd1 _0972_.CLK a_20543_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2736 vccd1 a_25382_23413# a_25309_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2737 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2738 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5724_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2740 a_21909_21807# _1021_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2741 _0994_.CLK a_21279_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2742 a_15036_18377# a_14637_18005# a_14910_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2743 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2744 vssd1 a_4403_22869# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2745 a_22181_1685# a_22015_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2746 a_2907_27613# a_2125_27247# a_2823_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2748 a_3298_17143# _0722_.C a_3435_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2749 io_out[2] _0753_.A2 a_2039_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2751 a_11490_3423# a_11322_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2752 vssd1 a_26835_11293# a_27003_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2753 vccd1 a_5015_28603# a_4931_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2754 a_14342_19061# a_14174_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2755 a_13403_1679# a_12539_1685# a_13146_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2756 a_17761_5487# _0622_.A1 a_17415_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2759 a_6741_14735# _0778_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2761 vccd1 _0784_.A1 a_7291_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2762 vccd1 _0582_.C a_20083_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2763 a_13437_3145# a_12447_2773# a_13311_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2764 vssd1 a_25899_6843# a_25857_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2765 vssd1 _0544_.C a_14011_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X2766 vccd1 _0745_.A1 _0791_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2767 _0945_.D a_17987_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2768 a_9489_5487# _0549_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2769 a_2198_6687# a_2030_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2770 a_17489_2473# _0969_.D a_17405_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2771 a_17657_13621# _0608_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X2773 a_25143_14441# _0648_.A2 a_25225_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2774 a_24386_2767# a_24113_2773# a_24301_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2775 vccd1 _0648_.A2 a_18065_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2776 vssd1 a_3155_21271# _0809_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2777 _0722_.A a_1591_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2779 a_23607_4765# a_22825_4399# a_23523_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2780 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8464_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2781 a_6062_3423# a_5894_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2782 vccd1 input2.X a_3523_6039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2784 a_7006_16911# _0833_.A a_6809_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2785 a_14174_19087# a_13901_19093# a_14089_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2786 a_11877_8213# a_11711_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2787 a_4065_31849# _0814_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2789 vccd1 _1053_.CLK a_12907_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2790 a_8102_21263# a_7829_21269# a_8017_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2791 a_19899_1385# _0516_.B1 a_19981_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2792 vccd1 a_20195_26677# a_20111_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2793 vssd1 _1017_.D a_20548_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2794 vssd1 a_13146_1653# a_13104_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2796 _0798_.A2 _0722_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2797 a_1757_6037# a_1591_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2798 a_15929_4399# _0497_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2799 vccd1 _0466_.A a_9895_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X2800 vccd1 io_in[5] a_1626_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2802 a_15511_23439# a_14729_23445# a_15427_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2803 vssd1 a_28015_2491# a_27973_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2804 a_2132_9295# a_1591_9301# a_2039_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X2805 vssd1 a_9043_12567# _0807_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2807 a_10785_19087# _0860_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2808 a_14536_28585# a_14287_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2809 _0574_.C _0472_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2810 a_22822_3677# a_22549_3311# a_22737_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2811 a_2752_1897# clkbuf_1_0__f_io_in[0].X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2812 a_8887_1679# a_8105_1685# a_8803_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2814 a_25156_16367# a_24757_16367# a_25030_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2816 _0584_.B1 a_22015_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2817 a_8464_30761# a_8215_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2818 _0869_.B1 a_2807_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2819 a_11776_31849# a_11527_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2820 vccd1 _0975_.CLK a_23947_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2821 a_27498_8863# a_27330_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2822 vccd1 fanout37.A a_23763_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2823 a_22438_26271# a_22270_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2824 temp1.capload\[13\].cap.Y temp1.capload\[13\].cap.A a_15017_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2828 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10212_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2829 a_12525_27791# a_12348_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2830 vssd1 _0778_.A2 a_6817_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X2831 vssd1 a_22695_26525# a_22863_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2833 a_25497_9839# _1068_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2834 vccd1 a_26099_3855# a_26267_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2835 _0572_.A1 a_26267_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2836 _0764_.A1 a_4170_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X2837 vccd1 _0614_.A a_15733_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2838 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2839 a_17857_15529# _0937_.Q a_17773_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2840 vssd1 a_16182_14303# a_16140_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2841 vssd1 a_10643_1679# a_10811_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2842 a_16853_9001# _0985_.D a_16771_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2843 a_4406_3829# a_4238_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2844 vssd1 _0999_.CLK a_25235_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2847 a_20598_20149# a_20430_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2850 a_11908_18543# a_11509_18543# a_11782_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2851 a_20717_10383# _0890_.D a_20635_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2852 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2853 vccd1 a_10735_2589# a_10903_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2854 vssd1 a_8270_21237# a_8228_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2856 a_14093_21263# _0863_.A1 _0864_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2857 a_13514_10357# a_13346_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2858 vccd1 _0735_.A2 a_11233_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2859 vccd1 a_18611_14191# _0931_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2860 a_13367_6575# _0604_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2862 vssd1 a_23082_20831# a_23040_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2863 a_14916_6825# _0565_.B1 a_14661_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2864 a_18409_9001# _0987_.D a_18325_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2865 a_17302_10383# a_16863_10389# a_17217_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2867 vssd1 a_27847_24349# a_28015_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2868 a_9577_4399# a_9411_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2869 a_7032_7663# _0657_.X _0694_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
X2870 a_10325_15055# _0770_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2871 a_20430_20175# a_20157_20181# a_20345_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2872 a_15848_7235# _0642_.C a_15753_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X2873 a_14599_19087# a_13901_19093# a_14342_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2874 a_23373_14191# a_22383_14191# a_23247_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2876 a_12610_21263# a_12337_21269# a_12525_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2877 a_14174_19087# a_13735_19093# a_14089_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2878 a_15354_14709# a_15186_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2879 vccd1 clkbuf_1_0__f_io_in[0].X a_1959_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2880 a_22273_2773# a_22107_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2881 a_13346_10383# a_13073_10389# a_13261_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2883 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_12999_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2884 a_27057_8751# a_26891_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2886 a_10160_14025# a_9761_13653# a_10034_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2887 a_12978_1679# a_12539_1685# a_12893_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2889 vssd1 a_2198_6005# a_2156_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2890 vssd1 _0565_.B1 a_17928_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2891 a_12150_11471# a_11711_11477# a_12065_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2892 a_19233_21641# a_18243_21269# a_19107_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2893 a_22990_3423# a_22822_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2894 vccd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_2686_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2895 a_4864_15797# _0807_.B a_5084_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2896 a_26133_6409# a_25143_6037# a_26007_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2898 a_9148_4233# a_8749_3861# a_9022_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2899 a_4802_27247# clkbuf_0__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2900 vccd1 _0893_.CLK a_22383_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2901 a_15186_14735# a_14913_14741# a_15101_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2903 a_10252_22729# a_9853_22357# a_10126_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2904 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2905 a_7642_4765# a_7203_4399# a_7557_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2906 vssd1 _0935_.CLK a_12171_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2907 a_27931_3677# a_27149_3311# a_27847_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2909 a_6736_30287# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2910 a_24462_22325# a_24294_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2911 a_11893_20175# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2912 vccd1 _0861_.X a_3326_2057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0672 ps=0.74 w=0.42 l=0.15
X2914 vccd1 _0702_.B1_N a_5210_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2915 a_21077_3677# a_20543_3311# a_20982_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2916 vccd1 _0722_.C a_5001_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2918 _0794_.A3 _0466_.A a_5909_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2919 _0860_.B a_11067_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X2920 a_25497_6031# _0506_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2921 vccd1 _1075_.Q a_14471_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2922 a_9949_13647# _0921_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2926 a_23006_7119# a_22733_7125# a_22921_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2928 a_24294_22351# a_24021_22357# a_24209_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2929 a_17930_6005# a_17762_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2930 vccd1 a_25915_8029# a_26083_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2931 _0612_.X a_19439_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2932 a_23936_13103# _0572_.A1 a_23361_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X2933 a_20671_14735# a_19973_14741# a_20414_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2934 a_15017_31599# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2936 a_6832_8527# _0689_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2939 a_27517_2589# a_26983_2223# a_27422_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2940 a_17865_12925# _0602_.A a_17783_12672# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2941 a_25198_21919# a_25030_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2942 vssd1 a_7623_10901# _0776_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2943 a_19659_13647# a_18795_13653# a_19402_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2944 a_24757_5487# a_24591_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2946 a_11697_20719# _0987_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2947 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2948 vccd1 _0590_.X a_18677_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2949 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_14536_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2950 vssd1 a_15667_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2953 _0963_.D a_20471_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2954 a_4590_1247# a_4422_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2955 a_7350_3829# a_7182_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2956 a_3643_4943# a_2861_4949# a_3559_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2957 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8464_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2958 a_13311_15823# a_12447_15829# a_13054_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2959 vccd1 a_21610_13215# a_21537_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2960 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11776_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2962 a_8749_3861# a_8583_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2964 a_20855_20175# a_20157_20181# a_20598_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2965 a_23070_18543# _1048_.D a_22980_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X2966 a_21357_23983# _1020_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2967 a_8301_27247# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2968 a_21081_27247# _1019_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2972 a_7479_29673# _0827_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2973 a_24278_11445# a_24110_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2974 a_5428_29429# _0445_.B a_5356_29429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X2975 a_13346_10383# a_12907_10389# a_13261_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2976 a_1945_6575# _0877_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2979 vccd1 a_25842_14709# a_25769_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2981 _1011_.D a_26267_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2982 a_23837_6031# a_23303_6037# a_23742_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2983 vssd1 _0847_.A3 a_11969_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X2984 _1012_.D a_25715_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2985 a_25589_25615# _0993_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2986 a_21859_18909# a_21077_18543# a_21775_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2987 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2988 a_6612_14709# _0793_.X a_6741_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2989 a_8033_10703# _0678_.Y _0746_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2990 a_2030_5853# a_1591_5487# a_1945_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2991 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2992 vssd1 a_24462_22325# a_24420_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2993 vccd1 a_7515_5853# a_7683_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2994 vccd1 _0847_.A2 a_11893_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2996 vccd1 a_17010_21919# a_16937_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
R8 vccd1 temp1.capload\[14\].cap_44.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2997 vccd1 a_3891_21263# _0814_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2998 vssd1 a_11950_20831# a_11908_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3001 a_12333_2223# _0945_.D a_11987_2473# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3002 vccd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_1674_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3005 vccd1 _0866_.B a_12725_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3006 vssd1 _0685_.B _0680_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3007 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_6651_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3008 a_12547_23145# a_12355_22901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X3009 a_14726_12381# a_14453_12015# a_14641_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3010 a_5549_17719# _0456_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3011 _0922_.CLK a_4259_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3012 vssd1 a_6487_3579# a_6445_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3013 _0829_.A1 a_5015_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3014 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3015 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3016 vssd1 a_22971_2767# a_23139_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3017 a_6559_15823# _0736_.B1 a_6737_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3018 a_4847_28701# a_4149_28335# a_4590_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3019 a_27149_15279# a_26983_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3020 vssd1 _0643_.B1 a_27513_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3022 a_8378_1679# a_7939_1685# a_8293_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3025 a_3240_14441# _0456_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X3026 a_21173_8751# _0940_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3027 a_7350_3829# a_7182_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3028 a_18600_7663# _1031_.Q a_18025_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X3030 a_11895_1385# _0850_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3031 vssd1 a_8123_20719# _0827_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3033 vssd1 a_26099_19087# a_26267_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3034 _0735_.A2 a_7111_13655# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3035 vccd1 a_12189_27001# a_12219_26742# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3037 vssd1 _0798_.X a_5361_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3039 a_15377_16367# _0990_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3040 vssd1 _0935_.CLK a_11343_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3041 _0869_.B1 a_2807_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3042 a_14453_7663# a_14287_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3043 a_23837_11477# a_23671_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3044 a_13901_19093# a_13735_19093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3046 vssd1 a_23691_9019# a_23649_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3047 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8944_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3048 a_20911_1385# _0645_.B1 a_20993_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3049 io_out[7] a_3983_31849# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3051 _0964_.CLK a_23855_15831# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3054 vccd1 a_21499_21085# a_21667_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3056 a_4530_9295# _0699_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3057 vccd1 _0625_.A1 a_10410_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X3058 _0599_.X a_14287_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3060 vccd1 _0717_.A2 a_6725_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X3062 a_11877_11477# a_11711_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3065 a_23776_21641# a_23377_21269# a_23650_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3066 vssd1 a_20471_17723# a_20429_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3067 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3068 a_7768_4399# a_7369_4399# a_7642_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3069 _1066_.D a_28015_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3070 a_7415_6941# a_6633_6575# a_7331_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3072 a_12150_6031# a_11877_6037# a_12065_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3073 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3074 a_20414_7775# a_20246_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3075 vccd1 _1024_.Q a_19846_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3077 vccd1 _0975_.CLK a_22383_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3080 vssd1 a_23247_14557# a_23415_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3081 vssd1 fanout27.A a_20819_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3082 temp1.capload\[8\].cap.Y temp1.capload\[8\].cap.A a_12441_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3083 _0854_.X a_25707_25321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X3084 vccd1 a_13571_1653# a_13487_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3086 a_21610_13215# a_21442_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3087 a_11793_2045# _0842_.A0 a_11711_1792# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3088 a_20414_7775# a_20246_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3089 a_12069_2473# _0902_.Q a_11987_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3090 a_20911_15936# _0995_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3091 a_8393_16617# _0735_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X3092 vssd1 _0529_.Y a_20385_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3093 vssd1 a_15023_28887# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3095 _0715_.X a_2693_15543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X3096 a_25198_15391# a_25030_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3097 a_20614_5853# a_20341_5487# a_20529_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3098 a_18455_1501# a_17673_1135# a_18371_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3099 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3100 a_12981_2767# a_12447_2773# a_12886_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3101 _0807_.C a_5639_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3102 vccd1 a_24554_2741# a_24481_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3104 a_9613_25045# _0816_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3105 _0472_.X a_8859_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3106 vssd1 a_9447_3855# a_9615_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3107 a_24315_10496# _0573_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3108 a_2686_28879# clkbuf_1_1__f__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3110 vssd1 a_27279_18811# a_27237_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3111 vssd1 a_10055_23983# _0847_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3112 a_22377_12015# _0892_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3114 a_25490_17821# a_25217_17455# a_25405_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3115 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3116 vssd1 _0908_.CLK a_4167_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3119 a_17670_23261# a_17397_22895# a_17585_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3121 vccd1 _0512_.X a_18225_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X3122 a_13882_4917# a_13714_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3123 vccd1 _0583_.A a_15943_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3124 vssd1 _0814_.A2 a_6559_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3125 a_18942_25589# a_18774_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3126 vccd1 _0861_.B1 a_12356_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3127 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3128 _0579_.X a_17231_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3129 a_12242_27791# a_12065_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3131 a_23303_16617# _0648_.B1 a_23385_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3132 vssd1 a_22990_1247# a_22948_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3133 vccd1 a_13054_15797# a_12981_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3134 a_6498_10089# _0778_.A2 a_6416_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3135 a_17946_11293# a_17507_10927# a_17861_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3138 vccd1 _0574_.C a_20911_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3139 vccd1 a_22990_3423# a_22917_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3140 vssd1 _0893_.CLK a_26983_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3142 a_7256_17429# _0812_.A2 a_7648_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3143 ANTENNA_7.DIODE a_3983_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3144 vccd1 temp1.capload\[4\].cap.A temp1.capload\[4\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3146 vccd1 _0848_.X a_12114_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X3147 vccd1 a_20471_15547# a_20387_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3148 _0589_.X a_19439_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X3149 a_14641_12015# _0897_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3150 a_24945_16367# _0938_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3153 _0531_.A1 a_27463_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3154 a_8485_12879# _0546_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3155 vccd1 a_8123_20719# _0827_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3156 a_6725_15823# _0440_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3157 vssd1 a_25623_2491# a_25581_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3159 vssd1 _0644_.A2 a_16105_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X3161 vssd1 a_25842_19061# a_25800_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3162 vccd1 a_18187_6031# a_18355_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3163 a_10218_4943# a_9945_4949# a_10133_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3164 a_2156_5487# a_1757_5487# a_2030_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3165 a_2455_6941# a_1591_6575# a_2198_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3166 a_27422_16733# a_26983_16367# a_27337_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3167 _0649_.B2 a_20563_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3168 _0721_.A a_2975_17461# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X3169 a_6354_2589# a_6081_2223# a_6269_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3171 a_19471_6603# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3172 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_4988_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3174 vssd1 a_25915_8029# a_26083_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3176 a_15005_5737# _0543_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3178 a_6559_27023# _0444_.B _0752_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3180 a_3134_4943# a_2695_4949# a_3049_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3181 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3182 a_8117_27023# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3183 vssd1 _0798_.A2 a_11044_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3184 vccd1 a_7607_3855# a_7775_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3185 _0861_.B1 a_3799_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3186 vccd1 a_4037_11989# _0791_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3187 _0863_.Y a_15576_21379# a_15777_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3188 vccd1 a_6423_8903# _0698_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X3189 vccd1 a_19770_26677# a_19697_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3190 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3191 a_13882_4917# a_13714_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3192 a_8504_2057# a_8105_1685# a_8378_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3193 _0634_.C1 a_19991_5056# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3195 a_18378_18543# _1053_.D a_18288_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3196 a_4621_16367# _0807_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3197 a_21445_2223# a_21279_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3199 a_23742_9295# a_23469_9301# a_23657_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3200 a_4356_23983# _0752_.Y io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3202 a_25674_3855# a_25235_3861# a_25589_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3204 vccd1 a_23487_15279# _0893_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3205 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3206 vssd1 _0739_.B1 a_7348_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3207 a_15737_3311# a_14747_3311# a_15611_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3208 vssd1 _0917_.CLK a_14287_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3209 vccd1 a_19183_20149# a_19099_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3210 vssd1 _1028_.CLK a_12539_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3213 a_27471_13469# a_26689_13103# a_27387_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3214 vssd1 a_26743_23261# a_26911_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3215 a_27149_14191# a_26983_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3216 vssd1 a_17727_2767# a_17895_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3218 a_8929_5321# a_7939_4949# a_8803_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3219 a_4993_11791# _0708_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3220 a_12557_19407# a_12356_19203# _0865_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3221 a_27548_25071# a_27149_25071# a_27422_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3223 a_4101_5515# _0695_.A1 a_4015_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3224 a_7389_25335# _0845_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3228 a_27847_10205# a_27149_9839# a_27590_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3229 vssd1 a_24703_11445# a_24661_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3230 a_20157_20181# a_19991_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3231 vccd1 a_22622_15797# a_22549_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3232 a_15005_5737# _0543_.B2 a_14921_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3234 a_8293_4943# _0538_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3236 a_15879_6603# _0504_.A a_15793_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3237 _0845_.Y _0845_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3238 vssd1 a_7810_4511# a_7768_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3239 vssd1 a_7515_5853# a_7683_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3240 vccd1 a_16101_18517# _0667_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3241 a_24481_2767# a_23947_2773# a_24386_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3243 a_8478_12265# _0684_.A2 a_8175_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X3245 vssd1 a_2991_27515# _1076_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3246 vssd1 a_13551_8215# _0582_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3248 a_17029_3861# a_16863_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3249 vccd1 a_2915_28701# a_3083_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3250 vssd1 a_13679_9295# a_13847_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R9 vccd1 temp1.capload\[0\].cap_39.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3254 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_14287_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3255 vccd1 _0819_.S temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3256 _1040_.Q a_19183_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3257 _0522_.B1 a_16897_16395# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X3258 a_24867_17999# _0662_.B1 a_24949_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3259 _0927_.D a_26083_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3260 a_9117_16917# a_8951_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3261 _0842_.A0 a_11435_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3262 a_21258_9117# a_20985_8751# a_21173_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3263 vssd1 a_4040_10901# _0745_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3264 a_25490_9117# a_25217_8751# a_25405_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3265 _0836_.Y _0845_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3266 _0933_.Q a_18263_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3267 a_25198_4511# a_25030_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3268 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3269 a_15630_16479# a_15462_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3271 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3273 a_15235_10205# a_14453_9839# a_15151_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3274 a_10998_19407# _0813_.A2 a_10703_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X3275 vccd1 a_17911_17821# a_18079_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3277 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A a_8760_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3278 a_1591_22057# _0752_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3279 vssd1 a_5234_4917# a_5192_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3280 a_7564_30287# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3281 vssd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_2686_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3282 a_22419_22173# a_21721_21807# a_22162_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3283 vssd1 a_7073_20149# _0789_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3284 a_19439_12675# _0576_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3289 vssd1 a_22035_13371# a_21993_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3290 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3291 a_2593_15325# _0460_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3293 a_25765_8585# a_24775_8213# a_25639_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3294 a_14542_20175# a_14103_20181# a_14457_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3295 _0660_.X a_25695_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3297 _0461_.A a_3983_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3298 vccd1 a_27590_12127# a_27517_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3299 vccd1 _0847_.A3 a_9687_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X3300 a_4663_3855# a_3799_3861# a_4406_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3301 a_2547_3855# a_1683_3861# a_2290_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3302 vssd1 clkbuf_1_0__f_io_in[0].X a_1591_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3304 a_2864_24893# a_2833_24759# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X3305 _0797_.B1 a_6876_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3307 vccd1 a_28015_17723# a_27931_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3308 _0574_.C a_11458_17429# a_11238_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3309 a_5635_20175# _0812_.B1 a_5417_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3310 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3311 a_5639_29967# _0798_.X a_5141_30199# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3312 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3313 vssd1 a_3028_14165# _0758_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3314 vssd1 _0472_.X a_12447_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X3317 vccd1 a_14524_6549# _0544_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3318 a_10788_25615# a_10515_25615# _0847_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3319 a_17581_3311# a_17415_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3321 vssd1 a_2198_5599# a_2156_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3324 a_21200_20719# a_20801_20719# a_21074_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3325 a_17139_18543# _1054_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3326 a_4337_2223# _0865_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3329 vssd1 a_4406_3829# a_4364_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3330 vssd1 a_2290_3829# a_2248_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3331 _0833_.A a_7939_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3332 _0596_.A1 a_5659_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3334 vccd1 fanout27.A a_17691_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3335 a_25800_21641# a_25401_21269# a_25674_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3336 vccd1 a_14139_4943# a_14307_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3337 a_3260_5321# a_2861_4949# a_3134_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3338 vssd1 _0778_.A2 a_7357_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3339 a_16029_20175# _0860_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X3341 _1031_.Q a_23783_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3342 a_27755_9117# a_26891_8751# a_27498_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3344 vssd1 _0439_.A a_5547_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3345 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3346 _0620_.X a_25143_14441# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3347 a_9393_7663# a_9227_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3348 a_6750_28918# _0825_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3349 vccd1 a_18555_11471# a_18723_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3350 _0726_.X a_6559_23552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3351 _0644_.A2 a_15975_10721# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3353 vssd1 _0472_.X _0838_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3355 a_25581_5487# a_24591_5487# a_25455_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3356 vccd1 _0829_.A1 a_14093_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3357 a_25800_4233# a_25401_3861# a_25674_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3358 a_13081_2473# _0535_.X a_13165_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3361 vssd1 _0836_.A a_11458_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3362 vssd1 a_18555_11471# a_18723_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3363 a_24803_20175# a_24021_20181# a_24719_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3364 a_12318_11445# a_12150_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3365 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3366 vssd1 _0584_.A2 a_18129_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X3367 vssd1 a_10719_6005# a_10677_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3368 a_9217_10089# _0653_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3369 a_15916_29673# a_15667_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3370 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13360_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3371 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3372 vssd1 a_12042_9951# a_12000_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3374 _0558_.X a_24867_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3375 vssd1 a_27111_18909# a_27279_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3376 a_10147_14735# _0770_.B1 a_10325_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3377 a_6612_8181# _0686_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3378 a_26099_4943# a_25235_4949# a_25842_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3380 a_10413_17999# _0749_.B1 a_10497_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3381 a_15115_9295# _0644_.X a_15369_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3382 _0531_.A1 a_27463_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3383 a_9284_10901# a_9495_11249# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X3384 a_16945_15101# _0521_.A a_16863_14848# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3385 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3386 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3387 a_26578_11039# a_26410_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3388 vssd1 fanout11.A a_11619_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3389 vccd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3390 vccd1 a_10689_21853# a_10789_22071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X3392 a_12150_11471# a_11877_11477# a_12065_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3393 vssd1 a_21023_20149# a_20981_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3394 _0901_.Q a_10259_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3395 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3396 a_17489_6037# a_17323_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 vssd1 _0574_.X a_23637_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3398 a_11582_13077# a_11435_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X3400 vccd1 fanout24.A a_27202_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X3402 _0918_.D a_12743_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3403 a_23006_7119# a_22567_7125# a_22921_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3404 a_2589_2767# _0852_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X3405 a_4705_2767# _0586_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3406 _0647_.X a_27167_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3408 _0918_.D a_12743_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3409 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3410 a_18059_4399# _1001_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3411 vccd1 a_10018_4511# a_9945_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3414 vssd1 _0662_.A3 a_22537_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3415 a_20267_6825# _0630_.A2 a_20349_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3416 a_6365_20719# _0845_.A1 a_6283_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3417 _0722_.C a_1867_15831# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3419 a_20429_15279# a_19439_15279# a_20303_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3420 vccd1 a_20782_5599# a_20709_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3421 vssd1 a_16745_6549# _0646_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3422 vssd1 a_13771_10383# a_13939_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3423 vssd1 a_6467_16367# _0717_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3424 a_3041_28335# a_2051_28335# a_2915_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3425 _0713_.A3 a_6600_11587# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3427 a_3167_24527# _0838_.A0 a_2655_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X3428 a_25769_3855# a_25235_3861# a_25674_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3429 a_17562_1653# a_17394_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3430 a_4035_25045# _0842_.A0 a_4244_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X3433 _1034_.Q a_26175_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3434 a_20709_4399# a_20543_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3435 a_22825_4399# a_22659_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3436 a_25857_11791# _0650_.A1 a_25511_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3437 a_17937_12925# _1026_.Q a_17865_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3439 a_11950_20831# a_11782_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3440 a_3435_17231# _0807_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3442 a_6809_16911# _0833_.A a_7006_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3443 a_7472_25077# _0850_.A a_7389_25335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3444 _0833_.A a_7939_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3445 vccd1 _0664_.A2 a_20717_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3446 vssd1 a_12318_11445# a_12276_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3447 vssd1 _0847_.A2 a_12355_22901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X3448 vssd1 _0636_.X a_12079_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 a_18114_11039# a_17946_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3451 vssd1 _0524_.X a_21213_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3452 a_25842_16885# a_25674_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3453 a_15703_2589# a_14839_2223# a_15446_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3454 a_12797_7913# _0646_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3455 a_18555_11471# a_17691_11477# a_18298_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3456 io_out[3] a_1585_24135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3457 a_26099_16911# a_25401_16917# a_25842_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3459 a_25382_23413# a_25214_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3461 vssd1 a_16055_16635# a_16013_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3462 a_26099_3855# a_25401_3861# a_25842_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3463 a_9853_6037# a_9687_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3464 io_out[4] _0774_.A2 a_4439_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3465 a_23886_12559# _0576_.D1 a_23637_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3467 a_15427_23439# a_14563_23445# a_15170_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3469 a_24945_4399# _0548_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3470 a_5821_13353# _0713_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3471 vssd1 _0768_.A1 a_4772_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3472 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3473 a_6611_25589# _0809_.B2 a_6893_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X3475 vccd1 _1019_.CLK a_17231_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3476 vssd1 _0735_.A2 a_5600_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X3477 vssd1 _1075_.Q a_12047_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X3478 a_21134_11177# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X3479 vssd1 _0845_.A2 a_4441_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3480 vssd1 _0545_.A1 a_10084_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3481 a_6646_10703# _0778_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X3482 vccd1 a_10386_4917# a_10313_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3483 vccd1 a_2623_6843# a_2539_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3485 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3488 _0643_.B1 a_20025_10955# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
R10 temp1.capload\[12\].cap_42.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3490 a_27590_24095# a_27422_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3491 a_22181_20181# a_22015_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3492 vccd1 a_6522_2335# a_6449_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3493 _0829_.A1 a_5015_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3494 a_15097_23439# a_14563_23445# a_15002_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3495 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3496 a_8763_14735# _0546_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3497 vssd1 a_13311_15823# a_13479_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3498 a_2455_6031# a_1757_6037# a_2198_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3499 _0681_.X a_7203_9408# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3500 a_6608_29111# _0825_.A0 a_6750_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3501 vssd1 a_26099_10383# a_26267_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3503 _0847_.A1 clkbuf_1_0__f_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3504 vssd1 a_24167_6031# a_24335_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3505 a_26919_11293# a_26137_10927# a_26835_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3506 a_10313_14735# _0807_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3507 vccd1 a_6795_14343# _0779_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X3508 a_12797_7913# _0924_.D a_12713_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3509 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15916_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3511 vssd1 clkbuf_1_0__f_io_in[0].X a_1959_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3512 _0746_.A2 _0678_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X3513 _0638_.X a_18059_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3514 vccd1 a_23910_9269# a_23837_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3515 vccd1 a_22990_14303# a_22917_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3516 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3518 _0931_.CLK a_18611_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3519 a_4915_25615# _0840_.A0 a_4403_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X3521 vccd1 a_23247_3677# a_23415_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3522 a_4517_2773# a_4351_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3523 vccd1 a_25842_19743# a_25769_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3524 vccd1 a_12318_8181# a_12245_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3525 vccd1 _0494_.X a_20025_10955# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3526 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3527 vccd1 _0483_.X a_19991_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3528 a_10129_13647# a_9595_13653# a_10034_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3529 vssd1 _0975_.CLK a_22383_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3530 a_25581_21807# a_24591_21807# a_25455_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3531 a_24719_22351# a_24021_22357# a_24462_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3533 a_2962_14735# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3534 a_15649_20719# a_15483_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3535 a_15949_6031# _0670_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3536 _0946_.Q a_15779_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3537 a_23358_8181# a_23190_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3538 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3539 a_4802_27247# clkbuf_0__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3540 a_10948_32143# a_10699_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3542 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3543 a_11877_6037# a_11711_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3544 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3545 a_25769_26159# a_25603_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3546 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12539_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3547 vssd1 a_25623_16635# a_25581_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3548 a_23132_7497# a_22733_7125# a_23006_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3549 a_27517_22173# a_26983_21807# a_27422_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3550 a_11893_20175# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3551 a_1735_29941# _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X3553 a_27847_17821# a_27149_17455# a_27590_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3554 a_22097_14013# _0521_.A a_22015_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3556 a_5541_29199# _0764_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3560 vccd1 a_4864_15797# _0795_.A1_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3562 a_23569_6575# _0552_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3565 a_18225_17999# _0933_.Q a_18141_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3567 vssd1 _0972_.CLK a_19163_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3570 vssd1 _0546_.A2 a_8477_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X3572 a_25198_5599# a_25030_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3573 _0988_.D a_12375_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3574 vccd1 a_21426_8863# a_21353_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3575 vccd1 _0812_.A2 a_10497_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X3576 vccd1 a_6516_18695# _0797_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X3577 a_12342_1385# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3578 a_7557_4399# _0907_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3579 a_4132_17429# a_3983_17455# a_4582_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X3580 a_5909_11791# _0768_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3581 vssd1 a_2122_12015# a_2228_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3583 vssd1 io_in[0] a_2962_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3584 a_22454_1679# a_22181_1685# a_22369_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3586 a_6633_6575# a_6467_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3587 a_19773_18689# _0584_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X3588 vssd1 _0529_.Y a_18087_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3589 vssd1 _0471_.X a_11435_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3590 a_22199_12015# _0563_.B1 a_22377_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3592 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3593 a_20671_8029# a_19807_7663# a_20414_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3594 a_16757_21807# _0933_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3595 a_10313_4943# a_9779_4949# a_10218_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3596 vccd1 _1028_.CLK a_9135_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3597 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3600 _0444_.B a_11803_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3601 vssd1 a_7900_14165# _0770_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X3603 a_13346_22351# a_12907_22357# a_13261_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3604 a_22733_7125# a_22567_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3605 vssd1 _0475_.X a_10335_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X3606 _0771_.C1 a_10147_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X3607 vccd1 a_2715_3829# a_2631_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3608 _0901_.Q a_10259_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3609 vccd1 a_4831_3829# a_4747_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3610 _1072_.D a_26267_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3611 vssd1 a_10811_4917# a_10769_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3614 _0847_.A3 a_10055_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3615 a_17635_19997# a_16771_19631# a_17378_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3616 a_15186_14735# a_14747_14741# a_15101_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3617 vssd1 a_2623_9019# a_2581_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3620 vssd1 _0860_.B a_15729_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3621 a_25401_16917# a_25235_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3622 _0587_.C1 a_12723_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3623 a_2566_1247# a_2398_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3625 a_14453_14557# a_14287_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X3626 vccd1 a_25750_9951# a_25677_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3627 a_8033_10703# _0679_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X3628 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3629 vccd1 _0964_.CLK a_26983_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3630 a_11697_15279# _0988_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3632 a_6958_21379# _0813_.A2 a_6876_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3633 a_4537_10927# _0698_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3634 a_9791_12015# _0833_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X3636 a_25455_4765# a_24591_4399# a_25198_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3637 vssd1 a_12318_6005# a_12276_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3638 a_25290_13215# a_25122_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3639 a_16123_25615# _0861_.B1 a_15905_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3640 a_10202_18517# a_10055_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X3641 a_6682_26409# _0819_.S a_6600_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3642 a_2953_25615# a_2419_25621# a_2858_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3643 a_25842_19743# a_25674_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3644 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3645 a_15777_21583# _0863_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3648 vccd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_1674_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3649 vssd1 a_15779_3579# a_15737_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3650 a_13395_2767# a_12613_2773# a_13311_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3651 _0444_.B a_11803_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3652 vssd1 a_23047_20149# a_23005_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3653 a_6336_15253# _0735_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3655 a_8338_20291# _0761_.B a_8256_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3656 a_12245_8207# a_11711_8213# a_12150_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3659 _0577_.C a_10202_18517# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3660 a_27697_6575# a_26707_6575# a_27571_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3661 _0753_.A2 a_9687_19881# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3662 a_8105_18793# _0833_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3663 vccd1 _0698_.B1 a_5727_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3665 vssd1 _0674_.C1 a_11527_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3667 vccd1 a_27923_9019# a_27839_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3668 a_25340_12937# a_24941_12565# a_25214_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3669 a_11509_18543# a_11343_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3670 a_11245_14191# _0747_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3672 a_23891_17999# a_23193_18005# a_23634_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3673 _0600_.X a_15943_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3674 vssd1 a_11685_25045# fanout11.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3675 a_25225_9295# _0506_.A2 a_25309_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3677 vccd1 a_14767_19061# a_14683_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3678 vccd1 a_3099_2767# a_3270_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X3679 vssd1 a_27847_2589# a_28015_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3680 vccd1 _0461_.A a_6467_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3681 vssd1 _0835_.A1 _0749_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3682 vccd1 a_8695_21237# a_8611_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3683 a_19517_6031# _0941_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3685 a_4153_3855# _0908_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3686 a_2037_3855# _0882_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3687 a_20985_8751# a_20819_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3688 _0837_.Y _0836_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3689 vccd1 a_22695_26525# a_22863_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3690 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3692 vccd1 a_26267_4917# a_26183_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3694 vccd1 a_14805_10357# _0614_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X3695 a_21357_23983# _1020_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3697 a_13714_4943# a_13275_4949# a_13629_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3698 a_23098_9117# a_22659_8751# a_23013_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3700 _0837_.A1 a_2991_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3701 a_24937_10927# _0562_.A1 a_24591_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3702 vssd1 _0444_.A a_2051_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3703 _0831_.D a_9811_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3704 a_15945_21263# _0863_.A2 _0863_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3705 a_18758_20149# a_18590_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3706 vssd1 _0491_.X a_12517_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X3707 _0611_.B a_5199_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3708 a_6403_3677# a_5621_3311# a_6319_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3709 a_21353_9117# a_20819_8751# a_21258_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3710 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3711 a_17210_19997# a_16937_19631# a_17125_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3712 vssd1 _0935_.CLK a_13735_19093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3714 a_15649_20719# a_15483_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3716 a_18213_4399# _1001_.Q a_18141_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3717 io_out[4] _0752_.Y a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3718 _0521_.A a_13459_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3719 vssd1 _0823_.A a_11746_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3720 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3721 _0588_.X a_15023_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3722 a_4931_26525# a_4149_26159# a_4847_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3723 _1052_.D a_17803_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3724 vssd1 clkbuf_1_0__f_io_in[0].X a_1591_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3725 vssd1 a_5692_13077# _0714_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3726 _0791_.A2 a_5091_12021# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X3729 vssd1 _0602_.A a_20635_13655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3730 a_18590_20175# a_18317_20181# a_18505_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3732 a_8464_32143# a_8215_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3733 a_2686_31055# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3734 vssd1 clkbuf_1_0__f_io_in[0].X a_1683_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3735 a_4852_5737# _0694_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3736 a_19693_8527# _1016_.D a_19347_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3737 vssd1 _0908_.CLK a_3799_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3738 a_12565_5515# _0842_.A0 a_12479_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3740 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3741 a_12337_21269# a_12171_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3742 vssd1 a_2658_25183# a_2616_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3743 vssd1 a_25455_22173# a_25623_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3744 vccd1 _0845_.A1 a_6283_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3745 a_25497_3311# _0505_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3746 vccd1 _0888_.CLK a_7939_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3747 vccd1 a_26007_6031# a_26175_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3748 a_17857_6031# a_17323_6037# a_17762_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3750 a_23565_21263# _1048_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3751 a_26325_10927# _1063_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3752 vssd1 a_10055_23983# _0847_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3754 a_3028_14165# a_2879_14191# a_3324_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3755 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3756 a_22085_7663# _1003_.Q a_21647_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3757 a_9687_23439# _0444_.B _0816_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X3758 vccd1 _0827_.A a_11977_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3760 vccd1 a_11950_20831# a_11877_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3762 a_8067_4765# a_7203_4399# a_7810_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3763 a_22015_5737# _0645_.B1 a_22097_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3764 a_18243_8751# _0667_.B1 a_18421_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3765 a_7203_10089# _0655_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3766 vccd1 _0602_.A a_24315_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3767 a_4036_30663# _0814_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X3768 a_2539_5853# a_1757_5487# a_2455_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3769 a_25639_8207# a_24775_8213# a_25382_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3770 a_25589_19087# _1067_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3771 vccd1 a_13939_10357# a_13855_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3772 a_7896_11703# _0836_.A a_8038_11510# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3773 vssd1 _0557_.X a_16829_12161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3774 vccd1 a_27698_4943# a_27804_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X3775 vssd1 _0917_.CLK a_11435_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3776 a_18065_8207# _0965_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3777 vccd1 a_21610_24095# a_21537_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3779 vssd1 a_5599_6263# _0694_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3780 vccd1 a_15871_2491# a_15787_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3781 a_18501_25621# a_18335_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3782 vssd1 a_6319_3677# a_6487_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3784 _0967_.Q a_26267_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3785 a_23009_21085# a_22475_20719# a_22914_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3788 vccd1 a_15779_14709# a_15695_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3789 a_22015_18112# _0928_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3790 a_14644_16143# _0471_.X a_14341_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3792 vccd1 _0533_.X a_17029_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X3794 a_14913_14741# a_14747_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3796 vccd1 a_25842_25589# a_25769_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3798 vssd1 a_12927_3829# a_12885_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3800 a_20004_15279# a_19605_15279# a_19878_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3801 a_14524_6549# _0531_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3802 a_19439_12015# _0894_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3803 temp1.capload\[7\].cap.Y temp1.capload\[7\].cap.A a_14373_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3804 a_17217_2767# _0622_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3805 a_7607_3855# a_6909_3861# a_7350_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3806 a_2214_4765# a_1775_4399# a_2129_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3807 a_21886_2335# a_21718_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3808 vssd1 a_15795_27791# a_15963_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3809 a_7385_27247# _0837_.A1 _0837_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3810 a_14736_24847# _0445_.B a_14433_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3812 _0963_.D a_20471_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3813 a_1945_9295# _1084_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X3815 a_14195_11471# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3820 a_21166_27613# a_20727_27247# a_21081_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3821 vccd1 a_24887_22325# a_24803_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3822 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3823 a_21886_2335# a_21718_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3824 vssd1 _0489_.X a_19439_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3826 vccd1 a_22587_22075# a_22503_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3827 vssd1 _0506_.A2 a_20245_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3828 a_26551_26525# a_25769_26159# a_26467_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3829 a_8155_16161# _0807_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3831 a_12018_17027# _0813_.A2 a_11936_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3833 vccd1 _0778_.A2 a_7203_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
R11 temp1.capload\[11\].cap_41.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3835 a_5823_28585# _0833_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3836 vssd1 _0761_.B a_6929_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3837 a_6612_8181# _0681_.X a_6832_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3838 a_1975_29967# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X3841 _0752_.Y _0444_.B a_6559_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3842 vccd1 _0558_.A2 a_24949_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3843 a_4356_23983# _0752_.Y io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3845 _0563_.C1 a_24591_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3846 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3847 vssd1 a_14710_20149# a_14668_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3848 vssd1 a_9003_15797# _0636_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3849 vssd1 _1078_.Q a_14287_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X3850 a_11149_19631# _0850_.A a_11067_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X3851 vccd1 _0745_.A2 a_6833_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3854 a_17470_10357# a_17302_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3855 _0954_.Q a_12743_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3856 a_11685_25045# _0825_.A1 a_11842_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3857 _0443_.A a_10789_22071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X3859 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3860 a_12441_17705# _0798_.A2 _0751_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3861 vccd1 a_15630_16479# a_15557_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3862 vssd1 _0922_.CLK a_9411_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3863 a_15016_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3864 a_10488_27497# a_10239_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3865 a_13840_5321# a_13441_4949# a_13714_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3866 a_23224_8751# a_22825_8751# a_23098_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3867 _0684_.A2 _0475_.X a_9217_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3868 a_27387_13469# a_26523_13103# a_27130_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3870 a_5813_25117# _0850_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3871 a_16937_19631# a_16771_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3872 a_22822_19087# a_22549_19093# a_22737_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3873 a_27422_5853# a_27149_5487# a_27337_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3874 _0945_.D a_17987_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3875 a_10564_20407# a_10714_20541# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X3876 _0845_.Y _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3877 a_6559_23552# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3878 a_21721_21807# a_21555_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3879 a_19973_7663# a_19807_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3880 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8464_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3883 vssd1 _0511_.D a_14875_18589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X3884 _0813_.A2 a_4132_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3886 a_9941_17289# a_8951_16917# a_9815_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3887 vccd1 _0999_.CLK a_23211_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3889 vccd1 _0583_.A a_23303_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3891 vccd1 _0577_.C a_15667_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3892 a_16685_11177# _0991_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3893 vccd1 a_5142_4511# a_5069_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3894 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_4811_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3896 vccd1 a_22659_19631# _0999_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3897 a_27057_13469# a_26523_13103# a_26962_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3898 a_17853_3145# a_16863_2773# a_17727_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3899 a_20145_5309# _0632_.B a_20073_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3900 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_11527_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3901 a_26183_14735# a_25401_14741# a_26099_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3902 a_21581_14219# _0842_.A0 a_21495_14219# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3903 a_9398_10383# _0475_.X a_9095_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X3904 vssd1 a_3270_2741# _0850_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X3905 vccd1 _0524_.X a_11711_1792# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3908 a_10068_11849# a_9669_11477# a_9942_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3909 vccd1 a_24075_21263# a_24243_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3910 vccd1 _0922_.CLK a_1959_4951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3911 _1076_.Q a_2991_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3912 vssd1 _0722_.A a_2975_17461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3913 vccd1 _0668_.X a_15641_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3915 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3916 vssd1 _0849_.X a_12433_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3917 vssd1 a_24075_21263# a_24243_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3919 _1034_.Q a_26175_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3920 a_6437_20719# _0869_.B1 a_6365_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3921 _0628_.X a_15667_15936# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3922 vccd1 _0959_.CLK a_9871_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3923 vssd1 a_16826_26271# a_16784_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3925 vccd1 a_22622_1653# a_22549_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3926 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3927 a_10294_22325# a_10126_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3928 vssd1 a_13203_21237# a_13161_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3929 vccd1 ANTENNA_7.DIODE a_3799_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3930 vccd1 a_3083_25339# a_2999_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3931 a_16929_17973# _0522_.B1 a_17086_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3932 a_18605_2473# _0594_.C a_18509_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3933 _0673_.B2 a_4831_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3934 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_7564_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3935 a_15285_27791# _1053_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3936 vssd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_2686_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3937 vssd1 a_23523_9117# a_23691_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3938 vccd1 _0844_.B a_3167_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X3939 a_2956_1956# a_2762_1801# a_3132_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.0687 ps=0.76 w=0.36 l=0.15
X3940 a_15563_9295# _0651_.X _0684_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3943 vssd1 a_16090_20831# a_16048_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3945 a_9911_12061# a_9595_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X3946 vccd1 _0752_.Y a_1591_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3947 vccd1 a_27590_24095# a_27517_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3948 vssd1 a_4132_17429# _0813_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3949 vssd1 a_20195_3829# a_20153_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3950 a_20521_3145# a_19531_2773# a_20395_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3951 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3952 vssd1 _0850_.Y a_14736_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3955 a_27590_12127# a_27422_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3956 a_6553_17705# _0812_.A2 _0749_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3957 vssd1 a_9963_17455# _0511_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3958 vccd1 a_23247_14557# a_23415_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3959 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3960 vssd1 a_19183_4917# a_19141_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3961 a_23515_7119# a_22733_7125# a_23431_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3962 vssd1 a_3451_25589# _1078_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3964 vssd1 _0580_.X a_19439_12675# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3965 a_12763_12879# _0833_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3966 vccd1 _0803_.X a_4843_19659# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3968 a_7544_25077# _0845_.A1 a_7472_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3969 a_11798_24847# _0847_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X3970 a_18274_7913# _0633_.X a_18025_7809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3971 _0652_.A a_15671_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X3973 a_8914_7093# a_8746_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3974 vccd1 a_20393_8545# _0523_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X3975 a_27422_10205# a_26983_9839# a_27337_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3976 a_26041_17455# a_25051_17455# a_25915_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3977 a_21568_13103# a_21169_13103# a_21442_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3978 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3979 a_8464_26409# a_8215_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3980 io_out[5] a_6611_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3981 a_20819_16617# _0564_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X3982 _0605_.D1 a_13367_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3983 vssd1 _0523_.B1 a_22729_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X3984 vssd1 _0722_.C _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3985 _0880_.A1 a_8155_16161# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3986 vccd1 a_4847_28701# a_5015_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3987 a_14139_4943# a_13441_4949# a_13882_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3988 a_17727_10383# a_17029_10389# a_17470_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3989 a_8292_14441# _0768_.B1 a_8037_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3990 a_3993_29673# _0845_.B1 a_4248_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3991 vccd1 a_25623_4667# a_25539_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3994 a_2340_4399# a_1941_4399# a_2214_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3995 a_6807_11177# _0746_.A2 a_6735_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3996 _0488_.B2 a_24335_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3997 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12355_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3998 vccd1 _0439_.A a_5797_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3999 vssd1 _0655_.X _0680_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4001 a_26961_10927# a_25971_10927# a_26835_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4002 _0583_.X a_20083_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4004 _0928_.D a_28015_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4005 _0758_.A1 a_3028_14165# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4006 vccd1 a_16035_4943# _1030_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4007 vssd1 a_10202_13621# a_10160_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4008 vssd1 _0505_.A2 a_26041_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4009 a_25789_25321# _0854_.B a_25707_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4010 a_20345_22351# _0932_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4011 a_25309_6037# a_25143_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4012 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_12788_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4013 vssd1 _0816_.S temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4014 vccd1 _0837_.A1 a_9718_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4015 vccd1 a_16439_4765# a_16607_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4016 a_3226_26703# a_2787_26709# a_3141_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4017 a_1591_22057# _0444_.A io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4018 vssd1 a_6336_15253# _0760_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4019 a_14726_12381# a_14287_12015# a_14641_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4021 a_22940_15279# _0648_.B1 a_22449_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4023 a_27337_21807# _0998_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4024 a_4958_2741# a_4790_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
R12 vssd1 temp1.capload\[3\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4025 a_2686_23439# clkbuf_1_1__f__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4026 a_12065_6031# _0954_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4027 a_24075_21263# a_23211_21269# a_23818_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4029 vccd1 _0824_.Y a_13183_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4030 a_22181_15829# a_22015_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4031 a_25769_26159# a_25603_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4032 a_21213_17249# _0504_.A a_21127_17249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4033 a_18645_7457# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4034 a_9171_7119# a_8473_7125# a_8914_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4035 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4036 a_5547_17027# _0873_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4038 vssd1 _0677_.A1 a_7663_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4039 vccd1 a_11815_12265# _0475_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4041 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4043 a_2313_2223# _0858_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4044 _0445_.X a_5273_29687# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X4045 a_4901_13647# _0791_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4047 a_22369_20175# _1022_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4048 vssd1 a_25455_2589# a_25623_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4049 vccd1 _0844_.B a_4915_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4050 vccd1 _0789_.A2 a_6809_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4051 a_27149_25071# a_26983_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4053 vccd1 _0597_.A2_N a_9495_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X4054 _0926_.D a_23047_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4055 vssd1 a_23266_8863# a_23224_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4056 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4057 a_24719_20175# a_23855_20181# a_24462_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4058 vssd1 _0524_.X a_23457_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4059 vssd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4061 vccd1 _0801_.X a_13367_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4062 a_20911_1385# _0645_.B1 a_20993_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4063 _1029_.Q a_18539_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4064 a_16753_26525# a_16219_26159# a_16658_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4066 _0538_.B2 a_7775_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4068 a_16897_12897# _0583_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4069 a_11040_29967# a_10791_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4073 a_8205_13967# _0626_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4074 _0954_.D a_10811_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4075 a_10497_17999# _0749_.B2 a_10413_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4076 _0622_.B2 a_10167_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4077 a_7291_20175# _0798_.A2 a_7073_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X4079 a_17217_10383# _0983_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4080 a_22833_17455# _0583_.A a_22751_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4081 _0544_.D a_14839_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4083 vccd1 a_5659_4917# a_5575_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4084 a_22821_26159# a_21831_26159# a_22695_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4085 vccd1 temp1.capload\[9\].cap_54.LO temp1.capload\[9\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4086 vccd1 a_8803_4943# a_8971_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4087 a_6633_6575# a_6467_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4088 a_11929_9633# _0479_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4089 a_21721_21807# a_21555_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4090 vccd1 _1062_.CLK a_22659_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4091 a_24389_20175# a_23855_20181# a_24294_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4093 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4094 a_12625_14441# _0735_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X4095 vssd1 a_27590_21919# a_27548_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4096 vssd1 _1028_.CLK a_11711_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4097 vssd1 a_12375_15547# a_12333_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4098 a_2566_2335# a_2398_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4099 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4100 vssd1 _0502_.X a_19557_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4101 vssd1 _0475_.X a_9313_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4102 a_22169_14013# _0893_.D a_22097_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4103 a_7360_31055# a_7111_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4104 vssd1 fanout10.A a_10791_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4105 a_16182_14303# a_16014_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4107 _0812_.A2 a_1775_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4108 _0768_.B1 a_4165_14455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X4109 a_12723_3561# _0532_.A2 a_12805_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4110 io_out[6] a_5141_30199# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4111 vssd1 a_21667_20987# a_21625_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4113 a_20709_3311# a_20543_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4115 _0641_.D1 a_11711_1792# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X4117 a_18317_20181# a_18151_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
R13 vssd1 temp1.capload\[8\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4120 a_20522_21263# a_20083_21269# a_20437_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4121 a_18758_4917# a_18590_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4122 vccd1 _1033_.CLK a_22567_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4123 a_27973_23983# a_26983_23983# a_27847_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4125 a_8479_16367# _0837_.A1 _0735_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X4126 a_12521_4399# a_12355_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4127 a_21166_27613# a_20893_27247# a_21081_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4128 a_12725_19087# _0866_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4129 a_23303_16617# _0648_.B1 a_23385_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4130 vccd1 a_8235_4667# a_8151_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4132 a_13161_21641# a_12171_21269# a_13035_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4133 vccd1 a_25807_8181# a_25723_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4135 vccd1 a_2455_9295# a_2626_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X4136 vssd1 a_24059_17973# a_24017_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4137 _1019_.Q a_21759_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4138 vssd1 _0472_.X _0518_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4140 a_25221_6575# _1003_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4141 a_16984_15529# _0577_.X a_16882_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4142 a_12613_2773# a_12447_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4143 vssd1 _0964_.CLK a_26983_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4145 vccd1 clkbuf_1_1__f_net57.A a_1674_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4146 a_17010_21919# a_16842_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4147 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A a_8464_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4149 a_16014_4765# a_15575_4399# a_15929_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4150 a_26689_13103# a_26523_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4151 vccd1 _0791_.A2 a_4901_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4152 a_21123_5853# a_20341_5487# a_21039_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4153 _0907_.Q a_8327_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4154 io_out[4] _0774_.A2 a_4439_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4155 vssd1 _0975_.CLK a_23855_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4156 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4157 a_4035_9813# _0807_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X4158 vccd1 _1019_.CLK a_19991_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4159 vccd1 _0959_.CLK a_14839_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4161 a_20299_12043# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4162 a_5820_14191# _0734_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X4163 vssd1 a_27739_6843# a_27697_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4164 a_27548_9839# a_27149_9839# a_27422_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4165 a_4882_19087# a_4705_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4166 vccd1 _0814_.A2 a_4065_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4167 _0845_.Y _0845_.A1 a_4441_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4168 vssd1 _1079_.Q a_9411_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4169 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE _0827_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4170 _0850_.A a_3270_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4171 vssd1 _1033_.CLK a_22751_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4172 vccd1 a_20855_22351# a_21023_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4173 a_11417_3677# a_10883_3311# a_11322_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4174 a_15588_16367# a_15189_16367# a_15462_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4176 a_12047_13103# _1076_.Q a_11956_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X4177 a_12995_16911# _0797_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4178 a_26870_4765# a_26431_4399# a_26785_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4179 vssd1 a_28015_12283# a_27973_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4181 a_2949_3311# a_1959_3311# a_2823_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4182 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4183 a_19617_9839# _0983_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4184 vssd1 a_20855_22351# a_21023_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4187 vssd1 a_21518_18655# a_21476_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4188 vccd1 _0764_.A1 a_6682_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4189 a_13261_10383# _0630_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4190 vccd1 _0999_.CLK a_22015_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4192 a_18555_11471# a_17857_11477# a_18298_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4193 vssd1 temp1.inv1_1.Y a_1766_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4194 vssd1 a_25707_25321# _0854_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4197 _0656_.Y _0655_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X4200 vssd1 _0868_.A2 a_6916_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4201 a_19605_15279# a_19439_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4203 _1053_.CLK a_8307_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4205 vssd1 _1080_.Q _0845_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4206 a_21533_4399# a_20543_4399# a_21407_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4208 a_27513_11791# _1068_.Q a_27167_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4209 a_9497_13353# _0735_.A2 _0747_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4210 a_22580_17289# a_22181_16917# a_22454_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4211 a_10183_12061# _0836_.A a_10083_12061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X4212 temp1.inv1_1.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4213 vccd1 a_16826_26271# a_16753_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4214 vssd1 a_13514_22325# a_13472_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4215 a_15101_14735# _0924_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4216 vccd1 a_11287_11293# a_11455_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4217 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11040_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4220 vssd1 _0444_.Y a_5428_29429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
X4221 a_22779_26525# a_21997_26159# a_22695_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4222 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4223 vccd1 _1075_.Q a_7939_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4224 a_8378_4943# a_8105_4949# a_8293_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4225 a_9558_16885# a_9390_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4226 vssd1 a_15354_14709# a_15312_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4227 a_25589_1135# _0552_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4229 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4230 a_9489_1135# _0646_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4231 a_25815_6941# a_25033_6575# a_25731_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4233 a_6427_11989# _0758_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X4234 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4235 a_15943_13760# _1050_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4236 vssd1 a_5015_1403# a_4973_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4237 vccd1 a_27590_5599# a_27517_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4238 vccd1 a_7258_5599# a_7185_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4239 vssd1 _0460_.C a_1945_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4240 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4242 a_20175_7119# _0516_.B1 a_20257_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4243 a_9547_25071# _0825_.A0 a_9184_25223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4244 _0814_.A1 clkbuf_1_1__f_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4246 a_24251_9295# a_23469_9301# a_24167_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4247 a_26007_12381# a_25143_12015# a_25750_12127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4248 a_25915_8029# a_25217_7663# a_25658_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4250 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_7360_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4252 vssd1 _1062_.CLK a_22659_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4253 a_2455_6031# a_1591_6037# a_2198_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4254 vccd1 a_28015_10107# a_27931_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4256 vccd1 temp1.capload\[0\].cap.A temp1.capload\[0\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4257 vccd1 _0845_.A2 a_4248_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4259 a_4382_17027# _0872_.A1 a_4300_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4260 vccd1 a_5215_2767# a_5383_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4261 vccd1 a_9095_20407# _0459_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X4262 vccd1 _0440_.A a_4249_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4263 vssd1 a_16439_4765# a_16607_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4264 vssd1 _0959_.CLK a_9779_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4265 a_2122_12015# a_1945_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X4266 vccd1 a_9503_19087# _0471_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4267 a_11316_27497# a_11067_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4268 _0662_.A1 a_18611_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4269 a_27981_4943# a_27804_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X4270 a_25589_10383# _1006_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4271 a_24113_2773# a_23947_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4272 a_25677_12381# a_25143_12015# a_25582_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4273 a_2030_6031# a_1591_6037# a_1945_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4274 vssd1 _0445_.A a_9897_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4275 a_17236_6575# _0645_.B1 a_16745_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4276 vccd1 _0662_.A3 a_15943_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4277 vssd1 a_13311_2767# a_13479_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4279 _0934_.Q a_17435_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4280 vssd1 _1053_.CLK a_7663_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4281 a_9312_14191# _0714_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.069875 pd=0.865 as=0.105625 ps=0.975 w=0.65 l=0.15
X4282 a_21134_11177# _1063_.Q a_20977_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4283 vssd1 a_12207_21085# a_12375_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4284 a_17221_18543# _0583_.A a_17139_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4285 a_22622_20149# a_22454_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4286 a_5823_28585# _0845_.A2 _0833_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4287 a_12575_6031# a_11877_6037# a_12318_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4288 vccd1 _0654_.Y _0768_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X4289 a_2033_27069# _0847_.A2 a_1933_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X4290 vssd1 a_6779_2589# a_6947_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4291 a_25723_12559# a_24941_12565# a_25639_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4292 a_20625_9839# _0504_.A a_20543_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4293 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_5639_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4294 a_14689_18589# a_14287_18543# a_14603_18589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X4295 a_27517_16733# a_26983_16367# a_27422_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4296 vccd1 a_11435_8751# _0842_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4297 vccd1 fanout13.A a_10977_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4298 vssd1 a_17378_19743# a_17336_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4300 vssd1 a_18187_6031# a_18355_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4303 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4304 vccd1 a_10110_21237# a_10037_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4305 a_16548_10901# _0565_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4306 a_23466_26703# a_23027_26709# a_23381_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4307 a_27931_15645# a_27149_15279# a_27847_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4308 a_10735_2589# a_10037_2223# a_10478_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4309 _0588_.A1 a_15319_12283# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4310 a_3129_17705# _0456_.B a_3057_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X4311 a_18087_12043# _0504_.A a_18001_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4312 a_16140_4399# a_15741_4399# a_16014_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4313 vccd1 a_4590_28447# a_4517_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4315 a_25309_9839# a_25143_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4316 vccd1 a_12743_11445# a_12659_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4318 vssd1 a_27590_9951# a_27548_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4319 vssd1 _0471_.X _0840_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X4320 vssd1 _0533_.X a_18600_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X4321 a_16565_7663# _1059_.D a_16127_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4324 vccd1 _0698_.B1 a_4621_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4326 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4327 vccd1 _1028_.CLK a_9227_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4328 vssd1 a_4590_26271# a_4548_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4329 a_7435_26324# _0817_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4330 a_2984_25993# a_2585_25621# a_2858_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4331 a_4931_2589# a_4149_2223# a_4847_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4332 vssd1 a_19827_1653# a_19785_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4335 vssd1 _0964_.CLK a_25235_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4339 a_20717_1679# _0645_.B1 a_20801_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4340 a_26996_4399# a_26597_4399# a_26870_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4341 a_25800_25993# a_25401_25621# a_25674_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4342 a_15186_3677# a_14747_3311# a_15101_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4343 a_19521_9001# _0517_.D a_19439_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X4344 vssd1 _0798_.A2 a_4414_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
X4345 vssd1 _0827_.A _0824_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4346 vccd1 _0511_.D a_14287_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4347 vccd1 _0975_.CLK a_24591_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4349 vssd1 a_9227_17455# _0995_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4350 a_25658_7775# a_25490_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4351 vccd1 a_11765_22325# _0858_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4353 _0505_.A2 a_19471_6603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4354 vccd1 a_2991_1403# _0840_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4355 a_25581_15279# a_24591_15279# a_25455_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4356 vccd1 a_23523_9117# a_23691_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4357 a_14894_12127# a_14726_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4359 a_14319_20747# _0829_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4360 _0652_.C a_12631_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4362 vccd1 _0922_.CLK a_9411_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4363 a_5081_23439# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4364 a_7185_5853# a_6651_5487# a_7090_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4365 a_18072_10927# a_17673_10927# a_17946_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4367 vccd1 clkbuf_1_1__f_net57.A a_1674_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4368 vccd1 a_19773_18689# _0584_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X4370 a_14825_17999# _1056_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4371 vssd1 _0761_.B a_9313_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4373 a_25677_6031# a_25143_6037# a_25582_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4374 a_13169_9295# _1026_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4376 a_15115_9295# _0652_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4378 _0749_.A1 _0835_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4379 a_15128_4233# a_14729_3861# a_15002_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4380 a_23487_6825# _0619_.B1 a_23569_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4381 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4383 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_7111_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4384 _0445_.A _0869_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4386 vccd1 _0845_.A1 _0866_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4387 a_19885_2767# _0970_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4388 vccd1 a_26267_16885# a_26183_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4389 a_15695_3677# a_14913_3311# a_15611_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4390 a_21994_22173# a_21721_21807# a_21909_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4391 vccd1 a_27847_24349# a_28015_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4393 a_19015_4943# a_18151_4949# a_18758_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4394 a_11601_9839# a_11435_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4395 _0564_.X a_20819_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X4396 a_7393_17705# _0869_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4397 a_3885_24847# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4399 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4401 vssd1 a_24811_2767# a_24979_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4402 a_6549_9001# _0657_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X4403 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11316_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4404 vccd1 _0815_.Y a_14011_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4405 a_20797_15113# a_19807_14741# a_20671_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4406 _0819_.S _0444_.B a_10055_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4407 a_5621_3311# a_5455_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4408 vssd1 a_12777_24501# fanout13.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4409 vccd1 a_15335_17999# a_15503_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4410 a_10401_4399# a_9411_4399# a_10275_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4411 a_2686_31055# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4413 vssd1 _0994_.CLK a_23855_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4414 a_8021_18793# _0798_.A2 a_7939_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4415 a_18497_1135# a_17507_1135# a_18371_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4422 a_25674_1501# a_25235_1135# a_25589_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4423 a_2129_4399# _0870_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4427 a_9574_1501# a_9135_1135# a_9489_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4428 a_4847_26525# a_3983_26159# a_4590_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4429 vssd1 a_3302_4917# a_3260_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4430 a_19709_11791# _0962_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4431 a_23266_4511# a_23098_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4432 a_9301_14441# _0714_.B2 a_9217_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4433 _0479_.Y _1079_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4435 a_2156_6409# a_1757_6037# a_2030_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4436 vssd1 a_26210_26271# a_26168_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4437 vccd1 _0745_.A1 _0713_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X4438 a_15277_7663# a_14287_7663# a_15151_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4439 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12355_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4440 a_20479_8545# _0582_.A a_20393_8545# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4441 a_12981_15823# a_12447_15829# a_12886_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4443 a_14729_3861# a_14563_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4444 a_18961_1685# a_18795_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4445 a_21809_8751# a_20819_8751# a_21683_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4446 vccd1 a_16863_11479# fanout27.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4447 vccd1 a_25731_6941# a_25899_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4449 a_21169_23983# a_21003_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4450 vssd1 a_22449_15253# _0561_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4451 vccd1 _0521_.A a_13551_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4452 a_13183_7232# _0611_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4453 a_2198_9269# a_2039_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4454 a_21127_11809# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4457 vccd1 _0908_.CLK a_7203_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4459 vssd1 fanout10.A a_10975_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4460 _0440_.C a_5547_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X4461 _0897_.Q a_18723_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4462 _0967_.Q a_26267_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4463 vccd1 a_16607_14459# a_16523_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4464 a_19439_4399# _0630_.A2 a_19617_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4465 a_1757_5487# a_1591_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4466 vccd1 _0655_.X a_7203_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X4468 vssd1 a_13367_17999# _0866_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4469 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4471 vssd1 a_3651_26703# a_3819_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4472 a_20989_20719# _1048_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4473 a_9583_15055# _0829_.A1 _0770_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X4474 a_13717_6031# _0538_.B2 a_13633_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4475 a_26183_19997# a_25401_19631# a_26099_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4477 a_11693_6825# _0921_.Q a_11609_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4478 _0897_.Q a_18723_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4479 _0725_.A a_3983_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4480 vssd1 _0506_.A2 a_20613_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4481 a_1639_7828# io_in[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4482 _1028_.CLK a_9135_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4483 _1031_.Q a_23783_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4484 a_2490_25437# a_2217_25071# a_2405_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4485 a_13441_4949# a_13275_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4487 vssd1 _0471_.X _0529_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4488 vccd1 _1019_.CLK a_18335_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4489 a_14655_2767# _0670_.A2 a_14737_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4491 vssd1 _1053_.CLK a_12907_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4492 vccd1 _0995_.CLK a_19439_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4493 a_4701_4399# a_4535_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4494 vccd1 a_26099_14735# a_26267_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R14 temp1.capload\[15\].cap_45.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4496 a_25539_15645# a_24757_15279# a_25455_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4498 vccd1 a_11950_15391# a_11877_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4499 vccd1 a_22143_2589# a_22311_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4500 a_23615_8207# a_22751_8213# a_23358_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4501 _0504_.A a_18703_12567# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4502 _0685_.X a_6651_12672# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X4503 vccd1 _0582_.A a_22015_18112# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4504 a_9497_14735# _0461_.A _0770_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4505 a_9850_4765# a_9577_4399# a_9765_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4507 vssd1 _0935_.CLK a_14747_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4509 a_10769_3145# a_9779_2773# a_10643_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4511 a_14457_20175# _0919_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4512 a_15312_3311# a_14913_3311# a_15186_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4513 a_8399_19407# _0763_.A2 a_8305_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4514 a_4422_26525# a_4149_26159# a_4337_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4515 a_20257_7119# _0649_.B2 a_20175_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4516 a_7843_14735# _0735_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4518 a_27847_2589# a_26983_2223# a_27590_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4519 a_21127_12043# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4520 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4521 a_25340_23817# a_24941_23445# a_25214_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4522 a_15335_17999# a_14471_18005# a_15078_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4523 _0845_.A1 a_2991_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4524 vccd1 _1015_.CLK a_23303_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4525 vccd1 _0696_.A1 a_4338_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X4527 _1024_.Q a_21851_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4528 a_10133_2767# _0673_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4529 vccd1 _0917_.CLK a_9319_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4530 _0671_.B2 a_20195_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4531 a_26467_26525# a_25603_26159# a_26210_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4534 vssd1 a_23910_9269# a_23868_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4536 vssd1 a_9926_9269# a_9884_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4537 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10416_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4538 a_15189_16367# a_15023_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4539 vssd1 a_27130_13215# a_27088_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4540 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4541 vssd1 a_2455_9117# a_2623_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4542 vccd1 _0563_.B1 a_27249_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4544 vccd1 _0833_.A a_5823_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X4545 a_6929_18543# a_6646_18865# a_6516_18695# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4546 vccd1 _0479_.Y a_14655_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4547 _0685_.B a_9284_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X4548 a_17401_17455# _1059_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4549 a_9390_16911# a_8951_16917# a_9305_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4550 vssd1 _0797_.A1 a_6287_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4552 a_3026_25589# a_2858_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4553 a_12604_26409# a_12355_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4554 vccd1 a_8546_4917# a_8473_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4556 a_18213_17277# _1061_.Q a_18141_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4557 _0842_.A0 a_11435_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4558 vccd1 a_16182_14303# a_16109_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4559 a_26137_26525# a_25603_26159# a_26042_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4560 a_2658_25183# a_2490_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4562 vccd1 a_3819_26677# _1075_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4564 _0874_.X a_4300_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4565 _0840_.A0 _0471_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4566 vssd1 a_21575_4667# a_21533_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4567 vssd1 a_25455_15645# a_25623_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4568 vccd1 _1019_.CLK a_21279_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4571 a_16829_12161# _0565_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X4573 io_out[1] a_4403_22869# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4574 a_9857_21263# _0988_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4575 a_8944_30287# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4576 a_17585_22895# _0932_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4578 a_9993_9839# _0545_.B2 a_10084_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4579 vssd1 _0583_.A a_19439_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4580 a_22097_18365# _0582_.A a_22015_18112# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4581 vssd1 _0791_.A3 a_5639_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4582 vccd1 a_2623_6005# a_2539_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4585 a_24110_11471# a_23671_11477# a_24025_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4586 _0791_.A1 _0745_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4587 a_9919_6740# _0854_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4589 a_16204_6031# _0565_.B1 a_15949_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4590 a_25800_1135# a_25401_1135# a_25674_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4592 _0809_.B2 a_3155_21271# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4593 _0872_.Y a_3141_19148# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X4594 a_7182_3855# a_6743_3861# a_7097_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4595 a_9700_1135# a_9301_1135# a_9574_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4596 a_5902_6031# _0680_.Y a_5599_6263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X4597 a_26091_10205# a_25309_9839# a_26007_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4598 a_21442_24349# a_21003_23983# a_21357_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4599 _0679_.A1 _0676_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4600 a_10594_15823# _0836_.A a_10397_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4601 a_7192_27497# _0845_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4602 a_27011_21085# a_26229_20719# a_26927_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4603 vssd1 a_12962_4511# a_12920_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4604 a_2566_27359# a_2398_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4606 _0508_.Y _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4607 vssd1 _0618_.C1 a_22751_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4608 a_5904_18543# _0783_.A1 a_5601_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4609 a_26099_14735# a_25235_14741# a_25842_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4610 vssd1 _0873_.A a_4300_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4611 vssd1 a_26099_3855# a_26267_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4612 a_11711_24527# _0840_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4613 a_2122_3855# a_1849_3861# a_2037_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4614 a_19709_16367# _0920_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4616 a_19689_9269# _0533_.X a_19846_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4618 a_22291_16617# _0643_.B1 a_22373_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4619 a_27149_3311# a_26983_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4620 a_10677_6409# a_9687_6037# a_10551_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4621 _0566_.B1 a_15115_5059# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X4622 a_16908_6575# _0662_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X4623 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8188_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4625 vccd1 _0602_.A a_18703_12567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4626 a_4065_31849# _0814_.B2 a_3983_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4627 _0854_.B a_11895_1385# a_12428_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4629 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4630 vccd1 a_25842_19061# a_25769_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4631 a_24696_14025# a_24297_13653# a_24570_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4632 vssd1 a_4403_22869# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4633 a_4250_10927# _0698_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X4634 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4635 vccd1 _0619_.X a_22653_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4636 a_24757_16367# a_24591_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4637 vccd1 _0814_.A2 a_2039_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4639 a_15005_17277# _1076_.Q a_14905_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X4640 vssd1 fanout23.X a_26983_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4641 vccd1 a_5323_29111# _0764_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X4643 _1078_.Q a_3451_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4644 a_20348_18543# _0934_.Q a_19773_18689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X4645 vssd1 _0558_.A2 a_24017_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X4646 a_10018_4511# a_9850_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4647 vccd1 _0821_.Y a_7755_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4648 a_23247_14557# a_22549_14191# a_22990_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4649 a_13219_4765# a_12521_4399# a_12962_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4650 vccd1 _0471_.X a_9911_12061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X4651 _0994_.D a_26267_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4653 a_23098_9117# a_22825_8751# a_23013_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4654 vssd1 a_5273_29687# _0445_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4655 _1078_.Q a_3451_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4658 a_27038_4511# a_26870_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4660 a_4843_19659# _0440_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4661 a_15380_10703# _0613_.A1 a_14805_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X4662 a_2405_28335# _0845_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4663 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_10033_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4664 _0629_.X a_18059_17024# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X4665 vccd1 _0768_.A2 a_8037_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4666 a_7006_16911# a_7226_16885# _0518_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4668 a_3993_29673# _0845_.C1 _0845_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4669 _0994_.D a_26267_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4670 a_19605_15279# a_19439_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4671 a_7520_23555# _0441_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4672 vssd1 _0773_.A2_N a_10714_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4673 vccd1 _0680_.Y _0710_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4674 a_21074_21085# a_20801_20719# a_20989_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4675 a_15285_1679# _1042_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4676 _0549_.C1 a_20267_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4678 a_15693_15307# _0521_.A a_15607_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4679 _0517_.D a_21647_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X4680 vssd1 _0662_.A3 a_14809_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4681 vccd1 _0513_.X a_15793_6603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4682 vssd1 fanout37.A a_16863_11479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4683 a_20981_22729# a_19991_22357# a_20855_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4684 _0999_.Q a_28015_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4685 _0798_.A2 _0722_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4686 vssd1 a_15354_3423# a_15312_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4688 a_4439_24233# _0814_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4689 a_13533_17455# _1078_.Q a_13433_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X4690 _0880_.A2 _0807_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4691 a_27337_9839# _0572_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4692 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4693 a_16902_6825# _0662_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X4694 vssd1 _0538_.C1 a_13551_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4695 a_8473_4943# a_7939_4949# a_8378_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4696 a_25225_9295# _0664_.X a_25143_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4697 a_22974_18793# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4701 a_2686_23439# clkbuf_1_1__f__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4702 a_26099_1501# a_25401_1135# a_25842_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4703 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_12604_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4704 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4706 a_15741_14191# a_15575_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4707 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4708 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A a_8004_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4709 vssd1 _0847_.A3 a_5466_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X4711 _0848_.X a_12547_23145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X4712 vccd1 a_8545_14709# _0546_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4713 a_25511_11471# _0664_.A2 a_25593_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4714 a_25800_16201# a_25401_15829# a_25674_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4715 vccd1 _1053_.CLK a_9503_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4716 _0648_.X a_23303_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4718 _0926_.D a_23047_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4721 a_23005_20553# a_22015_20181# a_22879_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4722 a_18405_3311# a_17415_3311# a_18279_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4723 a_12291_21085# a_11509_20719# a_12207_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4724 a_7074_6687# a_6906_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4726 vccd1 _0721_.A a_3155_21271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4728 vccd1 _0964_.CLK a_22015_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4729 a_4901_13647# _0791_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4731 a_27061_6575# _0562_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4732 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4733 vssd1 a_7435_26324# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4734 vssd1 _0460_.C a_2879_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X4737 _0662_.B1 a_21127_17249# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4738 a_11977_27497# fanout11.A fanout9.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4739 a_7074_6687# a_6906_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4740 vccd1 a_4958_2741# a_4885_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4741 _0684_.A1 _0652_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4742 vccd1 _0670_.A2 a_13165_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4744 a_9769_19881# _0798_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4746 a_13309_5515# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4747 a_6809_25615# _0787_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4748 vccd1 a_19659_1679# a_19827_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4749 vssd1 _0722_.C _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4750 vccd1 a_22879_15823# a_23047_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4751 a_24017_15055# _0999_.Q a_23579_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4752 a_7745_12559# _0684_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4753 a_18088_13647# _0606_.X a_17986_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4755 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4756 a_13360_27023# _0824_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4757 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10876_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4758 vccd1 a_26743_23261# a_26911_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4761 a_25217_8751# a_25051_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4763 vccd1 _0445_.X a_9779_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4764 a_5639_16367# _0873_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4765 a_27337_16367# _1012_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4766 vccd1 a_18371_11293# a_18539_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4768 a_10386_4917# a_10218_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4769 a_25217_7663# a_25051_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4770 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4771 a_17393_21807# a_16403_21807# a_17267_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4772 vssd1 a_23891_26703# a_24059_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4773 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4774 vccd1 a_8031_16911# _0836_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4775 a_12962_4511# a_12794_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4777 a_3367_25615# a_2585_25621# a_3283_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4778 a_21150_3423# a_20982_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4779 a_24293_6409# a_23303_6037# a_24167_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4780 a_23837_11477# a_23671_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4781 a_7308_4233# a_6909_3861# a_7182_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4782 temp1.capload\[9\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4783 clkbuf_0_temp1.i_precharge_n.A a_9779_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4784 a_26183_25615# a_25401_25621# a_26099_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4785 a_23097_3145# a_22107_2773# a_22971_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4787 vssd1 a_3083_25339# a_3041_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4788 _0761_.X a_9636_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4789 vccd1 _0845_.C1 a_11068_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4790 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A _0825_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4792 vccd1 _0873_.A a_4382_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4794 a_11685_25045# _0829_.A1 a_11938_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X4795 a_12318_13621# a_12150_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4796 vccd1 a_13309_5515# _0515_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X4797 a_23082_20831# a_22914_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4798 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_15667_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4799 a_19521_12015# _0582_.A a_19439_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4801 vssd1 _0553_.C1 a_18243_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4802 a_8393_9615# _0679_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4803 vccd1 a_18001_12043# _0667_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X4804 a_11908_15279# a_11509_15279# a_11782_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4805 a_15611_14735# a_14913_14741# a_15354_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4809 a_19045_15797# _0658_.B1 a_19202_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4810 a_19329_6037# a_19163_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4813 vccd1 a_20027_3855# a_20195_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4814 vssd1 a_6427_11989# _0768_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4815 a_17293_18543# _1054_.Q a_17221_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4816 a_3049_4943# _0673_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4819 a_10294_6005# a_10126_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4820 a_15097_1685# a_14931_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4821 _1017_.D a_23415_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4822 vccd1 clkbuf_1_1__f_net57.A a_1674_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4824 vccd1 _0814_.A2 a_4439_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4825 a_6817_5487# a_6651_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4826 a_13080_17231# _0836_.A a_12777_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4827 vssd1 a_25382_12533# a_25340_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4828 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X4829 a_6556_15279# _0758_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X4831 vccd1 a_8325_11769# a_8355_11510# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4832 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_13183_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4833 a_10221_22351# a_9687_22357# a_10126_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4834 vssd1 _0722_.C a_5642_19637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4835 a_6909_3861# a_6743_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4837 a_21169_13103# a_21003_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4838 _0648_.B1 a_21495_14219# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4839 vccd1 io_in[7] a_1591_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4840 vccd1 a_11068_16617# _0882_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4841 _0483_.X a_15115_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4842 a_4035_25045# _0829_.A1 a_4262_25393# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4843 a_17811_2767# a_17029_2773# a_17727_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4844 a_17301_7439# _1029_.Q a_16863_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4845 vccd1 a_5509_7093# _0695_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4846 vccd1 a_23783_8181# a_23699_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4849 vccd1 a_10202_13621# a_10129_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4850 a_16745_6549# _0645_.B1 a_16902_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4851 vssd1 a_20839_14709# a_20797_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4852 vccd1 _0456_.A a_5549_17719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4853 vccd1 a_24995_13647# a_25163_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4854 _0970_.Q a_17895_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4855 vssd1 a_2991_1403# _0840_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4858 vssd1 _0506_.X a_19439_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X4860 a_12249_3855# _0956_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4862 vssd1 _0572_.A2 a_22361_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4863 _0666_.X a_21831_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4864 vssd1 _0888_.CLK a_2695_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4865 vssd1 a_24995_13647# a_25163_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4867 vccd1 a_10564_20407# _0774_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X4868 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11888_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4871 vccd1 a_27590_17567# a_27517_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4872 a_22612_15279# _0662_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X4873 _1033_.CLK a_22015_8215# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4874 a_6646_18865# _0795_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X4875 _0611_.B a_5199_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4876 a_4885_2767# a_4351_2773# a_4790_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4877 a_27548_12015# a_27149_12015# a_27422_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4878 _0861_.A1 _0860_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4880 vccd1 _0739_.A2 a_7477_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4881 a_20617_21263# a_20083_21269# a_20522_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4883 a_26785_4399# _1008_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4884 vccd1 _0866_.Y a_6831_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4885 vccd1 _1030_.CLK a_19807_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4886 _0825_.A0 _0825_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4887 a_27590_2335# a_27422_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4888 vccd1 a_20635_13655# _0583_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4889 vccd1 _1081_.Q a_1591_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4890 a_6645_6351# _0689_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4891 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_12532_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4892 vccd1 a_10719_22325# a_10635_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4893 a_6892_9001# _0680_.Y a_6549_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X4894 a_4864_15797# _0456_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4895 vccd1 _0838_.A0 a_9003_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X4896 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4897 _0505_.X a_22659_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4898 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4899 vssd1 a_27590_15391# a_27548_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4900 _1059_.D a_16607_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4901 _0845_.B1 _1080_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4902 a_25455_22173# a_24591_21807# a_25198_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4903 vccd1 _0717_.A2 a_10313_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4904 vssd1 a_18539_1403# a_18497_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4905 vssd1 _0869_.Y a_5173_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4906 a_6081_2223# a_5915_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4907 vssd1 _0685_.X a_6612_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4909 a_23657_9295# _0894_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
R15 vccd1 temp1.capload\[13\].cap_43.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4910 vssd1 a_26007_6031# a_26175_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4912 a_9673_9295# _0899_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4913 a_19602_26703# a_19163_26709# a_19517_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4915 a_21350_18909# a_21077_18543# a_21265_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4917 vccd1 a_17470_10357# a_17397_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4918 vssd1 a_15319_7931# a_15277_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4919 a_12441_32463# temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4920 a_16017_21085# a_15483_20719# a_15922_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4921 a_2599_16911# _0874_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4924 vssd1 _0833_.Y _0835_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4925 _0963_.Q a_23507_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4926 a_25842_16885# a_25674_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4927 a_6938_14237# _0717_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4928 vccd1 a_2626_9269# a_2539_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4930 vccd1 _0845_.A1 a_4248_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4931 vssd1 a_21851_9019# a_21809_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4933 _1079_.Q a_5015_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4934 a_18282_18793# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4935 vssd1 a_11747_3677# a_11915_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4936 a_15569_8323# _0675_.C a_15473_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4937 a_11704_28335# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4938 a_25673_13103# a_24683_13103# a_25547_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4939 a_16902_6825# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4940 _0662_.A1 a_18611_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4941 _0839_.Y _0839_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4942 a_20157_20181# a_19991_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4943 a_12068_22671# _0856_.Y a_11765_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4945 a_25674_16911# a_25401_16917# a_25589_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4947 a_25674_16911# a_25235_16917# a_25589_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4949 vccd1 _0722_.A a_4165_14455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X4950 a_11865_2045# _0905_.Q a_11793_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4951 a_18022_3423# a_17854_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4952 vccd1 a_2290_3829# a_2217_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4953 a_5721_16367# _0439_.A a_5639_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4954 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4955 a_10324_30511# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4956 a_10068_21641# a_9669_21269# a_9942_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4957 vssd1 _0471_.X _0574_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4959 vssd1 _1081_.Q a_10515_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X4960 a_2599_16911# _0861_.B1 a_2381_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X4961 vccd1 a_2455_9117# a_2623_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4962 _0745_.A3 _0776_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4963 a_13254_9295# a_12815_9301# a_13169_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4964 a_9897_22923# _0850_.A a_9811_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4967 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4968 vssd1 a_17267_22173# a_17435_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4969 _0808_.A a_6559_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4970 _0972_.CLK a_15667_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4972 a_27590_16479# a_27422_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4973 a_15017_32463# temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4975 vccd1 _0511_.D a_14603_18589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X4976 a_15841_1385# _1042_.Q a_15759_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4977 vssd1 a_7607_3855# a_7775_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4978 a_12709_4399# _0951_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4979 a_22097_5737# _1045_.D a_22015_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4980 _0833_.Y _0845_.A2 a_5823_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4981 vccd1 a_10294_22325# a_10221_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4983 a_6929_18543# _0829_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4984 a_10410_10383# _0475_.X a_10107_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X4986 a_27973_3311# a_26983_3311# a_27847_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4987 vssd1 a_13882_4917# a_13840_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4989 a_10777_10927# _0588_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4990 vccd1 _0972_.CLK a_16863_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4991 a_12659_13647# a_11877_13653# a_12575_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4992 a_4170_20291# _0722_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
R16 vccd1 temp1.capload\[5\].cap_50.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4993 vccd1 _0829_.A1 a_7025_18865# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4994 a_27847_15645# a_26983_15279# a_27590_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4995 vssd1 a_27755_9117# a_27923_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4996 vssd1 a_2626_9269# _0835_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X4997 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_6559_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4998 vccd1 a_23266_8863# a_23193_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4999 a_21683_19997# a_20985_19631# a_21426_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5001 _0624_.D_N _0620_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X5002 vccd1 a_15151_12381# a_15319_12283# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5003 a_4981_21024# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5004 vccd1 _0847_.A2 _0850_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5005 a_5599_6263# _0689_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X5006 a_18682_21263# a_18243_21269# a_18597_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
D1 vssd1 _0865_.Y sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X5008 a_24294_1679# a_24021_1685# a_24209_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5009 a_25309_12559# a_24775_12565# a_25214_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5010 a_6725_15823# _0735_.Y a_6641_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R17 temp1.dac.vdac_single.einvp_batch\[0\].vref.TE vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5012 a_19141_20553# a_18151_20181# a_19015_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5013 vssd1 a_20046_17567# a_20004_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5014 a_19613_11471# _0489_.C1 a_19531_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5015 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5016 a_11044_20541# fanout13.A a_10564_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5017 a_15189_16367# a_15023_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5018 a_15667_15936# _1055_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5019 vccd1 _0662_.A1 _0654_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5020 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5816_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5021 a_7164_14191# _0845_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5022 a_5264_20969# _0869_.Y _0870_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X5025 _0954_.Q a_12743_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5028 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5029 _0648_.A2 a_17909_16395# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X5030 vccd1 _0821_.Y a_8583_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5031 a_12893_1679# _0604_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5032 a_12575_6031# a_11711_6037# a_12318_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5033 a_8473_7125# a_8307_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5034 a_2398_2589# a_2125_2223# a_2313_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5035 vccd1 a_21759_27515# a_21675_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5036 a_2658_25183# a_2490_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5037 _0618_.C1 a_22015_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5038 _0831_.B clkbuf_1_0__f_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5039 _1040_.Q a_19183_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5041 vssd1 _0845_.A2 a_5177_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5042 vccd1 clkbuf_1_1__f_net57.A a_1674_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5045 vssd1 a_2915_25437# a_3083_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5046 vssd1 a_13571_1653# a_13529_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5047 a_15101_3311# _0946_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5049 a_12150_6031# a_11711_6037# a_12065_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5050 vssd1 a_4863_23413# _0814_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5051 vssd1 a_27571_6941# a_27739_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5052 _0574_.C _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5053 vccd1 a_24979_2741# a_24895_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5054 vssd1 fanout27.A a_17691_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5055 a_12176_25071# _0825_.A1 a_11685_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5057 _0710_.B1 a_4015_5515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5058 a_15151_10205# a_14453_9839# a_14894_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5059 vccd1 _0797_.A1 a_8105_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X5060 a_5737_14441# _0768_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5061 a_27295_4765# a_26431_4399# a_27038_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5063 a_14483_18543# _1075_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X5064 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5066 a_10310_2589# a_9871_2223# a_10225_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5067 a_8270_21237# a_8102_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5068 vccd1 _0835_.A1 a_4984_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5070 a_24278_11445# a_24110_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5072 vssd1 _0579_.C a_18213_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5073 vssd1 a_27590_14303# a_27548_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5074 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15023_28887# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5075 vssd1 _0440_.A _0445_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5076 a_14913_3311# a_14747_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5077 a_9945_2773# a_9779_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5079 a_9600_15823# _0935_.Q a_9003_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X5080 a_27422_15645# a_27149_15279# a_27337_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5081 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A _0819_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5082 _1008_.Q a_28015_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5083 a_7900_14165# _0768_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X5084 vssd1 _1078_.Q a_9503_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X5085 vssd1 _0935_.CLK a_8951_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5090 a_26007_10205# a_25309_9839# a_25750_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5091 vccd1 _0917_.CLK a_11435_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5092 a_20982_4765# a_20709_4399# a_20897_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5094 vssd1 _0836_.A _0836_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5095 vssd1 a_25842_15797# a_25800_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5097 a_2956_1956# a_2752_1897# a_3138_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0693 ps=0.75 w=0.42 l=0.15
X5099 a_8393_12015# _0684_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5100 a_22169_18365# _0928_.Q a_22097_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5101 vssd1 _0653_.A1 a_9135_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5102 a_8305_19407# _0761_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X5103 vccd1 fanout27.A a_23487_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X5104 a_10218_1679# a_9945_1685# a_10133_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5105 a_25214_8207# a_24941_8213# a_25129_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5106 a_10055_24527# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5107 a_12557_19407# _0864_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5109 a_12631_7663# _0522_.B1 a_12809_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5110 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE a_8215_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5111 a_20303_17821# a_19439_17455# a_20046_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5113 a_22825_8751# a_22659_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5114 vssd1 fanout13.A _0828_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5115 vccd1 a_17727_3855# a_17895_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5116 vccd1 _0582_.A a_19991_5056# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5117 vccd1 a_25842_10357# a_25769_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5119 a_22181_1685# a_22015_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5120 a_24757_16367# a_24591_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5121 vccd1 a_9411_15279# _0602_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5122 a_12711_14191# _0840_.A1 _0760_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5123 a_23792_13353# _0572_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5124 a_25589_21263# _0992_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5125 _0667_.B1 a_18001_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5126 _0524_.X a_11582_13077# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5127 vccd1 _0512_.X a_22373_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5128 a_4517_1501# a_3983_1135# a_4422_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5130 vssd1 a_1757_26703# _0832_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X5131 a_9217_14441# _0717_.A2 _0717_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5132 a_6779_2589# a_5915_2223# a_6522_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5133 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5134 a_13380_9673# a_12981_9301# a_13254_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R18 temp1.capload\[1\].cap_46.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5135 vssd1 a_9558_16885# a_9516_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5136 vssd1 _0505_.A2 a_21257_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5137 a_23193_9117# a_22659_8751# a_23098_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5138 vssd1 a_4847_1501# a_5015_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5139 vccd1 a_14453_14557# _0662_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X5140 a_14894_9951# a_14726_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5141 vssd1 a_14139_4943# a_14307_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5142 a_25723_23439# a_24941_23445# a_25639_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5143 a_5142_4511# a_4974_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5145 a_13616_30761# a_13367_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5146 vssd1 a_18539_11195# a_18497_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5147 vssd1 a_25547_13469# a_25715_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5151 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5152 a_23373_19465# a_22383_19093# a_23247_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5153 a_6805_12925# _0685_.B a_6733_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5154 vccd1 _0788_.C a_5913_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5155 vssd1 a_2623_6005# a_2581_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5156 a_17167_26525# a_16385_26159# a_17083_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5157 a_8929_2057# a_7939_1685# a_8803_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5158 a_14433_24501# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X5159 a_25401_7125# a_25235_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5160 a_27517_8029# a_26983_7663# a_27422_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5162 a_16101_18517# _0662_.A1 a_16354_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X5163 vccd1 a_18079_17723# a_17995_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5164 a_20341_5487# a_20175_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5165 a_12778_21237# a_12610_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5166 vssd1 _0745_.A2 a_5731_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5168 a_11509_15279# a_11343_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5169 a_13219_4765# a_12355_4399# a_12962_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5170 vssd1 a_26099_14735# a_26267_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5171 a_12705_1685# a_12539_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5176 _0489_.C1 a_23119_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5177 vssd1 a_24278_11445# a_24236_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5178 a_19697_6031# a_19163_6037# a_19602_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5179 a_2752_1897# clkbuf_1_0__f_io_in[0].X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5180 a_26099_19997# a_25235_19631# a_25842_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5181 vssd1 _0722_.B _0798_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5182 vccd1 a_14621_8897# _0614_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X5183 a_24017_18377# a_23027_18005# a_23891_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5184 a_8293_1679# _0674_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5185 vccd1 _0518_.Y a_16897_12897# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5187 vssd1 a_28015_16635# a_27973_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5188 _0515_.B1 a_13309_5515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X5189 vccd1 _1076_.Q a_14637_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X5190 vssd1 _0975_.CLK a_23947_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5191 vssd1 a_26267_4917# a_26225_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5192 _0529_.Y _0471_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5194 a_2885_2057# a_2752_1897# a_2464_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X5197 a_1639_7338# io_in[2] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5198 a_15929_14191# _1057_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5199 a_12981_9301# a_12815_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5200 a_8135_11249# _0699_.A0 a_7623_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X5201 vssd1 a_18447_3579# a_18405_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5203 a_12065_13647# _0917_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5204 a_17720_13353# _0658_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5206 _0838_.A0 _0472_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5207 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5209 vccd1 _1075_.Q a_11582_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X5210 a_12995_24527# _0444_.B a_12777_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5212 a_27590_3423# a_27422_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5213 vccd1 _0565_.A1 a_17260_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5215 a_21426_19743# a_21258_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5216 _0580_.C1 a_16127_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5217 a_14741_14013# a_14471_13647# a_14637_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5218 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5220 a_24462_22325# a_24294_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5221 vssd1 a_1775_15279# _0812_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5222 a_14444_28879# a_14195_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5223 a_22181_20181# a_22015_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5224 a_12276_6409# a_11877_6037# a_12150_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5225 vssd1 a_17083_26525# a_17251_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5226 a_25915_9117# a_25051_8751# a_25658_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5228 a_25405_17455# _0926_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5229 a_10643_4943# a_9779_4949# a_10386_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5230 _0549_.X a_16127_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5231 a_9857_11471# _0985_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5232 a_18942_25589# a_18774_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5233 a_10779_13103# _0768_.A1 _0714_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5234 a_9489_5487# _0549_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5235 vssd1 a_3819_26677# _1075_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5236 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5237 vccd1 a_21407_4765# a_21575_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5240 vssd1 _1062_.CLK a_23855_15831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5241 a_12632_8751# _0472_.X a_12526_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X5242 vssd1 _0847_.A3 a_10872_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5243 a_25677_3677# a_25143_3311# a_25582_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5246 vccd1 a_13679_9295# a_13847_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5249 vccd1 _0445_.A a_10789_22071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5250 a_10436_2223# a_10037_2223# a_10310_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5251 _0625_.A1 a_9339_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5253 _0475_.X a_11815_12265# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X5254 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5256 a_22917_7913# _1014_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5258 a_27149_12015# a_26983_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5260 vccd1 _0494_.X a_19439_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X5261 vccd1 a_12355_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5262 vccd1 a_28015_14459# a_27931_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5263 a_6833_13353# _0745_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5264 a_1975_29967# _0847_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X5266 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5268 vssd1 _0599_.X a_14621_8897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X5269 _0708_.A2 a_4447_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X5271 _0717_.A2 a_6467_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5272 vssd1 a_20671_8029# a_20839_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5273 a_18236_27247# temp1.dac.vdac_single.einvp_batch\[0\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5274 vccd1 a_20195_3829# a_20111_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5277 _0609_.C1 a_19439_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5279 a_16115_20495# _0860_.A _0863_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5280 a_27149_2223# a_26983_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5282 vccd1 a_20046_17567# a_19973_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5283 a_10041_22351# _1055_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5284 a_13177_2223# _0908_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5285 a_12069_2473# _0945_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X5286 _0907_.Q a_8327_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5287 a_4521_1679# _0905_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5288 a_9497_16367# a_9305_16672# _0880_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5291 a_10397_15823# _0836_.A a_10594_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5292 a_5510_8527# _0694_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X5293 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_13616_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5294 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5295 a_26927_21085# a_26063_20719# a_26670_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5296 a_25401_4949# a_25235_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5297 a_22015_13760# _0893_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5298 a_22917_7913# _0618_.B2 a_22833_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5299 a_17397_2767# a_16863_2773# a_17302_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5301 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5302 a_19593_12015# _0894_.Q a_19521_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5304 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5305 a_8105_1685# a_7939_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5306 a_3685_5321# a_2695_4949# a_3559_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5308 a_17538_13353# _0605_.D1 a_17289_13249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5309 vccd1 a_18371_1501# a_18539_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5310 vssd1 _0577_.C a_14441_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5311 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5312 vssd1 _0655_.X _0656_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X5314 a_16897_16395# _0521_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5315 a_7734_6031# a_7295_6037# a_7649_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5316 vssd1 _0577_.C a_17293_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5317 a_1941_4399# a_1775_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5318 a_19402_13621# a_19234_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5319 _0845_.B1 _0844_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5320 a_26597_21085# a_26063_20719# a_26502_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5321 vccd1 _0722_.A a_4167_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5322 a_2398_3677# a_1959_3311# a_2313_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5325 vssd1 a_8695_21237# a_8653_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5326 vccd1 _0602_.A a_22383_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5327 vssd1 fanout23.X a_27521_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5329 a_12342_1385# _0850_.Y _0854_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X5330 vccd1 a_10423_3855# _0959_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5332 _0544_.C a_13551_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X5334 _0675_.D a_11527_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X5336 a_2039_22057# _0753_.A2 io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5337 a_20437_21263# _0930_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5338 _0512_.A a_19439_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X5339 a_18601_5487# _0504_.A a_18519_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5340 temp1.capload\[6\].cap.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5341 vccd1 a_24462_1653# a_24389_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5342 vccd1 _0471_.X a_11435_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5344 a_25455_22173# a_24757_21807# a_25198_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5345 a_20717_1679# _0660_.X a_20635_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5346 vssd1 a_22622_16885# a_22580_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5347 a_4774_1653# a_4606_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5348 vccd1 a_26099_25615# a_26267_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5349 a_18048_14191# _0630_.A1 a_17473_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X5351 a_26835_11293# a_25971_10927# a_26578_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5352 a_26007_12381# a_25309_12015# a_25750_12127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5355 a_27249_11791# _0619_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5356 a_27847_5853# a_27149_5487# a_27590_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5357 vccd1 a_14710_20149# a_14637_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5358 a_10594_15823# a_10814_15797# _0529_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5359 a_4889_4399# input3.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5360 _0647_.B2 a_26267_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5361 a_13361_17455# a_13091_17455# a_13257_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5362 _0518_.Y a_7226_16885# a_7006_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5363 vssd1 a_26099_25615# a_26267_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5364 a_16998_6575# _1049_.Q a_16908_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X5366 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5367 a_19149_1679# _0645_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5368 a_22369_22351# _1017_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5369 a_11950_18655# a_11782_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5370 a_14603_18589# a_14287_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X5371 vssd1 _0722_.C a_5089_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5372 a_2030_9117# a_1757_8751# a_1945_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5373 a_21951_13469# a_21169_13103# a_21867_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5374 vssd1 a_26267_3829# a_26225_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5376 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_14444_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5377 a_1674_31599# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5378 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5379 a_10313_14735# _0770_.B2 a_10229_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5380 a_16565_14191# a_15575_14191# a_16439_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5381 a_2907_3677# a_2125_3311# a_2823_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5382 vccd1 a_12743_6005# a_12659_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5383 vssd1 a_6612_8181# _0710_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5384 vssd1 a_27847_22173# a_28015_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5385 vssd1 a_2991_2491# a_2949_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5386 a_15837_20719# _0920_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5388 vccd1 a_2566_2335# a_2493_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5389 a_5819_18793# _0795_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5390 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X5391 a_17302_3855# a_16863_3861# a_17217_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5392 a_5717_9615# _0710_.A1 _0711_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5393 vssd1 _0746_.A2 a_9583_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X5394 vccd1 _0686_.A a_6807_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5396 vccd1 a_10643_2767# a_10811_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5398 a_10714_20291# _0773_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X5399 vccd1 _1030_.CLK a_19163_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5400 a_13763_9295# a_12981_9301# a_13679_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5401 a_6613_22325# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X5402 vssd1 _0888_.CLK a_7295_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5403 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5404 vssd1 a_23415_1403# a_23373_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5405 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5406 _0488_.B2 a_24335_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5408 vccd1 fanout27.A a_15575_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5409 a_10083_12061# a_9791_12015# a_9997_12061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5410 a_23465_20719# a_22475_20719# a_23339_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5411 a_3651_26703# a_2787_26709# a_3394_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5412 vccd1 a_27463_4667# a_27379_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5413 a_25030_5853# a_24757_5487# a_24945_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5414 _1020_.Q a_22863_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5415 vccd1 a_27755_9117# a_27923_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5416 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5417 vssd1 a_10478_2335# a_10436_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5418 vssd1 a_22879_15823# a_23047_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5419 a_17351_22173# a_16569_21807# a_17267_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5420 vssd1 a_23361_13249# _0572_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X5421 a_12613_15829# a_12447_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5422 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X5423 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13360_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5424 a_12207_21085# a_11343_20719# a_11950_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5425 _0882_.Y a_11068_16617# a_11269_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5426 vccd1 _0483_.X a_22325_6603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5427 vccd1 a_21407_3677# a_21575_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5428 vccd1 _0745_.A3 a_6427_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X5430 a_4337_28335# _0847_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5431 a_5819_18793# _0782_.X a_5601_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5432 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X5433 vssd1 _0825_.S a_5541_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X5436 vccd1 _0655_.X a_7203_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5437 vssd1 a_4035_13077# _0780_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5439 a_18141_17999# _0667_.X a_18059_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5440 io_out[4] _0752_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5442 a_25777_1679# _1035_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X5443 a_8033_10703# _0679_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5444 vccd1 a_8031_16911# _0836_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5445 _0921_.Q a_13479_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5446 a_10727_2767# a_9945_2773# a_10643_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5447 vccd1 a_16897_12897# _0533_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X5448 a_17486_17821# a_17047_17455# a_17401_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5449 a_20414_14709# a_20246_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5450 a_9574_5853# a_9135_5487# a_9489_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5451 _0807_.B a_9043_12567# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5452 vccd1 a_10386_1653# a_10313_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5453 a_26410_11293# a_26137_10927# a_26325_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5454 a_21081_27247# _1019_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5455 a_16592_18543# _0667_.B1 a_16101_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5456 vccd1 a_25382_8181# a_25309_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5457 a_1945_6575# _0877_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5458 vccd1 _0630_.X a_15921_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X5460 vccd1 a_21851_19899# a_21767_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5461 vccd1 _1077_.Q a_8859_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5462 vssd1 _0717_.A2 a_8101_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X5463 a_12291_15645# a_11509_15279# a_12207_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5464 a_17761_2223# _0956_.Q a_17323_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5465 _0621_.A1 a_25623_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5467 a_20027_3855# a_19329_3861# a_19770_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5468 a_5299_2767# a_4517_2773# a_5215_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5469 _0512_.A a_19439_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5470 vssd1 _0583_.C a_19041_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5471 a_22606_15529# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5472 vssd1 a_11760_26935# _0823_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5473 vssd1 _0789_.B1 a_6611_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X5474 a_26099_25615# a_25235_25621# a_25842_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5475 vssd1 a_5549_17719# _0797_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X5476 a_20246_14735# a_19973_14741# a_20161_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5478 a_17670_23261# a_17231_22895# a_17585_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5479 a_21518_18655# a_21350_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5481 vccd1 a_25455_15645# a_25623_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5482 vccd1 a_6947_2491# a_6863_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5483 vccd1 a_4036_30663# _0798_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5484 _1067_.Q a_26267_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5485 vssd1 _0456_.B _0722_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X5486 vccd1 a_2823_1501# a_2991_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5487 _0872_.A1 a_4386_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X5488 vssd1 a_21775_18909# a_21943_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5489 a_5793_16367# _0873_.A a_5721_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5491 vssd1 a_21407_4765# a_21575_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5492 vssd1 _0745_.A2 _0756_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5494 a_11269_16367# _0882_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5495 vssd1 a_1591_14191# _0456_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5498 a_22549_14191# a_22383_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5499 a_6522_2335# a_6354_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5500 vssd1 a_25842_25589# a_25800_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5501 a_25401_3861# a_25235_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5504 a_12337_21269# a_12171_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5505 a_7860_6409# a_7461_6037# a_7734_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5506 vssd1 _0505_.A2 a_23005_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5507 vccd1 fanout13.A a_15667_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X5509 _0893_.Q a_28015_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5510 a_2524_3311# a_2125_3311# a_2398_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5511 vccd1 _0842_.A0 a_11711_1792# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5512 _0908_.Q a_8235_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5513 _0763_.A2 a_7663_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5514 a_22974_18793# _0994_.D a_22817_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5517 vccd1 a_13387_4667# a_13303_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5518 a_4253_9839# _0807_.B a_4035_9813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5520 a_22837_10927# _0926_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5521 vccd1 a_27847_10205# a_28015_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5522 a_14637_13647# a_14471_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X5524 _0597_.A1_N a_15759_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X5525 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5526 a_8653_21641# a_7663_21269# a_8527_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5528 a_24867_17999# _0662_.B1 a_24949_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5530 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10140_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5533 a_1639_7828# io_in[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5534 a_2493_2589# a_1959_2223# a_2398_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5535 vssd1 _0502_.X a_22169_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5538 vssd1 a_25198_16479# a_25156_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5540 vccd1 _0888_.CLK a_8307_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5542 a_14726_10205# a_14453_9839# a_14641_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5543 vccd1 a_15703_2589# a_15871_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5544 _0882_.Y a_11068_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5545 vccd1 a_15795_1679# a_15963_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5546 a_23745_21263# a_23211_21269# a_23650_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5547 a_17092_18319# _0577_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X5548 a_23557_7497# a_22567_7125# a_23431_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5549 vssd1 _0816_.S a_6416_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5552 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_12316_24135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5553 a_8105_18793# _0719_.B2 a_8021_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5554 a_13395_15823# a_12613_15829# a_13311_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5555 vccd1 _0662_.B1 a_25225_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5556 a_5399_4765# a_4535_4399# a_5142_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5557 vssd1 a_5659_4917# a_5617_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5561 vccd1 a_27279_18811# a_27195_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5562 vccd1 a_15319_7931# a_15235_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5563 _0585_.X a_19439_12675# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5564 a_2490_28701# a_2051_28335# a_2405_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5565 a_17428_4233# a_17029_3861# a_17302_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5566 a_18313_6409# a_17323_6037# a_18187_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5567 temp1.capload\[10\].cap.Y temp1.capload\[10\].cap.A a_8301_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5568 vccd1 a_12356_19203# _0865_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5569 a_17904_14441# _0630_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5570 _0860_.A a_2114_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5571 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5572 _0548_.B2 a_23139_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5573 vccd1 a_12042_9951# a_11969_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5574 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_9135_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5575 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_6368_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5576 vssd1 a_11950_18655# a_11908_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5577 vccd1 a_10811_4917# a_10727_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5578 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5580 a_10140_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5581 a_22879_1679# a_22015_1685# a_22622_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5582 a_4769_23145# _0742_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5583 a_17428_10761# a_17029_10389# a_17302_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5585 a_17378_19743# a_17210_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5587 a_6600_11587# _0745_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5589 a_26183_19087# a_25401_19093# a_26099_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5591 a_10313_1679# a_9779_1685# a_10218_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5592 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5593 vssd1 _1019_.CLK a_21003_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5594 vssd1 _0828_.Y a_12176_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5595 vssd1 a_17635_19997# a_17803_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5596 vssd1 a_16439_14557# a_16607_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5597 temp1.capload\[12\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5598 vssd1 a_7625_14709# _0793_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5599 a_14300_19465# a_13901_19093# a_14174_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5600 _1064_.Q a_27003_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5601 vccd1 _0827_.A a_7469_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5602 vccd1 a_2991_27515# a_2907_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5603 a_8159_6031# a_7461_6037# a_7902_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5604 vccd1 a_2198_8863# a_2125_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5605 _0572_.D1 a_23303_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5606 vssd1 a_2623_5755# a_2581_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5608 a_22825_11177# _0506_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5609 vccd1 a_21667_20987# a_21583_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5610 a_11067_19631# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X5611 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11704_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5614 vccd1 _0840_.A0 a_9600_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X5615 vccd1 a_11435_8751# _0842_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5617 vssd1 _0460_.C a_1867_15831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5619 vssd1 _0524_.X a_18213_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5620 a_12276_11849# a_11877_11477# a_12150_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5621 vssd1 a_22622_1653# a_22580_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5622 a_9700_5487# a_9301_5487# a_9574_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5623 a_26041_8751# a_25051_8751# a_25915_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5624 vccd1 _0707_.A1 a_6001_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X5626 vccd1 a_18279_3677# a_18447_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5627 vssd1 a_2715_3829# a_2673_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5628 _0532_.A2 a_12479_5515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5629 vssd1 a_4831_3829# a_4789_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5630 _0651_.X a_22199_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5633 a_9312_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5634 a_4590_26271# a_4422_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5635 vssd1 a_23339_21085# a_23507_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5636 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_11711_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5637 a_17029_3861# a_16863_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5638 vccd1 a_2626_9269# _0835_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5639 a_25455_16733# a_24591_16367# a_25198_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5640 a_9919_6740# _0854_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5641 vssd1 a_4847_26525# a_5015_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5642 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10324_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5643 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5646 vssd1 a_9613_25045# a_9547_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5647 a_15741_4399# a_15575_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5648 vssd1 _0999_.CLK a_23211_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5649 a_27149_7663# a_26983_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5651 vssd1 _0845_.C1 _0839_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5652 _0860_.A a_2114_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X5654 vccd1 a_25198_5599# a_25125_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5656 a_11509_15279# a_11343_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5657 vccd1 fanout24.A a_25235_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5658 a_22963_15823# a_22181_15829# a_22879_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5659 _0674_.A1 a_9615_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5660 a_24757_2223# a_24591_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5662 vssd1 a_25842_7093# a_25800_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5663 a_6563_12015# _0745_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X5665 vssd1 a_20782_5599# a_20740_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5666 a_20801_20719# a_20635_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5667 _0517_.B a_19439_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X5668 vssd1 _1015_.CLK a_26983_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5669 vssd1 a_2566_3423# a_2524_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5670 a_4793_4949# a_4627_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5671 a_19846_9295# _0590_.B2 a_19689_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5672 a_21334_27359# a_21166_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5673 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_6559_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5674 a_6639_17455# _0873_.A _0749_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5676 vccd1 _0995_.CLK a_8307_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5677 vssd1 a_25382_23413# a_25340_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5678 vccd1 a_24059_17973# a_23975_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5679 a_25589_4943# _0531_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5680 vccd1 a_20977_10901# _0496_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5681 vssd1 _0778_.A2 a_6805_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5682 vssd1 a_7389_25335# _0825_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
R19 temp1.capload\[3\].cap_48.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5684 a_23193_18005# a_23027_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5686 _1013_.Q a_28015_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5687 vccd1 _0917_.CLK a_12815_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5688 a_23891_26703# a_23027_26709# a_23634_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5690 a_1775_28879# _0845_.A2 _0836_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5691 vccd1 a_23818_21237# a_23745_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5693 a_14655_11177# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5694 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5696 a_7203_10089# _0685_.B a_7457_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5697 _0850_.Y _0847_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5698 _0621_.A1 a_25623_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5699 a_18025_7809# _0634_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5700 a_13472_10761# a_13073_10389# a_13346_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5702 a_25769_1501# a_25235_1135# a_25674_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5703 a_1757_9301# a_1591_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5704 a_26053_13967# _0928_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5705 a_9669_1501# a_9135_1135# a_9574_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5710 a_9815_16911# a_9117_16917# a_9558_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5712 vccd1 a_17289_13249# _0605_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X5714 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5715 a_23561_26703# a_23027_26709# a_23466_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5716 a_21242_20831# a_21074_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5718 vccd1 _0814_.A2 a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5719 vccd1 a_12759_3855# a_12927_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5720 vccd1 _0504_.A a_15667_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5721 a_17486_17821# a_17213_17455# a_17401_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5722 _0722_.B _0456_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5723 a_22373_16617# _1019_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X5724 vccd1 _0505_.A2 a_17497_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
D2 vssd1 _0858_.X sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X5726 a_26210_26271# a_26042_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5727 a_7843_14735# _0461_.A a_7625_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5728 vssd1 a_8546_4917# a_8504_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5729 vccd1 a_4864_11445# _0745_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X5730 _0835_.Y _0835_.A1 a_5177_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5731 vssd1 a_19689_9269# _0590_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X5732 a_27149_12015# a_26983_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5733 a_4547_25393# _0842_.A0 a_4035_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X5735 vssd1 _0659_.X a_21831_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5736 vssd1 a_6151_21781# _0809_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5737 a_3965_3861# a_3799_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5738 a_1849_3861# a_1683_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5739 a_27146_6941# a_26873_6575# a_27061_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5742 a_18282_18793# _0932_.Q a_18125_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5743 a_2125_9117# a_1591_8751# a_2030_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5744 _0696_.A1 _0734_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5745 _0678_.Y _0472_.X a_8485_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5746 vccd1 a_12375_18811# a_12291_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5747 a_19149_13647# _1025_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5748 vccd1 _0847_.A2 a_6559_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5750 a_19697_11471# _1057_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5751 a_14195_11471# _0474_.X _0630_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5752 _0675_.C a_16863_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5754 vssd1 _0845_.C1 _1078_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5756 a_21345_15253# _0558_.A2 a_21502_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5757 vccd1 fanout23.X a_26431_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5758 a_20855_22351# a_19991_22357# a_20598_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5759 a_20901_16617# _0564_.D a_20819_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
R20 temp1.capload\[8\].cap_53.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5760 vssd1 _0831_.D a_2033_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X5761 vccd1 fanout23.X a_25235_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5762 vccd1 _0908_.CLK a_9135_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5764 a_14287_14557# _0511_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5765 vssd1 a_2823_27613# a_2991_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5766 a_2975_17461# _0456_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5767 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5768 a_13629_4943# _0670_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5770 a_11747_3677# a_10883_3311# a_11490_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5771 a_22822_3677# a_22383_3311# a_22737_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5772 a_25125_5853# a_24591_5487# a_25030_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5773 vssd1 _0572_.A2 a_21625_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5774 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_3983_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5775 a_9895_10089# _0545_.B2 a_10089_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X5776 a_15753_7235# a_15565_7235# a_15671_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X5777 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_15667_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5778 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5779 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5780 a_7283_20719# _0845_.A1 _0869_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5781 _0819_.S _0837_.A1 a_10142_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5782 _1059_.D a_16607_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5783 a_17473_14337# _0627_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5785 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5786 vccd1 a_5031_1679# a_5199_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5787 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI a_14188_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5788 _0998_.D a_26911_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5790 vssd1 _0864_.Y a_12557_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5791 a_26835_11293# a_26137_10927# a_26578_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5792 a_12219_26742# _0825_.A0 a_11760_26935# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X5793 _0828_.Y fanout13.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5795 vssd1 _0872_.A1 a_3327_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X5796 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5797 vssd1 a_18371_1501# a_18539_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5798 a_6151_21781# _0764_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X5799 _0813_.A2 a_4132_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5800 vssd1 fanout24.A a_22015_8215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5801 _0602_.A a_9411_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5803 vccd1 _1053_.CLK a_14471_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5804 _0511_.D a_9963_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5805 a_18677_2473# _0591_.X a_18605_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5808 a_11895_1135# _0835_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X5809 vssd1 _0542_.X a_14839_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5810 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X5811 vccd1 _0908_.CLK a_5915_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5812 vccd1 a_27590_9951# a_27517_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5813 a_20111_10955# _0602_.A a_20025_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5814 a_5466_22895# _0788_.C a_4403_22869# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.08775 ps=0.92 w=0.65 l=0.15
X5815 vssd1 a_15151_8029# a_15319_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5816 vccd1 _0512_.X a_19429_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5817 vssd1 _0529_.Y a_19593_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5818 _0444_.B a_11803_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X5820 a_27130_13215# a_26962_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5821 a_4160_32463# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5822 a_19281_18337# _0512_.A a_19195_18337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5823 a_16945_7119# _0487_.X a_17029_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5824 _1080_.Q a_3083_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5825 a_20801_20719# a_20635_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5826 a_18317_20181# a_18151_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5827 vccd1 _0975_.CLK a_22107_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5829 vccd1 a_21943_18811# a_21859_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5830 a_14905_17277# _0511_.D a_14833_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X5832 vssd1 _0995_.CLK a_8307_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5834 a_25589_15823# _0892_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5835 vccd1 _1033_.CLK a_25051_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5836 a_10876_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5837 a_27422_2589# a_27149_2223# a_27337_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5843 vssd1 _0491_.X a_19877_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X5844 a_13349_9295# a_12815_9301# a_13254_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5845 a_18298_11445# a_18130_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5846 vccd1 a_23634_26677# a_23561_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5847 a_14839_5487# _0645_.B1 a_15017_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5848 _0837_.Y _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5849 _0814_.A2 a_3891_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5850 a_10033_19631# _0798_.A2 a_9687_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5851 _0674_.C1 a_11987_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5852 a_25309_23439# a_24775_23445# a_25214_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5853 vccd1 _0814_.A2 _0752_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5854 a_25999_8029# a_25217_7663# a_25915_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5855 a_15115_13103# _1076_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5857 a_12843_3855# a_12061_3861# a_12759_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5858 a_1766_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5859 io_out[2] _0444_.A a_1591_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5860 a_12207_21085# a_11509_20719# a_11950_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5861 a_6728_15529# _0758_.B1 a_6473_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5864 a_25582_10205# a_25143_9839# a_25497_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5865 a_1775_27791# _0843_.B _0843_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5866 vssd1 _0722_.B a_4132_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X5867 a_10862_11293# a_10423_10927# a_10777_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5868 _0954_.D a_10811_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5869 _0676_.B a_15391_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5870 a_22695_26525# a_21997_26159# a_22438_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5871 a_12701_14025# a_11711_13653# a_12575_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5872 vssd1 _0494_.X a_18731_7457# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X5873 vccd1 a_23047_20149# a_22963_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5874 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X5875 vssd1 _1019_.CLK a_19991_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5876 a_9305_16911# _0986_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5878 vssd1 _0572_.X a_19439_12675# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5879 a_13433_17455# _1075_.Q a_13361_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X5880 vssd1 a_8803_4943# a_8971_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5882 vssd1 _0753_.A2 a_1591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
X5883 a_27548_16367# a_27149_16367# a_27422_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5884 vccd1 a_5567_4667# a_5483_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5885 a_5915_13103# _0791_.A2 a_5821_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5888 a_9531_3855# a_8749_3861# a_9447_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5889 _0791_.A1 _0745_.A1 a_3333_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5891 a_25474_6687# a_25306_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5893 vssd1 a_19659_1679# a_19827_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5895 vccd1 a_13403_1679# a_13571_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5896 a_2539_9295# a_1757_9301# a_2455_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X5897 a_16090_20831# a_15922_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5899 _0863_.Y _0863_.A2 a_15945_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5901 a_23742_6031# a_23469_6037# a_23657_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5902 a_8325_11769# _0466_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5903 a_17865_9845# _0624_.D_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5904 a_11582_13077# _1076_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5905 a_25474_6687# a_25306_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5910 _0816_.S _0835_.A1 a_9774_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5911 a_8176_19061# _0813_.A2 a_8399_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5912 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5913 _0835_.A1 a_2626_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X5914 vssd1 _0710_.B2 a_4451_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5916 a_10714_20541# _0773_.A2_N a_10714_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X5917 a_23247_3677# a_22383_3311# a_22990_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5919 a_27847_24349# a_27149_23983# a_27590_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5920 vssd1 _0999_.CLK a_22015_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5921 a_9786_26486# _0819_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5923 a_4517_2773# a_4351_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5924 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5925 a_11149_14441# _0747_.B1 a_11233_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5926 a_13035_21263# a_12337_21269# a_12778_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5928 _0937_.Q a_14767_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5929 vssd1 _0487_.X a_15380_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X5932 vccd1 fanout37.A a_4259_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X5934 vccd1 ANTENNA_7.DIODE a_4811_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5935 a_25401_10389# a_25235_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5937 a_2455_6941# a_1757_6575# a_2198_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5938 vssd1 a_27590_25183# a_27548_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5939 a_17857_11477# a_17691_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5940 a_10120_31849# a_9871_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5943 vccd1 _0444_.A a_2419_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5944 vssd1 a_12743_6005# a_12701_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5945 a_22948_3311# a_22549_3311# a_22822_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5946 a_19846_9295# _0582_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X5948 vssd1 fanout37.A a_23763_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X5949 vccd1 a_2915_25437# a_3083_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5950 _0631_.B a_22311_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5951 _0572_.A1 a_26267_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5952 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5953 a_7025_18865# _0761_.B a_6516_18695# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X5954 vccd1 _0931_.CLK a_18151_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5955 a_24293_9673# a_23303_9301# a_24167_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5956 a_22737_19087# _1016_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5957 a_24945_4399# _0548_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5959 a_9786_26159# _0819_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X5960 _1054_.Q a_15595_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5961 vssd1 a_3270_2741# _0850_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X5962 vssd1 _0988_.D a_16592_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5963 _0669_.X a_21279_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5964 vccd1 a_25842_21237# a_25769_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5965 _0695_.A1 _0656_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5966 _0645_.B1 a_15793_6603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X5967 a_2765_4399# a_1775_4399# a_2639_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5968 _1068_.Q a_27279_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5969 _0518_.Y _0472_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5971 a_22369_1679# _0618_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5972 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5973 vccd1 clkbuf_0__0390_.A a_4802_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5974 vccd1 a_21683_19997# a_21851_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5975 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_12532_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5976 vccd1 a_9184_25223# _0817_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5977 temp1.capload\[1\].cap.Y temp1.capload\[1\].cap_46.LO a_4529_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5978 vssd1 a_7256_17429# _0719_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5979 a_27337_17455# _0927_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5981 a_10789_22071# _0441_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X5983 a_23637_12533# _0576_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5984 a_27973_7663# a_26983_7663# a_27847_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5986 vssd1 _0872_.A1 a_5793_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5987 vccd1 _0521_.A a_22015_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5989 vccd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_1766_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5990 vccd1 _0602_.A a_17783_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5991 a_21361_6825# _0669_.B2 a_21279_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5993 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11152_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X5994 vssd1 _0658_.B1 a_19969_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X5997 vccd1 a_15538_1653# a_15465_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5998 a_18961_13653# a_18795_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5999 a_14668_20553# a_14269_20181# a_14542_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6000 a_25589_7119# _0573_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6002 vssd1 a_23783_8181# a_23741_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6003 _0985_.D a_13939_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6004 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6005 a_27590_21919# a_27422_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6006 a_22741_11791# _0992_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6007 vccd1 a_7348_17973# _0742_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X6008 _0604_.B a_10811_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6009 _0505_.A1 a_25807_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6010 vssd1 _0776_.A2 _0745_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6011 vccd1 a_24703_11445# a_24619_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6012 a_2313_3311# _0868_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6013 _0920_.Q a_16515_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6014 vssd1 a_17473_14337# _0630_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X6015 _0513_.X a_9911_12061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X6016 vccd1 a_8803_1679# a_8971_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6017 a_12978_1679# a_12705_1685# a_12893_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6018 vssd1 _0836_.A _0518_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6019 a_25708_9839# a_25309_9839# a_25582_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6020 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6021 a_5031_1679# a_4167_1685# a_4774_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6022 a_8004_27791# a_7755_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6023 vssd1 _0825_.A0 _0815_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6024 vssd1 _0515_.B1 a_16105_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6025 a_26318_23261# a_26045_22895# a_26233_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6026 a_25842_7093# a_25674_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6027 a_1674_31599# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X6029 a_22015_6144# _0575_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6030 a_17618_13353# _0605_.C1 a_17538_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X6031 _0664_.X a_25971_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6033 vccd1 _0873_.A a_3241_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X6034 vssd1 a_15319_12283# a_15277_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6035 vccd1 a_11803_23439# _0444_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X6036 a_18758_20149# a_18590_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6037 a_19439_9839# _0630_.A2 a_19617_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6038 vssd1 a_3523_6039# fanout37.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6039 _0868_.A2 a_7244_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6041 a_4771_12791# _0758_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6042 a_26183_10383# a_25401_10389# a_26099_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6043 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6044 _0608_.X a_20083_15936# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6045 vssd1 a_5215_2767# a_5383_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6046 a_18639_11471# a_17857_11477# a_18555_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6047 a_21867_13469# a_21003_13103# a_21610_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6049 vccd1 _0511_.D a_13257_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X6050 vccd1 a_27314_6687# a_27241_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6052 a_9644_26311# _0825_.A0 a_9786_26486# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6053 a_10229_14735# _0812_.A2 a_10147_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6054 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6055 a_25581_2223# a_24591_2223# a_25455_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6056 a_14464_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6057 a_4149_2223# a_3983_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6058 _0621_.X a_23303_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6059 _0768_.A1 a_3523_13655# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6060 a_8392_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6061 a_17397_22895# a_17231_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6062 vssd1 _0995_.CLK a_15667_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6063 a_7557_4399# _0907_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6065 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X6067 a_5621_6575# _0698_.B1 a_5537_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6068 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10120_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6069 a_21537_13469# a_21003_13103# a_21442_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6070 vssd1 _0827_.A temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6073 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6074 a_22369_16911# _1062_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6075 a_12334_3855# a_11895_3861# a_12249_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6076 a_12610_21807# a_12433_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6077 a_8293_4943# _0538_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6079 vssd1 clkbuf_1_0__f_io_in[0].X a_3983_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6081 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6082 vccd1 _0999_.CLK a_22383_19093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6083 a_14910_17999# a_14637_18005# a_14825_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6084 _0921_.Q a_13479_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6085 a_19613_16617# _0561_.C1 a_19531_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6086 vccd1 a_4221_8725# _0699_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6089 a_17267_22173# a_16403_21807# a_17010_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6090 a_26686_18909# a_26413_18543# a_26601_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6091 vccd1 a_11455_11195# a_11371_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6092 vccd1 _0935_.CLK a_12447_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6093 vssd1 a_26267_10357# a_26225_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6094 vssd1 a_6651_28335# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6095 vssd1 a_18723_11445# a_18681_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6097 vccd1 a_28015_25339# a_27931_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6098 vccd1 a_11915_3579# a_11831_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6100 vssd1 _0717_.B1 a_7256_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X6101 a_25769_14735# a_25235_14741# a_25674_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6102 vssd1 _0646_.C1 a_12631_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6103 a_25490_17821# a_25051_17455# a_25405_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6105 vssd1 _0670_.A2 a_14920_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6106 vssd1 _0662_.A3 a_16981_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6108 vccd1 _0791_.A3 a_5074_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X6110 _0850_.Y _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6111 vccd1 a_2787_7119# _0888_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6113 vccd1 a_17083_26525# a_17251_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6114 a_9492_18543# _0840_.A1 a_9189_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X6115 a_27422_5853# a_26983_5487# a_27337_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6117 vccd1 a_13311_15823# a_13479_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6118 a_11490_3423# a_11322_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6119 a_25382_8181# a_25214_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6120 a_25225_14441# _0996_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6123 _0474_.X a_10147_15529# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X6126 vccd1 _0441_.B a_11435_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6127 vccd1 a_2381_16885# _0875_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6129 vccd1 a_12316_24135# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6130 a_12207_15645# a_11343_15279# a_11950_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6131 a_1757_8751# a_1591_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6132 vssd1 a_12189_27001# a_12123_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6133 a_9003_15797# _0508_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6135 a_23098_4765# a_22825_4399# a_23013_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6136 _0601_.B1 a_14655_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6137 a_4414_30511# _0798_.A1 a_4036_30663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X6138 vssd1 _0888_.CLK a_7939_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6139 a_13432_25615# a_13183_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6142 a_15465_1679# a_14931_1685# a_15370_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6143 a_22270_26525# a_21997_26159# a_22185_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6144 vssd1 ANTENNA_7.DIODE a_3799_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6146 _0624_.C a_22751_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X6147 _0797_.A1 a_5549_17719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X6148 a_25455_15645# a_24757_15279# a_25198_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6149 vccd1 _0466_.A _0546_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6150 a_21491_4765# a_20709_4399# a_21407_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6151 a_8102_21263# a_7663_21269# a_8017_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6153 vccd1 a_26099_19087# a_26267_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6154 _0919_.D a_12375_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6155 vccd1 _0917_.CLK a_11711_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6156 vccd1 a_21150_3423# a_21077_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6158 a_20697_9839# _1025_.Q a_20625_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6159 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_14195_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6161 vssd1 _0882_.A2 a_11269_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6162 vccd1 a_6704_13077# _0747_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X6163 a_4324_20291# _0722_.B a_4252_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6164 _0456_.B a_1591_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6166 a_4606_1679# a_4167_1685# a_4521_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6167 vssd1 _0831_.D a_10055_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6168 a_6813_19087# _0440_.C _0445_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6169 a_8378_1679# a_8105_1685# a_8293_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6170 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_11746_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6171 a_27590_15391# a_27422_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6172 _0749_.B1 a_11067_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X6173 a_26873_6575# a_26707_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6176 vccd1 a_19367_25589# a_19283_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6178 a_18141_17999# _0584_.A2 a_18225_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6179 vccd1 _0964_.CLK a_26983_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6181 vssd1 _1028_.CLK a_12355_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6183 vssd1 a_27847_15645# a_28015_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6184 vccd1 a_27590_2335# a_27517_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6185 vssd1 _0648_.A2 a_19969_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X6186 _0842_.A0 a_11435_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6187 a_11789_9839# _0625_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6188 a_10198_7351# _0565_.X a_10412_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6189 a_17128_15279# _0580_.A1 a_16553_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X6190 a_4537_10927# a_4251_11249# a_4040_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6191 _0843_.B a_4035_25045# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6192 a_23266_8863# a_23098_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6193 a_27167_10383# _0619_.B1 a_27249_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6194 vccd1 fanout10.A a_10975_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6195 a_23634_17973# a_23466_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6196 a_2382_4511# a_2214_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6197 a_27241_6941# a_26707_6575# a_27146_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6198 _0920_.D a_15135_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6199 vccd1 _0464_.X a_3523_13655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6200 _0850_.A a_3270_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X6201 _0694_.A2 _0689_.X a_6463_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6202 vssd1 a_25750_9951# a_25708_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6203 a_21039_5853# a_20175_5487# a_20782_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6204 a_11030_11039# a_10862_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6206 vccd1 a_22622_22325# a_22549_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6207 a_8325_11769# _0466_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6208 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6209 a_24209_20175# _0965_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6211 a_20246_14735# a_19807_14741# a_20161_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6212 vssd1 _0535_.X a_13069_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6213 a_21951_24349# a_21169_23983# a_21867_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6214 a_2290_3829# a_2122_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6215 a_27590_7775# a_27422_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6216 a_8485_13103# _0546_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6219 a_23466_17999# a_23193_18005# a_23381_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6220 a_16209_7913# _0644_.A2 a_16293_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6222 a_18597_21263# _1060_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6223 a_3983_31849# _0814_.B1 a_4065_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6224 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6226 vssd1 a_8123_13647# _0778_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X6227 a_6416_24233# _0764_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6228 a_6938_14237# _0717_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X6229 a_9945_4949# a_9779_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6230 a_5325_8181# _0710_.A2 a_5829_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6231 vssd1 fanout23.X a_25235_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6232 vccd1 _0888_.CLK a_4535_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6233 vssd1 _0908_.CLK a_9135_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6234 vccd1 a_23910_6005# a_23837_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6235 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_7295_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6237 a_13735_3968# _0639_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6238 a_22714_2741# a_22546_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6240 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6241 a_20430_20175# a_19991_20181# a_20345_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6242 vssd1 a_19439_14191# _1062_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6243 vssd1 a_2626_9269# a_2584_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X6244 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_7939_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6245 vccd1 _0630_.A1 a_17904_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6246 a_15671_7235# _0634_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6247 vssd1 _0438_.A a_9043_12567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6248 vccd1 a_23415_3579# a_23331_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6252 vssd1 _0850_.A a_8256_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6255 a_4149_1135# a_3983_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6256 _1026_.Q a_19827_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6257 a_27149_16367# a_26983_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6258 a_12460_4233# a_12061_3861# a_12334_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6259 _0639_.X a_13735_3968# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6262 a_26743_23261# a_26045_22895# a_26486_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6263 a_22606_15529# _0927_.D a_22449_15253# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6264 vccd1 a_2455_5853# a_2623_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6265 _0801_.X a_14319_20747# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6266 vssd1 fanout37.A a_9227_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6267 a_22990_3423# a_22822_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6268 vccd1 a_23763_10927# _1015_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6270 vccd1 _0662_.A3 a_14655_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6271 vssd1 fanout24.A a_27202_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6273 _1026_.Q a_19827_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6274 a_1975_30287# _0847_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6275 vccd1 a_5199_1653# a_5115_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6276 a_4342_30761# _0814_.A2 a_4036_30663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6277 a_15016_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6278 a_26099_19087# a_25235_19093# a_25842_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6279 vssd1 a_22015_3855# _0975_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6281 a_2869_17501# _0722_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6282 vssd1 a_15667_2767# _0972_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6284 a_16565_4399# a_15575_4399# a_16439_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6285 vccd1 _0803_.X a_5264_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X6286 a_15737_15113# a_14747_14741# a_15611_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6287 vssd1 a_2823_2589# a_2991_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6289 a_15844_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6290 vssd1 _0805_.A a_4386_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6291 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6292 a_19605_4649# _0497_.B2 a_19521_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6293 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9312_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6294 a_17217_10383# _0983_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6295 vccd1 a_26083_7931# a_25999_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6296 vccd1 _0466_.A _0684_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X6297 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6298 a_22917_1501# a_22383_1135# a_22822_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6299 a_11782_18909# a_11509_18543# a_11697_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6300 a_27548_5487# a_27149_5487# a_27422_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6303 a_20027_26703# a_19163_26709# a_19770_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6304 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13432_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6305 _0723_.X a_6416_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6306 a_4406_3829# a_4238_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6307 a_2290_3829# a_2122_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6308 vccd1 a_21591_27613# a_21759_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6309 a_25198_2335# a_25030_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6310 vssd1 a_4259_6031# _0922_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6311 vccd1 _0523_.X a_14261_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X6312 fanout27.A a_16863_11479# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6314 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6315 vssd1 a_23247_1501# a_23415_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6317 _1020_.Q a_22863_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6318 a_15051_20175# a_14269_20181# a_14967_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6319 a_21825_7663# _0967_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6320 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6321 a_15971_16733# a_15189_16367# a_15887_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6322 a_22281_10499# _0650_.X a_22199_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6323 a_4422_28701# a_3983_28335# a_4337_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6325 vssd1 a_25382_8181# a_25340_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6326 vssd1 _0563_.C1 a_22291_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6327 vccd1 a_15795_27791# a_15963_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6328 vccd1 _1023_.Q a_19202_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6329 _0702_.B1_N a_4852_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6331 a_19697_26703# a_19163_26709# a_19602_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6335 vccd1 _0863_.A1 a_15945_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6336 _0866_.B a_13367_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6337 a_9926_9269# a_9758_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6340 vssd1 fanout10.A a_11803_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6341 a_4590_1247# a_4422_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6342 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6343 a_3134_4943# a_2861_4949# a_3049_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6344 a_15002_3855# a_14729_3861# a_14917_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6345 vccd1 a_26007_12381# a_26175_12283# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6346 a_11251_5737# _0667_.B1 a_11333_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6347 _0633_.X a_20543_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6348 a_22879_15823# a_22015_15829# a_22622_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6354 a_15661_31599# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6355 a_4732_2057# a_4333_1685# a_4606_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6356 vssd1 _0931_.CLK a_20635_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6357 a_8159_6031# a_7295_6037# a_7902_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6358 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10948_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6362 a_20393_8545# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6363 vssd1 clkbuf_1_1__f_net57.A a_1674_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6364 _0805_.A a_4843_19659# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6365 vccd1 _1078_.Q a_14287_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6366 a_25674_3855# a_25401_3861# a_25589_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6367 a_5325_8181# _0734_.A2 a_5612_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X6368 vccd1 a_18022_3423# a_17949_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6369 vccd1 a_4811_10383# _0845_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6370 _0556_.B a_17323_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6372 a_13472_22729# a_13073_22357# a_13346_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6373 a_22549_15823# a_22015_15829# a_22454_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6375 _0930_.Q a_25623_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6376 a_6283_20719# _0869_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6378 a_27590_14303# a_27422_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6379 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6380 a_14729_16911# a_14563_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X6382 vssd1 _0827_.A fanout9.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6383 _0825_.A1 a_7389_25335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X6384 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6385 vssd1 _0964_.CLK a_23027_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6388 a_15312_15113# a_14913_14741# a_15186_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6389 vssd1 a_27847_14557# a_28015_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6391 a_7900_14165# _0768_.A1 a_8120_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6392 vccd1 _0931_.CLK a_20819_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6393 vssd1 _0652_.C _0684_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6395 _0710_.B2 a_5128_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6397 a_19743_1679# a_18961_1685# a_19659_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6398 vssd1 _0643_.B1 a_25581_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X6399 vssd1 _0523_.B1 a_17117_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6400 vssd1 _0847_.A2 _0788_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6401 a_7457_10089# _0685_.B a_7203_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6403 vccd1 _0798_.A2 _0814_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6405 vccd1 _0708_.A2 a_4993_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X6406 _0739_.A2 a_6559_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X6407 vccd1 a_20839_14709# a_20755_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6408 _0625_.A1 a_9339_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6410 a_10007_26159# _0825_.A0 a_9644_26311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6411 vccd1 a_15667_21807# _1019_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6412 a_16984_15529# _0522_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6413 a_1863_24233# _0444_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X6414 vssd1 _0472_.X _0529_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6415 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_11527_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6416 a_22622_20149# a_22454_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6417 a_13261_10383# _0630_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6419 vccd1 _0866_.B a_6283_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6420 a_8393_9615# _0678_.Y a_8175_9527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6423 _1075_.Q a_3819_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6424 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6425 a_1591_21807# _0752_.Y io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6426 a_19785_14025# a_18795_13653# a_19659_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6427 a_15729_19453# _0860_.A a_15657_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6428 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6429 vssd1 a_9644_26311# _0820_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6430 a_20057_16885# _0662_.A1 a_20310_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X6431 a_4533_7913# a_4259_7669# a_4451_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6432 a_21610_24095# a_21442_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6433 a_10175_8029# a_9393_7663# a_10091_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6435 a_22454_20175# a_22181_20181# a_22369_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6436 vccd1 _0483_.X a_24315_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6438 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6439 a_4984_26703# _0833_.Y a_4729_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6440 a_4973_2223# a_3983_2223# a_4847_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6441 vssd1 a_1591_9839# _0466_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6442 _1053_.Q a_15963_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6444 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6445 a_27517_12381# a_26983_12015# a_27422_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6446 vssd1 _0722_.C a_3983_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6447 a_25030_15645# a_24757_15279# a_24945_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6449 a_14637_13647# _0511_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X6451 _0783_.A1 _0779_.X a_5731_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6452 _0555_.C1 a_11987_2473# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6454 _0630_.A2 _0474_.X a_14195_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6455 vccd1 a_8175_11989# _0655_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X6456 a_24995_13647# a_24131_13653# a_24738_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6457 a_1861_27069# a_1591_26703# a_1757_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6458 _0627_.X a_20911_15936# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6459 _0668_.X a_18059_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X6460 a_4621_16367# a_4429_16672# _0877_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6461 vccd1 _0583_.C a_16897_16395# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6462 a_25455_4765# a_24757_4399# a_25198_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6463 _1078_.D _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6464 vssd1 _1019_.CLK a_17231_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6465 vssd1 _1053_.CLK a_9503_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6466 a_15749_16189# _0504_.A a_15667_15936# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6467 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6468 vssd1 a_2807_4667# a_2765_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6470 vccd1 a_2547_3855# a_2715_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6473 vssd1 a_9503_19087# _0471_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6474 vssd1 io_in[1] a_3983_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6475 _0595_.D a_18427_2473# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6476 vssd1 _0445_.X a_9779_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6478 vssd1 a_2869_17501# a_2975_17461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6479 vccd1 _0959_.CLK a_10883_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6480 _0946_.Q a_15779_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6481 vssd1 a_27590_5599# a_27548_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6482 a_24665_13647# a_24131_13653# a_24570_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6484 a_10977_20175# a_10714_20541# a_10564_20407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6485 a_15553_4233# a_14563_3861# a_15427_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6486 vccd1 _0994_.CLK a_26983_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6488 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6489 vccd1 _0722_.A _0456_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6490 a_5821_13103# _0713_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X6491 a_9577_4399# a_9411_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6492 _0445_.B a_7520_23555# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6493 clkbuf_0_temp1.i_precharge_n.A a_9779_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6494 a_22737_3311# _0632_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6495 _0644_.X a_15667_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6496 a_15812_6005# _0669_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X6498 a_5078_30511# temp1.dcdc.Z vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X6499 a_20855_22351# a_20157_22357# a_20598_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6500 a_12801_15823# _0920_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6501 vccd1 a_16439_14557# a_16607_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6502 vccd1 a_23266_4511# a_23193_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6503 temp1.capload\[9\].cap.Y temp1.capload\[9\].cap_54.LO a_11797_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6504 vccd1 _0908_.CLK a_5455_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6505 a_25589_10383# _1006_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6506 temp1.capload\[7\].cap.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6507 a_1916_23983# _0764_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.209625 ps=1.295 w=0.65 l=0.15
X6508 a_14483_18543# _1075_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X6511 vccd1 _1033_.CLK a_23303_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6512 a_21809_19631# a_20819_19631# a_21683_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6513 a_22199_10499# _0648_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6514 a_13146_1653# a_12978_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6515 vssd1 a_23910_6005# a_23868_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6517 a_8175_9527# _0678_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6518 a_20819_16617# _0559_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6519 vssd1 a_4132_17429# _0813_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6520 temp1.dcdc.Z temp1.dcdc.A a_4160_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6521 vssd1 a_28015_3579# a_27973_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6523 a_23377_21269# a_23211_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6524 vssd1 a_2455_5853# a_2623_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6525 a_23303_12015# _1000_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6526 vssd1 _0840_.X _1078_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6527 _0445_.X a_5273_29687# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X6529 _0647_.B2 a_26267_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6530 a_25309_3311# a_25143_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6531 vccd1 _0972_.CLK a_19531_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6532 a_16182_4511# a_16014_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6533 a_16473_20719# a_15483_20719# a_16347_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6534 a_4403_22869# _0788_.C a_5466_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6535 vccd1 a_8546_1653# a_8473_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6536 _0637_.A1 a_10443_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R21 temp1.capload\[9\].cap_54.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6539 vssd1 _0582_.C a_21581_14219# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6540 _0994_.Q a_26635_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6541 a_26133_12015# a_25143_12015# a_26007_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6542 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9319_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6543 vccd1 a_4847_26525# a_5015_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6544 a_22879_20175# a_22181_20181# a_22622_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6545 vssd1 a_9999_1501# a_10167_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6546 _1048_.Q a_24243_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6548 a_25321_9615# _0665_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6551 a_11049_3311# a_10883_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6553 a_22454_20175# a_22015_20181# a_22369_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6554 vccd1 _0931_.CLK a_20635_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6555 clkbuf_0__0390_.A a_4075_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6556 vccd1 a_26099_4943# a_26267_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6558 a_25695_1679# _0619_.B1 a_25777_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6559 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_6808_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6561 _0998_.Q a_28015_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6562 _0814_.A2 a_3891_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6563 _1048_.Q a_24243_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6564 a_11067_19631# _0837_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X6565 vssd1 fanout23.X a_25143_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6567 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_12631_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6569 a_1766_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6570 _1072_.D a_26267_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6572 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_15023_28887# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6573 vssd1 _0740_.X a_4769_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6574 vccd1 a_21207_5755# a_21123_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6575 a_1945_6031# _0872_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6576 a_13403_1679# a_12705_1685# a_13146_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6577 vccd1 _0524_.X a_23303_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6578 a_19602_3855# a_19163_3861# a_19517_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6579 a_17267_22173# a_16569_21807# a_17010_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6580 vssd1 a_12299_10205# a_12467_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6581 vssd1 _0847_.A3 a_9945_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X6582 a_16061_10721# _0842_.A0 a_15975_10721# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6583 a_4132_17429# _0722_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6584 a_18059_17024# _1061_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6585 a_14737_2767# _0952_.Q a_14655_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6586 a_8067_4765# a_7369_4399# a_7810_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6587 vssd1 _0511_.D a_9595_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6588 _0940_.Q a_23415_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6589 a_2581_8751# a_1591_8751# a_2455_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6592 vccd1 _0702_.B1_N a_4259_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6595 a_21292_27247# a_20893_27247# a_21166_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6597 a_25497_9839# _1068_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6598 _0605_.C1 a_17783_12672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6599 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6600 _0684_.A2 _0466_.A a_9135_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6601 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6604 vccd1 temp1.dcdc.Z a_5078_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6607 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6610 a_17911_17821# a_17213_17455# a_17654_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6611 a_27057_8751# a_26891_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6613 _0650_.A1 a_28015_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6614 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6615 _0888_.CLK a_2787_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6616 _1081_.Q a_5015_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6617 a_5445_9615# _0710_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6618 a_2198_6005# a_2030_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6620 vccd1 _0456_.A a_3983_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6621 vccd1 a_27847_2589# a_28015_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6622 a_12150_8207# a_11877_8213# a_12065_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6623 a_18037_17455# a_17047_17455# a_17911_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6624 vccd1 _0975_.CLK a_22383_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6625 a_19234_1679# a_18795_1685# a_19149_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6626 vssd1 a_16929_17973# _0522_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X6627 a_12517_7439# _0637_.A1 a_12079_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6628 vssd1 a_20027_3855# a_20195_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6629 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10140_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6632 vssd1 _0922_.CLK a_1959_4951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6633 vssd1 _0511_.D a_14875_15325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X6634 a_25221_6575# _1003_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6635 vccd1 a_24738_13621# a_24665_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6636 vccd1 a_4882_19087# a_4988_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6637 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6638 a_17125_19631# _1050_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6639 a_15929_14191# _1057_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6640 a_8038_11837# _0466_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X6641 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10968_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6642 a_23193_4765# a_22659_4399# a_23098_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6643 a_21077_4765# a_20543_4399# a_20982_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6644 _0988_.Q a_10535_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6645 vccd1 _1076_.Q a_14453_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X6646 vccd1 _1015_.CLK a_25235_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6647 _1067_.D a_27555_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6648 a_17497_5487# _0622_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6649 a_20977_10901# _0662_.A1 a_21230_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X6650 vssd1 a_22035_24251# a_21993_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6651 a_24159_21263# a_23377_21269# a_24075_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6652 a_15052_9001# _0601_.B1 a_14950_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6654 a_25777_1999# _1072_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6656 vssd1 _0574_.C a_21213_17249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6657 _0670_.A1 a_13387_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6658 _0643_.B1 a_20025_10955# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X6660 a_5323_29111# _0809_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6661 a_27973_21807# a_26983_21807# a_27847_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6662 vccd1 a_26099_10383# a_26267_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6664 vccd1 a_12643_12559# a_12763_12879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X6665 a_22829_20719# _0963_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6667 a_27517_3677# a_26983_3311# a_27422_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6668 a_2039_9295# a_1591_9301# a_1945_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6669 vssd1 _0664_.A2 a_26317_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6670 vccd1 _0917_.CLK a_11711_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6671 vccd1 a_18539_11195# a_18455_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6672 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6673 a_8473_1679# a_7939_1685# a_8378_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6674 a_26873_6575# a_26707_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6675 a_15391_8323# _0675_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6676 a_4065_14237# _0460_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6677 a_9926_9269# a_9758_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6678 a_15236_10383# _0610_.X a_15134_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6681 a_26854_18655# a_26686_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6682 a_21345_15253# _0662_.A1 a_21598_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X6683 a_10862_11293# a_10589_10927# a_10777_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6684 a_19521_10089# _0588_.X a_19439_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6685 a_4590_2335# a_4422_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6686 a_5234_4917# a_5066_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6687 vssd1 _0479_.Y a_13459_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6689 vccd1 _0577_.C a_17139_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6690 vccd1 _0888_.CLK a_6651_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6691 vssd1 a_27698_4943# a_27804_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6693 _0487_.X a_17725_15073# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X6694 a_22917_14557# a_22383_14191# a_22822_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6695 vccd1 a_3302_4917# a_3229_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6696 a_5692_13077# _0768_.A1 a_5821_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6697 a_23193_26709# a_23027_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6698 a_4529_24847# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6699 a_10693_13353# _0735_.A2 _0714_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6700 a_25769_19997# a_25235_19631# a_25674_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6702 vssd1 _0821_.B a_11067_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6703 vssd1 a_24243_21237# a_24201_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6704 a_19973_15645# a_19439_15279# a_19878_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6705 vssd1 a_15795_1679# a_15963_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6706 vccd1 a_8327_6005# a_8243_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6707 a_4802_27247# clkbuf_0__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6708 a_22373_16367# _1067_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6709 a_17762_6031# a_17489_6037# a_17677_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6710 _0569_.X a_22383_14848# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6711 vccd1 a_25842_3829# a_25769_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6712 vccd1 a_25842_15797# a_25769_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6713 _0995_.Q a_24059_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6716 _0623_.D a_17415_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6719 a_9313_10703# _0596_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6720 a_3229_4943# a_2695_4949# a_3134_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6721 a_19325_25993# a_18335_25621# a_19199_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6723 a_17673_10927# a_17507_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6724 a_2915_28701# a_2217_28335# a_2658_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6725 a_2030_6941# a_1591_6575# a_1945_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6726 vssd1 a_5141_30199# io_out[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6728 _0523_.X a_17691_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6729 vccd1 fanout27.A a_18795_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6731 a_12625_14441# _0717_.A2 _0760_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6732 a_9669_5853# a_9135_5487# a_9574_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6733 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X6735 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_12631_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6736 _0860_.B a_11067_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X6737 vccd1 a_6319_3677# a_6487_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6738 a_10386_1653# a_10218_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6739 _0506_.A1 a_24335_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6740 a_25382_8181# a_25214_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6741 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6742 vssd1 a_15779_14709# a_15737_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6744 vccd1 a_16897_16395# _0522_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X6745 a_7663_15279# _0760_.B1 a_7841_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6747 a_4614_9615# _0696_.A1 a_4447_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X6748 vssd1 a_21610_13215# a_21568_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6749 a_6151_21781# _0797_.A2 a_6369_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X6750 a_22971_2767# a_22107_2773# a_22714_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6752 a_19728_4233# a_19329_3861# a_19602_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6753 a_10451_21263# a_9669_21269# a_10367_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6755 vssd1 a_16347_21085# a_16515_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6756 _0518_.Y _0836_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6758 a_4149_1135# a_3983_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6759 a_27149_16367# a_26983_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6760 a_18774_25615# a_18501_25621# a_18689_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6761 a_4847_1501# a_3983_1135# a_4590_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6762 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6763 _0815_.Y _0825_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6764 vssd1 a_14342_19061# a_14300_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6765 a_25547_13469# a_24849_13103# a_25290_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6767 vssd1 _0456_.A a_5642_19637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6768 vssd1 _1033_.CLK a_24775_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6769 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_14464_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6771 a_21901_18543# a_20911_18543# a_21775_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6772 a_21718_2589# a_21279_2223# a_21633_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6775 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8392_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6776 a_20157_22357# a_19991_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6777 vssd1 _0722_.C a_4137_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6778 a_23339_21085# a_22475_20719# a_23082_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6781 a_17029_7119# _0897_.Q a_16945_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6782 vccd1 _0529_.Y a_20299_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6783 a_3352_27081# a_2953_26709# a_3226_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6784 vccd1 a_13203_21237# a_13119_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6785 a_26099_10383# a_25235_10389# a_25842_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6786 a_24025_11471# _1014_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6787 a_14852_12015# a_14453_12015# a_14726_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6788 a_1674_26159# clkbuf_1_1__f_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6789 vssd1 a_22714_2741# a_22672_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6790 vssd1 a_16607_4667# a_16565_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6791 a_7561_12265# _0685_.B _0758_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6792 _0637_.A1 a_10443_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6793 vssd1 _0721_.A a_3155_21271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6794 vssd1 _0827_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6795 a_7097_3855# _0622_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6796 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X6798 a_27847_8029# a_26983_7663# a_27590_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6799 vssd1 a_10551_6031# a_10719_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6800 vccd1 _0515_.B1 a_20801_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X6801 _0932_.Q a_21023_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6803 a_19360_2057# a_18961_1685# a_19234_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6804 a_26007_10205# a_25143_9839# a_25750_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6808 vccd1 a_23361_13249# _0572_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6810 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6811 _0932_.Q a_21023_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6813 vccd1 a_7074_6687# a_7001_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6815 a_25401_21269# a_25235_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6816 a_15101_3311# _0946_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6818 a_7476_17455# _0717_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6819 a_2125_2223# a_1959_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6821 a_20161_14735# _1024_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6824 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6825 a_9718_20969# _0761_.B a_9636_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6826 vssd1 a_22587_22075# a_22545_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6827 a_25677_10205# a_25143_9839# a_25582_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6828 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10876_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6830 a_2198_8863# a_2030_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6831 a_2313_27247# _0837_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6832 vccd1 a_18125_18517# _0559_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X6833 vssd1 a_20414_14709# a_20372_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6834 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6835 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_6651_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6836 _0993_.D a_26267_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6837 vccd1 a_8307_17455# _1053_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6839 a_25842_1247# a_25674_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6842 a_25198_16479# a_25030_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6843 a_9742_1247# a_9574_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6845 a_4863_23413# _0813_.C1 a_5294_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X6847 a_19015_20175# a_18317_20181# a_18758_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6848 _0899_.Q a_11455_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6849 vccd1 a_18114_1247# a_18041_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6850 vssd1 _0533_.X a_23649_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6851 a_17083_26525# a_16385_26159# a_16826_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6852 _0993_.D a_26267_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6853 a_5165_19087# a_4988_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6854 vccd1 _0444_.A a_3983_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6855 a_15285_27791# _1053_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6856 a_10635_6031# a_9853_6037# a_10551_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6857 a_22465_15101# _0602_.A a_22383_14848# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6858 a_20349_6825# _0548_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6859 a_10335_7439# _0565_.X a_10198_7351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X6860 vccd1 _0745_.A2 a_5353_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6861 a_18509_2473# _0594_.D a_18427_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6863 a_11895_1135# _0850_.Y a_11895_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6864 _0639_.B a_13479_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6865 vssd1 a_20598_20149# a_20556_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6866 vssd1 _0524_.X a_11865_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6867 a_14559_17705# _0797_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6868 vccd1 a_27590_14303# a_27517_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6869 a_15354_3423# a_15186_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6870 a_17720_13353# _0602_.X a_17618_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6871 vssd1 _0685_.B _0686_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6872 a_22990_19061# a_22822_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6873 a_27337_5487# _0650_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6874 vssd1 _0797_.A1 a_10331_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6875 a_19697_16617# _0963_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6876 a_18961_1685# a_18795_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6878 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6880 a_8079_28500# _0820_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6881 a_20648_21641# a_20249_21269# a_20522_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6882 a_27498_8863# a_27330_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6883 vssd1 a_19827_13621# a_19785_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6885 a_7733_4233# a_6743_3861# a_7607_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6886 a_9581_7663# _0613_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6887 vssd1 _0917_.CLK a_10423_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6888 _0847_.A2 a_11435_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6889 a_17761_19631# a_16771_19631# a_17635_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6890 vssd1 a_13735_12925# _0572_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X6891 _0599_.X a_14287_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6892 a_13432_28585# a_13183_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6893 vssd1 a_12207_18909# a_12375_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6894 a_6641_15823# _0812_.A2 a_6559_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6895 a_15196_8751# _0961_.D a_14621_8897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X6896 vssd1 a_8031_16911# _0836_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6898 a_24201_21641# a_23211_21269# a_24075_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6899 a_22702_15279# _1047_.D a_22612_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X6900 vccd1 a_12777_16885# _0739_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6901 a_23657_6031# _0607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6903 _0445_.A _0440_.C a_6813_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6904 a_14559_17705# _0798_.A2 a_14341_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6905 a_2156_6575# a_1757_6575# a_2030_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6907 a_27422_17821# a_26983_17455# a_27337_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6908 vccd1 _0847_.A3 a_11842_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6909 _0670_.A1 a_13387_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6910 a_12052_30761# a_11803_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6911 vssd1 a_16035_4943# _1030_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6912 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_4988_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6913 a_12069_2223# _0902_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6914 a_22143_2589# a_21279_2223# a_21886_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6915 vssd1 a_25915_9117# a_26083_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6916 _0545_.B1 a_19439_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X6917 a_17673_10927# a_17507_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6920 vssd1 _0549_.X a_15115_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6921 a_5356_29429# _0445_.A a_5273_29687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6922 vccd1 a_14967_20175# a_15135_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6924 a_4973_26159# a_3983_26159# a_4847_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6925 a_18519_5487# _0631_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6927 vccd1 a_5491_4943# a_5659_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6929 a_27249_10383# _0647_.B2 a_27167_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6930 a_10977_20175# _0798_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6932 a_27337_12015# _1013_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6933 vccd1 a_15319_12283# a_15235_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6934 a_22751_7663# _0506_.A2 a_22929_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6935 vssd1 a_14967_20175# a_15135_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6936 a_12318_13621# a_12150_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6937 vccd1 _1030_.CLK a_20175_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6939 vssd1 a_15630_16479# a_15588_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6940 a_9666_8029# a_9227_7663# a_9581_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6941 a_21844_2223# a_21445_2223# a_21718_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6942 _0861_.B1 a_3799_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6943 a_25674_4943# a_25235_4949# a_25589_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6945 a_16123_25615# _0861_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6946 a_26183_21263# a_25401_21269# a_26099_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6947 vccd1 _0711_.A a_5245_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X6948 a_21867_24349# a_21003_23983# a_21610_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6949 vccd1 _0648_.A2 a_23385_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6950 a_2129_4399# _0870_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6951 vccd1 temp1.capload\[15\].cap_45.LO temp1.capload\[15\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6952 a_27053_20719# a_26063_20719# a_26927_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6953 vssd1 a_17727_3855# a_17895_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6955 a_19613_11471# _0648_.A2 a_19697_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6956 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6957 a_11877_21085# a_11343_20719# a_11782_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6958 _0778_.A2 a_8123_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6959 a_12150_13647# a_11877_13653# a_12065_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6960 a_17673_1135# a_17507_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6961 vssd1 a_21023_22325# a_20981_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6962 a_22009_10089# _0663_.X a_21913_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6963 _0445_.A _0440_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6964 _0751_.B1 a_10331_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X6965 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10791_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6966 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12355_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6968 a_8038_11510# _0466_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6970 a_7829_15529# _0439_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6971 ANTENNA_7.DIODE a_3983_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6972 a_2401_2773# a_2235_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6973 a_22917_8213# a_22751_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6974 a_6737_16143# _0735_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6975 a_11965_6575# _0674_.A1 a_11527_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6977 vccd1 a_22622_16885# a_22549_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6978 a_21537_24349# a_21003_23983# a_21442_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6979 a_9407_18793# _0797_.A1 a_9189_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6980 _1062_.CLK a_19439_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6981 a_2823_1501# a_2125_1135# a_2566_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6983 _0553_.C1 a_23487_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6984 a_8256_20291# _0761_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6985 vccd1 a_19659_13647# a_19827_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6986 a_18041_1501# a_17507_1135# a_17946_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6987 a_9297_7497# a_8307_7125# a_9171_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6988 a_12316_24135# _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6989 a_23247_19087# a_22549_19093# a_22990_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6990 _0680_.Y _0778_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6991 a_23361_13249# _0572_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X6992 _0870_.Y a_4981_21024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X6993 a_20395_2767# a_19531_2773# a_20138_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6994 fanout37.A a_3523_6039# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6995 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6996 vccd1 a_25455_2589# a_25623_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6998 a_24251_6031# a_23469_6037# a_24167_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6999 a_4035_13077# _0758_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X7000 vccd1 _0511_.D a_10202_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X7001 vccd1 a_20025_10955# _0643_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X7002 vssd1 a_19659_13647# a_19827_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7003 a_1933_27069# _0831_.B a_1861_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X7004 vssd1 a_26267_21237# a_26225_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7005 io_out[6] a_5141_30199# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7007 a_4439_9001# _0711_.A a_4221_8725# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X7008 _1035_.Q a_24979_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7009 vssd1 _0672_.C1 a_16863_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7010 vccd1 _0863_.A1 a_14319_20747# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7011 vccd1 _0572_.A1 a_23792_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7012 a_25769_25615# a_25235_25621# a_25674_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7013 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7014 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7015 a_13080_24847# _0829_.A1 a_12777_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7017 a_2125_1135# a_1959_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7018 _0946_.D a_15871_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7019 a_25198_5599# a_25030_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7020 vssd1 a_4037_11989# _0791_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7022 a_9313_20495# _0847_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7023 a_24719_1679# a_23855_1685# a_24462_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7024 a_13551_6031# _0644_.A2 a_13729_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7025 a_12995_24527# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7026 a_23466_17999# a_23027_18005# a_23381_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7027 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7030 a_7067_28918# _0825_.A1 a_6608_29111# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7031 a_23331_1501# a_22549_1135# a_23247_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7033 vssd1 a_8123_20719# _0827_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7035 vccd1 clkbuf_1_0__f_io_in[0].X a_1591_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7036 vccd1 _0506_.A2 a_22825_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7037 vssd1 _0869_.B1 _0445_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7039 a_16523_14557# a_15741_14191# a_16439_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7040 vssd1 a_20138_2741# a_20096_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7041 a_10048_31599# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7042 vssd1 clkbuf_1_1__f__0390_.A a_2686_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7044 a_26593_26159# a_25603_26159# a_26467_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7045 a_25842_19061# a_25674_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7047 a_15703_2589# a_15005_2223# a_15446_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7049 _0928_.Q a_28015_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7050 vccd1 _0797_.B1 a_6151_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X7052 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X7054 a_15887_16733# a_15023_16367# a_15630_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7055 _0634_.B1 a_18519_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7056 vccd1 a_16495_5487# fanout24.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7057 a_19521_12675# _0584_.X a_19439_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X7058 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7059 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_13432_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7060 _0658_.B1 a_17539_16161# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7061 a_14689_15325# a_14287_15279# a_14603_15325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X7062 vssd1 _0580_.C1 a_16553_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X7063 temp1.capload\[11\].cap.Y temp1.capload\[11\].cap_41.LO a_3885_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7064 a_15833_12559# _0918_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7066 a_20525_20175# a_19991_20181# a_20430_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7067 a_10055_24527# _0444_.B _0819_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X7068 vssd1 a_24462_1653# a_24420_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7069 _0545_.A1 a_5567_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7071 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14563_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7073 a_15369_9295# _0652_.C a_15563_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7074 a_15557_16733# a_15023_16367# a_15462_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7075 vccd1 a_17930_6005# a_17857_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7076 a_4985_12061# _0807_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7077 vssd1 clkbuf_1_1__f_net57.A a_1674_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7078 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_12052_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7079 a_22181_22357# a_22015_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7080 _0932_.D a_21115_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7081 vssd1 a_16101_18517# _0667_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X7082 a_23592_27081# a_23193_26709# a_23466_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7084 vccd1 _0917_.CLK a_10423_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7085 vssd1 a_23358_8181# a_23316_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7086 a_20245_1135# _0976_.Q a_19899_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7087 a_17401_17455# _1059_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7088 a_9217_14441# _0714_.B1 a_9301_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7089 a_19852_9615# _0582_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7090 vccd1 _1079_.Q _0479_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7091 vssd1 a_2198_6687# a_2156_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7092 vssd1 a_13403_1679# a_13571_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7093 a_20046_15391# a_19878_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7095 _1018_.D a_23047_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7097 a_8259_11837# _0836_.A a_7896_11703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7098 a_11913_13336# _0511_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X7099 vccd1 _0572_.A2 a_21813_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7101 a_16548_10901# _0991_.D a_16768_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7102 _0832_.A a_1757_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X7103 _1018_.D a_23047_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7104 vssd1 _0797_.A1 a_12527_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X7106 a_11884_13103# a_11435_13103# a_11582_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7107 vccd1 _0527_.X a_21127_11809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7108 a_26225_7497# a_25235_7125# a_26099_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7109 _0662_.A3 a_14453_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X7110 a_22825_4399# a_22659_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7111 a_20709_4399# a_20543_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7112 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10048_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7113 a_9792_7663# a_9393_7663# a_9666_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7116 _0814_.B1 _0827_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7117 vccd1 a_18850_21237# a_18777_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7120 vccd1 temp1.capload\[2\].cap_47.LO temp1.capload\[2\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7121 vssd1 a_21886_2335# a_21844_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7122 a_25800_5321# a_25401_4949# a_25674_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7123 _1075_.Q a_3819_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7124 vccd1 a_22863_26427# a_22779_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7126 a_18497_18319# _1018_.D a_18059_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7127 vccd1 a_27847_15645# a_28015_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7130 _0778_.B1 a_5089_14851# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X7131 _0839_.B a_2655_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7132 vccd1 _0580_.A1 a_16984_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7133 a_22547_9295# _0621_.X a_22465_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X7134 _0529_.Y _0472_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7135 a_11322_3677# a_11049_3311# a_11237_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7136 a_13487_1679# a_12705_1685# a_13403_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7137 _0672_.C1 a_14747_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7139 a_12069_4943# _0673_.B2 a_11987_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7140 a_25750_3423# a_25582_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7141 _0835_.Y _0845_.C1 a_4729_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7142 a_25225_14191# _0966_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7143 vssd1 a_18703_12567# _0504_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7144 a_27513_13103# a_26523_13103# a_27387_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7145 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_12355_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7146 vccd1 _0836_.A a_1775_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7147 a_27517_24349# a_26983_23983# a_27422_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7148 a_24673_11177# _1011_.D a_24591_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7149 vssd1 a_18114_11039# a_18072_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7150 a_10791_17705# _0472_.X a_11041_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7151 a_13805_9673# a_12815_9301# a_13679_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7152 vccd1 a_3651_26703# a_3819_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7153 io_out[2] _0752_.Y a_1591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7154 a_17909_16395# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7155 vccd1 _0959_.CLK a_12447_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7156 _0778_.Y _0778_.B1 a_5455_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7157 a_2547_3855# a_1849_3861# a_2290_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7158 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7159 a_14917_23439# _1053_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7160 vccd1 a_8123_20719# _0827_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7161 a_4663_3855# a_3965_3861# a_4406_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7162 vccd1 a_4811_10383# _0845_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7165 a_23690_13353# _0570_.X a_23610_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7167 vssd1 a_10791_16919# _0935_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7169 a_6423_8903# _0681_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X7170 vssd1 _0513_.X a_13889_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7171 a_22461_2767# _0497_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7172 a_22737_14191# _0939_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7174 _1046_.D a_23599_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7175 vccd1 a_9095_10615# _0597_.A2_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X7176 a_14453_12015# a_14287_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7177 vssd1 a_19367_25589# a_19325_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7178 a_21031_21263# a_20249_21269# a_20947_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7180 a_5731_13967# _0778_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7181 a_10183_9295# a_9319_9301# a_9926_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7182 vccd1 _0524_.X a_21127_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7183 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7184 vssd1 a_26927_21085# a_27095_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7185 a_18456_7913# _0533_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7186 vssd1 a_20057_16885# _0557_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X7187 a_26486_23007# a_26318_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7188 a_5491_4943# a_4627_4949# a_5234_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7190 a_5509_7093# _0656_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X7192 a_25129_12559# _1000_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7193 a_18590_20175# a_18151_20181# a_18505_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7194 a_24021_20181# a_23855_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7195 vssd1 _0717_.A2 a_6639_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X7196 _0497_.A1 a_15595_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7197 _1001_.Q a_25807_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7199 a_25769_4943# a_25235_4949# a_25674_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7200 vccd1 _0479_.Y a_13459_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7201 a_2405_28335# _0845_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7202 vccd1 _0582_.C a_22015_18112# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7203 vccd1 a_9284_10901# _0685_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7204 a_13432_29967# a_13183_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7205 a_12788_29673# a_12539_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7206 _1001_.Q a_25807_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7207 _0580_.A1 a_10627_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7208 vccd1 _0831_.B a_1757_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X7209 io_out[3] a_1585_24135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7210 vccd1 _0861_.B1 a_15576_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X7213 a_12999_2223# _0535_.X a_13177_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7214 vssd1 _0522_.B1 a_18232_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X7216 vccd1 a_20598_20149# a_20525_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7217 _0456_.A _0722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7218 vccd1 a_10110_11445# a_10037_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7219 vccd1 _0529_.Y a_19439_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7220 vccd1 _0582_.C a_17783_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7222 a_10416_27247# _0821_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7223 _0444_.Y _0444_.A a_1775_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7224 a_1591_21807# _0444_.A io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X7225 a_16431_21085# a_15649_20719# a_16347_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7226 vssd1 _0522_.X a_17691_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7227 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7228 _0580_.A1 a_10627_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7229 _0892_.D a_25623_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7230 a_16439_14557# a_15741_14191# a_16182_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7231 a_13257_17821# _1078_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X7232 _0604_.B a_10811_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7233 _0505_.A1 a_25807_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7234 a_2198_6005# a_2030_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7235 a_16771_9001# _0630_.A2 a_16853_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7236 a_4253_9839# _0696_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7237 a_11797_30287# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7238 a_16014_4765# a_15741_4399# a_15929_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7239 a_16014_14557# a_15575_14191# a_15929_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7241 vccd1 _1015_.CLK a_26891_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7243 vssd1 a_8803_1679# a_8971_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7244 a_12355_8751# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X7245 vssd1 _0651_.C a_22199_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X7246 vccd1 a_25715_13371# a_25631_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7247 a_10643_1679# a_9779_1685# a_10386_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7248 _0594_.D a_19899_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7249 a_26099_4943# a_25401_4949# a_25842_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7250 a_22097_5737# _1008_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7254 a_8270_21237# a_8102_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7255 a_15097_1685# a_14931_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7256 a_11760_26935# _0825_.A0 a_11902_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7257 a_24945_5487# _1031_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7258 vccd1 _0445_.A a_5273_29687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7259 a_6795_14343# a_6938_14237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7260 vssd1 a_10643_2767# a_10811_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7261 a_26041_1999# _1035_.Q a_25695_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7262 vccd1 _0524_.X a_18059_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7263 vccd1 a_6779_2589# a_6947_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7264 a_17946_11293# a_17673_10927# a_17861_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7265 a_23339_21085# a_22641_20719# a_23082_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7266 vssd1 _0708_.B1 a_4864_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X7267 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X7268 vssd1 a_3298_17143# _0812_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7269 a_10083_1501# a_9301_1135# a_9999_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7270 _0529_.Y a_10814_15797# a_10594_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7271 vssd1 a_23047_22325# a_23005_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7272 a_8937_3855# _0902_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7273 vccd1 _0745_.A2 a_4255_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7274 vssd1 _0836_.A _0508_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7275 vssd1 a_26467_26525# a_26635_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7276 a_25030_4765# a_24591_4399# a_24945_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7278 a_18673_5487# _0631_.B a_18601_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7279 a_27590_25183# a_27422_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7280 vccd1 a_22311_2491# a_22227_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7282 vssd1 a_10386_1653# a_10344_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7284 vssd1 a_27847_25437# a_28015_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7285 vssd1 _0524_.X a_13337_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7286 vssd1 _0590_.X a_18427_2473# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7287 _0616_.B1 a_16771_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7288 a_11969_24847# _0840_.A1 _0825_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X7290 vccd1 _0491_.X a_14737_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7291 a_9774_23759# _0847_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X7292 a_2683_2767# a_2401_2773# a_2589_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X7293 a_16209_7913# _0549_.C1 a_16127_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7294 a_3983_31849# _0814_.B1 a_4065_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7295 vccd1 _0814_.A2 a_6559_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7296 vssd1 a_11435_8751# _0842_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X7297 vssd1 _1019_.CLK a_21279_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7298 vssd1 _0670_.A2 a_15277_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X7299 a_4769_22895# _0740_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7301 vssd1 clkbuf_1_0__f_io_in[0].X a_1959_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7302 a_2686_15823# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7303 vssd1 a_9834_7775# a_9792_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7305 a_20057_16885# _0512_.X a_20214_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X7306 a_2039_22057# _0814_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7307 vssd1 _1028_.CLK a_9135_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7308 a_13809_4943# a_13275_4949# a_13714_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7309 vccd1 _0872_.A1 a_4705_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7312 a_17309_1679# _0515_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7313 a_6635_7913# _0689_.X _0694_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7314 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7315 vccd1 a_3451_25589# _1078_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7316 vccd1 a_10567_19061# _0773_.A1_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7317 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X7318 vccd1 temp1.dcdc.Z a_5078_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
D3 vssd1 _0849_.X sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X7320 _0545_.A1 a_5567_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7321 vssd1 a_1959_4951# _0908_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7322 vssd1 _0710_.A2 a_5717_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
X7323 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7324 a_4988_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7325 a_25915_17821# a_25217_17455# a_25658_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7326 a_19045_15797# _0512_.A a_19298_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7327 vccd1 a_27847_14557# a_28015_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7328 a_14569_1385# _0641_.D1 _0642_.D_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.755 ps=3.51 w=1 l=0.15
X7329 a_10543_13647# a_9761_13653# a_10459_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7330 vccd1 _0961_.D a_15052_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7332 vccd1 _0873_.A _0873_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7333 a_6559_10383# _0685_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7334 vccd1 _1021_.Q a_21502_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7335 vssd1 _0850_.A a_7520_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7336 _1003_.Q a_26083_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7337 a_5692_13077# _0713_.A1 a_5915_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7338 vccd1 _0758_.A1 a_7561_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7339 vccd1 a_25290_13215# a_25217_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7340 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_12532_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7341 vssd1 _0518_.Y a_15693_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7342 vccd1 _1030_.CLK a_17323_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7343 vssd1 _1028_.CLK a_10423_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7344 a_12778_21237# a_12610_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7346 _0784_.A1 a_11936_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7347 a_9516_17289# a_9117_16917# a_9390_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7348 vccd1 _0529_.Y a_18001_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7349 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7350 a_17838_23007# a_17670_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7351 vssd1 a_17930_6005# a_17888_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7353 vccd1 a_9999_5853# a_10167_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7355 vssd1 _0444_.A a_3983_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7356 vccd1 _0845_.C1 a_1775_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7357 a_19329_26709# a_19163_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7358 vssd1 _0807_.A _0880_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7359 vssd1 _0613_.C1 a_14805_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X7360 vccd1 a_20563_2741# a_20479_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7361 vssd1 _0763_.B1 a_8176_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X7362 a_7090_5853# a_6817_5487# a_7005_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7363 vccd1 a_25915_9117# a_26083_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7364 a_27314_6687# a_27146_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7366 a_27931_22173# a_27149_21807# a_27847_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7367 _0833_.A a_7939_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X7373 vccd1 a_10367_21263# a_10535_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7374 vccd1 _0472_.X a_12441_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X7375 a_14189_7235# _0544_.C a_14093_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X7376 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13432_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7377 a_25582_6031# a_25309_6037# a_25497_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7378 vssd1 a_25842_19743# a_25800_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7380 a_8527_21263# a_7829_21269# a_8270_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7381 a_27314_6687# a_27146_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7383 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_13183_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7384 a_5466_22895# _0847_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7385 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7386 vssd1 a_27387_13469# a_27555_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7387 a_9669_21269# a_9503_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7388 vssd1 a_10367_21263# a_10535_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7390 vccd1 a_24887_1653# a_24803_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7391 _0891_.D a_22035_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7393 a_15391_13103# _1076_.Q a_15285_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7394 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15844_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7395 a_7291_20175# _0784_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7396 a_24236_11849# a_23837_11477# a_24110_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7398 a_11950_15391# a_11782_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7401 _0564_.D a_22291_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X7402 a_18758_4917# a_18590_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7403 vssd1 _0527_.X a_23457_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7404 a_21568_23983# a_21169_23983# a_21442_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7405 vccd1 _0850_.Y a_11895_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X7406 a_25589_21263# _0992_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7407 a_22537_15101# _1048_.Q a_22465_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7408 a_17945_2057# a_16955_1685# a_17819_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7409 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7410 _0566_.A1 a_7683_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7411 a_2455_9117# a_1591_8751# a_2198_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7412 _0438_.A a_2715_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7413 a_17811_10383# a_17029_10389# a_17727_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7414 a_14772_1385# _0638_.X a_14668_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X7416 a_10693_13353# _0546_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X7417 a_9644_26311# _0825_.A1 a_9786_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7418 _0998_.D a_26911_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7419 vssd1 a_21759_27515# a_21717_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7420 a_14737_4399# _0479_.Y a_14655_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7421 vccd1 _0659_.X a_22081_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7422 vccd1 a_28015_5755# a_27931_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7423 a_4802_27247# clkbuf_0__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X7424 _0995_.Q a_24059_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7426 a_20993_1385# _1040_.Q a_20911_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7427 a_22411_6603# _0504_.A a_22325_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7428 _0548_.B2 a_23139_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7429 vccd1 _0845_.A1 a_5635_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7430 vccd1 a_25623_15547# a_25539_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7431 vccd1 io_in[6] a_1591_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7432 a_25030_2589# a_24757_2223# a_24945_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7433 a_26785_4399# _1008_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7434 vccd1 _0995_.CLK a_23027_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7435 a_2566_2335# a_2398_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7436 vccd1 _0662_.A3 a_16895_5281# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7437 vssd1 _0972_.CLK a_16863_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7438 vssd1 a_12778_21237# a_12736_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7439 a_20214_16911# _1017_.D a_20057_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7441 vccd1 _0835_.A1 a_11895_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7442 vssd1 a_17987_1653# a_17945_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7443 vccd1 fanout9.A a_12999_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7444 vccd1 a_4170_20291# _0764_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X7445 vccd1 a_15611_3677# a_15779_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7446 a_18317_4949# a_18151_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7448 vccd1 _0999_.CLK a_26983_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7449 a_14089_19087# _0936_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7450 a_25156_4399# a_24757_4399# a_25030_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7451 a_25455_5853# a_24591_5487# a_25198_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7452 a_12318_6005# a_12150_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7453 a_24209_1679# _0976_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7454 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7455 vccd1 a_23891_26703# a_24059_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7456 a_11269_16367# _0827_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7457 _0613_.C1 a_13183_7232# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7459 a_15511_3855# a_14729_3861# a_15427_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7460 vssd1 fanout27.A a_17507_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7461 vccd1 a_5325_8181# _0711_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X7462 a_19605_10089# _0940_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7463 a_13514_10357# a_13346_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7464 vssd1 a_6516_18695# _0797_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7465 vccd1 a_13054_2741# a_12981_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7466 vssd1 _0835_.A1 a_12428_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7468 vccd1 _0679_.A1 a_8116_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X7470 a_17673_1135# a_17507_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7471 _0865_.Y a_12356_19203# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7472 a_23105_8207# _0590_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7473 vccd1 a_2455_6031# a_2623_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7474 a_9095_20407# _0813_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X7476 a_21173_19631# _1023_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7477 vssd1 a_27847_3677# a_28015_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7478 vssd1 _0535_.X a_11597_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7479 a_13514_22325# a_13346_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7480 a_26183_3855# a_25401_3861# a_26099_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7481 _0917_.D a_12743_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7484 a_10367_21263# a_9503_21269# a_10110_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7485 a_14453_7663# a_14287_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7486 _0825_.A0 _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7487 vccd1 _0742_.A2 a_4769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7488 _0833_.A a_7939_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7489 a_22549_1135# a_22383_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7490 a_14870_9001# _0600_.X a_14621_8897# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7491 a_1674_26159# clkbuf_1_1__f_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X7492 a_20985_8751# a_20819_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7493 _0572_.A2 a_13735_12925# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X7494 a_17415_5737# _0535_.X a_17497_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7495 _0615_.A1 a_20195_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7496 a_23358_8181# a_23190_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7497 vssd1 _1063_.Q a_21468_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X7498 a_5642_19637# _0456_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7499 a_26601_18543# _1067_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7500 vccd1 a_11490_3423# a_11417_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7504 vssd1 _0523_.B1 a_19877_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X7505 a_13346_22351# a_13073_22357# a_13261_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7508 a_14668_1385# _0639_.X a_14569_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.1725 ps=1.345 w=1 l=0.15
X7509 a_10037_21263# a_9503_21269# a_9942_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7510 a_8848_15055# _0833_.A a_8545_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7511 vccd1 a_26835_11293# a_27003_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7513 vssd1 a_23891_17999# a_24059_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7514 _0845_.A1 a_2991_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7515 vccd1 _0479_.Y a_11435_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7516 a_19402_13621# a_19234_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7517 a_24462_1653# a_24294_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7518 a_16029_20175# _0840_.A1 _0863_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7519 _0527_.X a_14603_15325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7520 a_9857_11471# _0985_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7521 a_21633_2223# _0575_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7522 a_2125_1135# a_1959_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7523 _1047_.D a_25163_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7524 a_4517_28701# a_3983_28335# a_4422_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7525 a_2823_1501# a_1959_1135# a_2566_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7526 vssd1 _0522_.B1 a_17128_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X7527 a_27973_15279# a_26983_15279# a_27847_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7530 vccd1 a_6062_3423# a_5989_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7531 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7532 a_8205_13647# _1080_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7533 vssd1 _0998_.D a_21836_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X7534 _1047_.D a_25163_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7537 a_3141_26703# _0835_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7538 vssd1 clkbuf_1_0__f_io_in[0].X a_1591_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7539 a_12709_4399# _0951_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7540 a_23385_12015# _0583_.A a_23303_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7541 a_19234_13647# a_18961_13653# a_19149_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7542 a_11987_4943# _0535_.X a_12069_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7543 vccd1 _1028_.CLK a_13275_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7544 vccd1 a_10351_9269# a_10267_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7545 a_20345_20175# _1061_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7546 _0489_.C1 a_23119_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7547 a_25842_10357# a_25674_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7548 a_12525_21263# _0934_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7549 vccd1 _0999_.CLK a_25235_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7550 vssd1 _0512_.A a_18611_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X7551 a_4530_9295# a_4259_9295# a_4447_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7552 vccd1 _0860_.A _0861_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7553 a_5001_15823# _0807_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7554 a_11040_29673# a_10791_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7555 _0839_.Y _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7556 _0753_.A2 a_9687_19881# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X7557 a_8377_18543# _0833_.A a_7939_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7559 vssd1 _0825_.A1 _0825_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7560 a_4769_23145# _0809_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.585 pd=2.17 as=0.135 ps=1.27 w=1 l=0.15
X7561 a_1757_26703# a_1591_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X7562 vccd1 a_3983_3311# ANTENNA_7.DIODE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7563 a_18130_11471# a_17691_11477# a_18045_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7564 a_13104_2057# a_12705_1685# a_12978_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7565 a_15921_28169# a_14931_27797# a_15795_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7566 a_15105_11471# _0988_.Q a_15023_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7567 vccd1 a_26099_21263# a_26267_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7568 vccd1 a_11619_29423# fanout10.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7569 vssd1 a_18263_23163# a_18221_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7570 a_25539_22173# a_24757_21807# a_25455_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7571 vssd1 _0860_.A a_10703_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7573 a_24719_1679# a_24021_1685# a_24462_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7574 _0991_.D a_16055_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7575 a_23385_16617# _0966_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7576 _0515_.B2 a_18355_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7577 a_10041_22351# _1055_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7578 a_5173_20719# _0803_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7579 vccd1 a_7037_29177# a_7067_28918# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7580 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X7581 _0842_.A0 a_11435_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X7582 vssd1 a_26099_21263# a_26267_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7583 a_2539_6941# a_1757_6575# a_2455_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7585 a_18689_25615# _1061_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7586 a_25401_15829# a_25235_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7587 a_2593_15325# _0460_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7588 vccd1 _0572_.A2 a_25593_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7589 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7590 _0642_.C a_12079_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X7591 vssd1 a_28015_7931# a_27973_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7592 vssd1 _0847_.A3 a_12694_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
X7593 vssd1 a_12759_3855# a_12927_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7594 _1003_.Q a_26083_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7595 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_15667_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7597 a_23615_8207# a_22917_8213# a_23358_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7598 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_18308_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7599 vssd1 a_11950_15391# a_11908_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7601 vccd1 a_10811_1653# a_10727_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7602 _0847_.A2 a_11435_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7603 vssd1 _0821_.Y a_7755_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7604 _0893_.D a_26267_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7606 vssd1 a_9999_5853# a_10167_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7607 a_3713_16911# _0456_.B a_3298_17143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X7608 a_10147_15529# _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X7609 a_24209_22351# _0928_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7610 a_17182_18319# _1052_.D a_17092_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X7611 vssd1 a_8031_16911# _0836_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7612 a_14260_29967# a_14011_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7614 vccd1 a_17473_14337# _0630_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X7615 vccd1 _1028_.CLK a_14563_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7616 vssd1 _0535_.X a_13069_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X7617 vccd1 _0512_.A a_14655_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7618 a_13616_29673# a_13367_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7620 a_19347_8207# _0515_.B1 a_19429_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7621 a_16258_18793# _0577_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X7623 a_20717_10703# _0890_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7625 vssd1 _0839_.B _0839_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7626 a_20220_17231# _0582_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7627 _0893_.CLK a_23487_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7628 _0791_.A2 a_5091_12021# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X7629 a_17217_3855# _0671_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7630 vssd1 a_25198_4511# a_25156_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7631 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7632 a_23381_17999# _0963_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7633 a_12705_1685# a_12539_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7634 a_19981_1385# _0970_.Q a_19899_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7635 a_20437_21263# _0930_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7636 a_7737_4765# a_7203_4399# a_7642_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7637 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7638 a_4534_25071# _0829_.A1 a_4035_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X7639 clkbuf_0__0390_.A a_4075_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7640 a_25079_13647# a_24297_13653# a_24995_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7641 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7644 a_27337_23983# _0928_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7645 vccd1 _0722_.A a_4324_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7646 vssd1 a_23634_17973# a_23592_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7647 vccd1 _0776_.A2 _0745_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7648 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7649 vssd1 _0471_.X a_7226_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7650 vssd1 _0695_.A2 a_4101_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7651 vssd1 _0758_.A1 a_5455_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7653 a_26099_7119# a_25235_7125# a_25842_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7654 _0814_.A2 a_3891_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7656 a_10769_18319# _0749_.A1 a_10331_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7657 vccd1 _0975_.CLK a_21279_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7659 a_17473_14337# _0629_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7660 _0961_.D a_10903_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7661 vccd1 fanout27.A a_17507_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7662 a_11764_20149# _0837_.A1 a_11893_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7664 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A _0816_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7665 _0566_.A1 a_7683_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7666 a_11956_13103# a_11913_13336# a_11884_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X7668 a_22369_22351# _1017_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7669 vccd1 _0917_.CLK a_9503_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7670 vccd1 a_11067_19631# _0860_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X7671 vccd1 _0836_.A a_11458_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7672 vssd1 _0624_.C a_17971_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7674 a_10133_1679# _0639_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7675 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7676 vccd1 a_25198_2335# a_25125_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7677 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE a_8215_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7679 vssd1 a_22162_21919# a_22120_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7680 vssd1 _0735_.A2 a_9573_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.099125 ps=0.955 w=0.65 l=0.15
X7682 _0789_.B1 a_5913_25335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7683 a_14655_11177# _0474_.X _0565_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7684 a_6750_29245# _0825_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7686 _0538_.C1 a_11251_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7687 a_12161_7119# _0487_.X a_12245_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7688 a_14453_12015# a_14287_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7689 a_26099_21263# a_25235_21269# a_25842_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7690 vccd1 _0658_.B1 a_16293_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7692 vccd1 a_7435_26324# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7694 vssd1 a_27590_12127# a_27548_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7695 a_16937_22173# a_16403_21807# a_16842_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7697 a_6641_15823# _0736_.B1 a_6725_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7698 a_19697_11471# _0962_.D a_19613_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7699 a_25306_6941# a_25033_6575# a_25221_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7700 a_9581_7663# _0613_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7701 a_13165_2473# _0951_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7702 vccd1 a_3451_25589# a_3367_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R22 vccd1 temp1.capload\[15\].cap_45.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7704 vccd1 _0847_.A3 a_10055_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X7705 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7706 vssd1 _0487_.X a_15369_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7707 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11040_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7709 a_6906_6941# a_6467_6575# a_6821_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7710 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_4811_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7711 a_17853_4233# a_16863_3861# a_17727_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7712 a_26183_15823# a_25401_15829# a_26099_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7713 a_27973_14191# a_26983_14191# a_27847_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7715 a_11333_5737# _0986_.D a_11251_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7716 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X7717 vccd1 _0722_.C a_5549_17719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X7718 a_19429_8527# _0515_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7719 a_5816_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7720 vccd1 a_25750_6005# a_25677_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7722 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7723 a_19728_27081# a_19329_26709# a_19602_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7724 a_19793_17455# _0937_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7725 a_11877_15645# a_11343_15279# a_11782_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7727 a_24554_2741# a_24386_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7729 a_10202_18517# _1078_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7730 _1077_.Q a_3083_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7731 a_4747_3855# a_3965_3861# a_4663_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7732 a_1757_6037# a_1591_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7734 a_17677_6031# _0615_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7735 _0825_.S _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7737 vccd1 a_23615_8207# a_23783_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7738 a_20982_3677# a_20543_3311# a_20897_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7739 a_25401_10389# a_25235_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7740 _0861_.A2 a_16904_24643# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X7741 vssd1 _0833_.A _0574_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7742 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7743 vssd1 _0833_.A _0833_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7744 a_17857_11477# a_17691_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7745 vssd1 clkbuf_1_1__f__0390_.A a_2686_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7746 a_5704_17461# _0456_.B a_5632_17461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X7747 a_1735_29941# _0847_.A1 a_2073_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X7748 a_12794_4765# a_12355_4399# a_12709_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7749 a_12575_13647# a_11877_13653# a_12318_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7750 vccd1 _0954_.D a_14772_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.29 ps=1.58 w=1 l=0.15
X7751 a_20111_6031# a_19329_6037# a_20027_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7752 a_20613_6575# _0548_.A1 a_20267_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7753 a_6927_13103# _0745_.A2 a_6833_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7754 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7755 a_14875_18589# _1076_.Q a_14775_18589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X7756 vccd1 a_2623_9019# a_2539_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7757 a_25800_17289# a_25401_16917# a_25674_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7758 vccd1 a_27590_25183# a_27517_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7759 vccd1 a_15023_28887# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7760 _0983_.D a_21207_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7761 vssd1 _0931_.CLK a_18151_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7762 a_24949_17999# _0993_.D a_24867_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7763 a_25401_4949# a_25235_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7765 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_14260_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7766 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13616_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7768 a_2398_27613# a_1959_27247# a_2313_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7769 _0835_.A1 a_2626_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X7770 vssd1 a_10903_2491# a_10861_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7772 vccd1 _0931_.CLK a_20083_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7774 a_25401_14741# a_25235_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7775 a_8105_1685# a_7939_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7776 a_17581_3311# a_17415_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7777 vccd1 a_23174_7093# a_23101_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7778 a_27839_9117# a_27057_8751# a_27755_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7779 _0685_.B a_9284_10901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X7781 vccd1 _0746_.A2 a_6549_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X7783 a_15667_12559# _0667_.B1 a_15845_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7785 a_16109_14557# a_15575_14191# a_16014_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7786 a_5813_13647# _0780_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7787 _0752_.Y _0814_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7788 vssd1 _0866_.B a_12557_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7789 vccd1 _1033_.CLK a_26983_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7790 vccd1 a_20947_21263# a_21115_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7791 a_20387_17821# a_19605_17455# a_20303_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7792 _0515_.X a_19347_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X7793 vssd1 a_23637_12533# _0576_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X7794 a_12189_27001# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7796 a_25405_17455# _0926_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7797 a_23266_4511# a_23098_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7798 vssd1 a_22659_19631# _0999_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7799 a_17086_17999# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X7800 vccd1 a_25623_5755# a_25539_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7801 a_4999_23759# _0813_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X7804 a_17585_22895# _0932_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7805 vccd1 _0768_.B1 a_7111_13655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7807 vssd1 a_20947_21263# a_21115_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7808 vssd1 a_18758_20149# a_18716_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7809 _0502_.X a_12763_12879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7810 vccd1 _0994_.CLK a_22015_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7813 vccd1 a_11582_13077# _0524_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X7814 vssd1 a_6612_14709# _0795_.A2_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X7815 a_21150_4511# a_20982_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7817 a_22281_12265# _0658_.X a_22199_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7818 a_25125_2589# a_24591_2223# a_25030_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7822 a_18808_21641# a_18409_21269# a_18682_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7823 vccd1 a_22879_22351# a_23047_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7824 a_24949_17999# _0998_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7825 vccd1 _0959_.CLK a_9779_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7827 a_23381_26703# _0994_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7828 a_13817_12925# _0602_.A a_13735_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X7829 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7830 a_18271_6031# a_17489_6037# a_18187_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7833 a_11765_22325# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X7834 vssd1 a_17727_10383# a_17895_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7835 vssd1 a_22879_22351# a_23047_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7836 a_22181_16917# a_22015_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7837 _0959_.CLK a_10423_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7838 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7839 a_26869_22895# a_25879_22895# a_26743_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7840 _0664_.A2 a_21127_11809# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X7841 a_10325_10703# _0625_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7842 vssd1 _0699_.A0 a_4614_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
X7843 a_2313_3311# _0868_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7844 a_25497_12015# _0893_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7845 a_14287_13103# _1056_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7847 a_11233_14441# _0747_.B2 a_11149_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7850 a_13081_2473# _0555_.C1 a_12999_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7852 a_15278_2589# a_14839_2223# a_15193_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7853 a_8188_31055# a_7939_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7854 a_6937_27497# _0836_.Y a_7192_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7855 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7856 vccd1 _0444_.B _0752_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7857 temp1.capload\[2\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7858 _1063_.Q a_23047_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7859 a_11711_24527# _0444_.B _0825_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X7860 a_7691_3855# a_6909_3861# a_7607_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7861 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_9135_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7862 a_19942_9615# _1024_.Q a_19852_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X7863 a_4993_11471# _0807_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7864 vccd1 a_5417_20149# _0813_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7865 a_25769_19087# a_25235_19093# a_25674_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7866 _0917_.CLK a_9411_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7867 vccd1 _1053_.CLK a_14931_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7868 a_26670_20831# a_26502_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7872 vssd1 a_20303_17821# a_20471_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7873 vccd1 a_23415_19061# a_23331_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7874 vccd1 fanout24.A a_22015_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7875 a_15186_3677# a_14913_3311# a_15101_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7876 _0523_.B1 a_20393_8545# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X7877 _0634_.C1 a_19991_5056# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7878 vccd1 a_9339_7093# a_9255_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7879 _1052_.D a_17803_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7880 vccd1 a_2991_1403# a_2907_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7881 vssd1 _0814_.A2 a_1591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7882 a_21073_1999# _0946_.D a_20635_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7885 vssd1 a_5600_14165# _0736_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X7886 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7887 a_21407_3677# a_20543_3311# a_21150_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7888 vssd1 _0845_.B1 _0845_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7889 a_4790_2767# a_4517_2773# a_4705_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7890 vccd1 a_18611_14735# _0662_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7891 a_15538_27765# a_15370_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7893 a_2566_3423# a_2398_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7894 vccd1 a_15427_23439# a_15595_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7895 _0497_.B2 a_23047_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7896 a_9742_5599# a_9574_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7897 vssd1 _0644_.A2 a_15093_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7898 a_21258_19997# a_20985_19631# a_21173_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7899 a_17260_12265# _0533_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7901 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_12716_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7902 a_15787_2589# a_15005_2223# a_15703_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7903 vssd1 a_15427_23439# a_15595_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7904 a_18282_18793# _0577_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X7905 _0464_.X a_2051_14848# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7906 vccd1 _0917_.CLK a_14287_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7907 a_14744_6575# _0532_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X7908 vssd1 _0837_.A1 a_9636_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7909 _0579_.X a_17231_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7910 vssd1 _0999_.CLK a_22383_19093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7912 _1053_.D a_17251_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7913 a_24554_2741# a_24386_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7914 a_23101_7119# a_22567_7125# a_23006_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7915 a_4524_8751# _0695_.A1 a_4221_8725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7917 vccd1 a_25639_12559# a_25807_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7918 a_26317_13967# _1012_.D a_25971_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7919 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7920 a_12920_4399# a_12521_4399# a_12794_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7921 a_13989_6351# _1027_.Q a_13551_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7923 vccd1 a_11747_3677# a_11915_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7924 a_14621_8897# _0600_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7925 a_4889_4399# input3.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7926 vssd1 a_11815_12265# _0475_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7929 a_9666_8029# a_9393_7663# a_9581_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7930 vccd1 a_12743_13621# a_12659_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7931 a_27295_4765# a_26597_4399# a_27038_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7932 vssd1 a_25639_12559# a_25807_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7933 vccd1 _0445_.A a_7389_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X7934 vccd1 a_10459_13647# a_10627_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7935 vssd1 _0999_.CLK a_26983_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7938 a_15097_3855# a_14563_3861# a_15002_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7940 a_3298_17143# _0456_.A a_3512_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X7941 _0836_.Y _0845_.A2 a_1775_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7942 a_22457_12559# _0938_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7943 a_16347_21085# a_15483_20719# a_16090_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7944 vssd1 a_10459_13647# a_10627_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7945 vccd1 _0722_.A a_4167_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7946 a_8079_28500# _0820_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7947 vssd1 a_15611_3677# a_15779_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7948 a_25401_3861# a_25235_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7950 a_2953_26709# a_2787_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7951 a_14453_14557# _1075_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X7953 a_4238_3855# a_3799_3861# a_4153_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7954 a_2122_3855# a_1683_3861# a_2037_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7956 a_17802_14441# _0628_.X a_17722_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7957 vccd1 _0845_.C1 a_12629_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7958 _0651_.C a_20175_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7959 _0618_.B2 a_23415_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7960 vccd1 a_3270_2741# a_3183_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X7961 vssd1 _0553_.X a_15115_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X7963 a_12643_12559# _0836_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X7964 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7967 vccd1 _1079_.Q a_9411_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7968 a_23742_6031# a_23303_6037# a_23657_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7969 vccd1 _0847_.A2 a_10788_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7971 vssd1 a_2842_2741# a_2780_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X7972 vccd1 _1030_.CLK a_15667_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7973 a_22549_1135# a_22383_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7974 vccd1 _1033_.CLK a_25143_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7976 vssd1 a_11455_11195# a_11413_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7977 vccd1 a_26267_7093# a_26183_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7979 vssd1 a_25750_6005# a_25708_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7980 a_23818_21237# a_23650_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7981 a_7197_20969# _0866_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X7982 vssd1 _0821_.Y a_8583_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7983 a_15795_27791# a_14931_27797# a_15538_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7984 _1048_.D a_26267_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7985 a_4337_28335# _0847_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7987 a_25511_11471# _0664_.A2 a_25593_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7989 a_2686_15823# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X7990 _0995_.CLK a_9227_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X7991 vssd1 a_10198_7351# _0567_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7992 vccd1 a_20761_9633# _0506_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X7993 vccd1 _0861_.B1 a_3141_19148# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7995 _1061_.D a_19275_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7997 vccd1 _1078_.Q a_14453_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X7998 _0983_.D a_21207_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7999 vssd1 _0844_.B _0845_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8000 a_6735_11177# _0685_.X a_6653_10933# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8001 a_17078_12265# _0564_.X a_16829_12161# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8002 temp1.dcdc.A a_1674_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8003 a_4167_17999# _0722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8004 a_2723_4765# a_1941_4399# a_2639_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8005 vssd1 _0833_.A a_10814_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8006 a_22383_14848# _1048_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8007 a_23201_10089# _0488_.B2 a_23119_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8008 a_15465_27791# a_14931_27797# a_15370_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8009 a_5341_3145# a_4351_2773# a_5215_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8011 a_15404_2223# a_15005_2223# a_15278_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8013 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8014 _0643_.X a_22291_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X8015 vccd1 temp1.capload\[6\].cap_51.LO temp1.capload\[6\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8017 vssd1 a_2114_1653# _0860_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X8019 a_4244_25071# a_4213_25223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X8020 _0854_.B _0850_.Y a_12342_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X8021 a_12437_8751# _0582_.A a_12355_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X8022 vssd1 a_5015_2491# a_4973_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8023 vccd1 a_25474_6687# a_25401_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8024 a_25309_9295# _1066_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8026 a_25750_9951# a_25582_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8027 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8028 a_10459_13647# a_9595_13653# a_10202_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8029 a_12318_6005# a_12150_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8030 a_2398_27613# a_2125_27247# a_2313_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8031 _0873_.Y _0872_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8035 a_25915_9117# a_25217_8751# a_25658_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8036 a_5089_14851# _0722_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8038 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_7295_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8039 _1076_.Q a_2991_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8040 vssd1 _0975_.CLK a_24591_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8042 a_10229_14735# _0770_.B1 a_10313_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8043 vccd1 _0662_.A3 a_22383_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8044 a_20755_8029# a_19973_7663# a_20671_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8045 a_18298_11445# a_18130_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8046 a_15277_9839# a_14287_9839# a_15151_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8047 a_18001_12043# _0504_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8048 a_4251_11249# _0698_.A2_N a_4250_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X8049 a_3138_1679# a_2885_2057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.178875 ps=1.26 w=0.42 l=0.15
X8050 a_10412_7119# _0566_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X8051 a_12383_10205# a_11601_9839# a_12299_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8052 a_23457_12015# _1000_.Q a_23385_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8056 a_10335_7439# _0566_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8058 a_27847_22173# a_26983_21807# a_27590_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8059 a_11344_19631# _0837_.A1 a_11238_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X8060 a_16802_15529# _0579_.X a_16553_15425# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8061 _0663_.X a_23579_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X8062 a_18279_3677# a_17415_3311# a_18022_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8063 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_3983_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8064 a_25129_23439# _0995_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8065 a_18130_11471# a_17857_11477# a_18045_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8066 a_5294_23759# _0809_.B2 a_4999_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X8067 _0996_.Q a_25807_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8068 a_21610_13215# a_21442_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8069 a_3735_26703# a_2953_26709# a_3651_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8070 vssd1 a_8971_4917# a_8929_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8071 a_23649_10703# _0621_.A1 a_23303_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8072 a_20204_18793# _0584_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X8073 a_12065_11471# _0580_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8074 a_7896_11703# _0567_.A1 a_8038_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8076 vssd1 a_21867_13469# a_22035_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8077 _0747_.B2 _0735_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X8078 vccd1 a_3155_21271# _0809_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8079 a_19613_16617# _0522_.B1 a_19697_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8081 temp1.inv1_1.Y temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8082 _0996_.Q a_25807_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8083 _0694_.A2 _0657_.X a_7271_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8084 a_27517_17821# a_26983_17455# a_27422_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8085 a_25539_4765# a_24757_4399# a_25455_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8087 a_11269_16367# a_11068_16617# _0882_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8088 a_15461_18377# a_14471_18005# a_15335_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8089 vssd1 a_23047_15797# a_23005_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8090 vccd1 a_17251_26427# a_17167_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8093 vssd1 _1075_.Q a_7939_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X8094 a_27931_16733# a_27149_16367# a_27847_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8095 a_26133_3311# a_25143_3311# a_26007_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8096 a_19191_21263# a_18409_21269# a_19107_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8097 a_9305_16672# _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8098 vccd1 _0845_.A2 a_7192_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8099 a_6427_11989# _0758_.A1 a_6858_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X8100 a_6971_29245# _0825_.A0 a_6608_29111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8104 a_17727_10383# a_16863_10389# a_17470_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8106 _0650_.X a_25511_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8107 vccd1 a_27739_6843# a_27655_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8110 vccd1 a_9043_12567# _0807_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8112 a_10018_4511# a_9850_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8113 vssd1 _0582_.C a_20697_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8114 _0843_.Y _0843_.B a_1775_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8115 vccd1 a_14341_17429# _0773_.A2_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8117 a_22361_5487# _1008_.Q a_22015_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8118 a_4439_24233# _0774_.A2 io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8119 a_18114_1247# a_17946_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8120 a_18681_8751# _0897_.D a_18243_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8122 vccd1 a_4847_1501# a_5015_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8123 a_2248_4233# a_1849_3861# a_2122_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8124 a_27698_4943# a_27521_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8125 a_4793_4949# a_4627_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8126 a_5074_12559# _0756_.A2 a_4771_12791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X8127 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8129 a_4364_4233# a_3965_3861# a_4238_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8130 _0584_.B1 a_22015_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8131 vccd1 _0807_.B a_3713_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8132 a_12189_27001# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X8133 a_4422_1501# a_4149_1135# a_4337_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8134 a_4974_4765# a_4535_4399# a_4889_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8135 a_15921_2057# a_14931_1685# a_15795_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8136 a_18114_1247# a_17946_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8138 a_4441_29423# _0845_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8139 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8140 vssd1 _0471_.X a_13035_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X8141 vccd1 temp1.capload\[13\].cap.A temp1.capload\[13\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8142 a_17397_10383# a_16863_10389# a_17302_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8144 vccd1 fanout10.A a_11803_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8145 a_23868_6409# a_23469_6037# a_23742_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8146 a_5817_6351# _0689_.X a_5599_6263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X8147 a_14894_7775# a_14726_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8148 a_2122_12015# a_1945_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8149 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15088_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8150 vssd1 a_12610_21807# a_12716_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8151 vssd1 _1060_.D a_19536_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X8152 vssd1 a_18298_11445# a_18256_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8154 a_27847_2589# a_27149_2223# a_27590_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8155 a_15921_7235# _0634_.X a_15848_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X8156 _0892_.D a_25623_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8157 vccd1 _1033_.CLK a_24591_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8158 _0764_.A1 a_4170_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X8159 a_7326_22057# _0866_.B a_7244_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8160 a_12701_8585# a_11711_8213# a_12575_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8161 a_14894_7775# a_14726_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8162 _0992_.D a_21943_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8163 vccd1 a_2991_2491# _0837_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8164 vssd1 _0827_.A a_11269_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8165 a_25581_16367# a_24591_16367# a_25455_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8166 a_27422_22173# a_27149_21807# a_27337_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8167 vccd1 a_15538_27765# a_15465_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8168 a_2833_24759# _0844_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8169 a_27422_8029# a_27149_7663# a_27337_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8170 a_21426_8863# a_21258_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8172 vssd1 _0644_.X _0684_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8173 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X8174 a_25401_6941# a_24867_6575# a_25306_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8175 vssd1 _0845_.A2 _0833_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8176 vccd1 _0872_.A1 a_5639_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8178 a_4517_2589# a_3983_2223# a_4422_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8179 vssd1 _0908_.CLK a_7203_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8180 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8181 vssd1 a_14599_19087# a_14767_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8182 vccd1 _0975_.CLK a_22015_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8183 vccd1 _0444_.A a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8184 a_26225_15113# a_25235_14741# a_26099_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8185 a_19602_6031# a_19329_6037# a_19517_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8186 a_25593_11471# _0650_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8187 a_10567_19061# _0761_.B a_10785_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X8188 a_1757_5487# a_1591_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8189 vssd1 a_25731_6941# a_25899_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8190 vccd1 a_23139_2741# a_23055_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8191 a_10091_8029# a_9393_7663# a_9834_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8193 vccd1 a_8859_17999# _0472_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8194 vssd1 a_15446_2335# a_15404_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8195 _0650_.A1 a_28015_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8196 vccd1 a_26467_26525# a_26635_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8198 vccd1 a_17819_1679# a_17987_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8199 a_1849_3861# a_1683_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8200 vssd1 _0694_.A1 a_4852_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8203 a_3965_3861# a_3799_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8204 vssd1 _0524_.X a_12565_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8205 a_19846_9295# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X8206 _1015_.CLK a_23763_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8207 vccd1 _0893_.CLK a_24683_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8208 a_5813_25117# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8210 _0548_.A1 a_26175_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8211 _0990_.D a_12375_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8212 vccd1 a_15354_3423# a_15281_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8213 vccd1 a_27847_25437# a_28015_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8216 a_9022_3855# a_8749_3861# a_8937_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8217 vccd1 a_26911_23163# a_26827_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8218 a_24811_2767# a_23947_2773# a_24554_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8219 a_2291_29967# _0847_.B1 a_1975_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X8220 a_15391_8323# _0675_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8221 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8222 a_4590_28447# a_4422_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8224 a_18320_8207# _0565_.B1 a_18065_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X8225 vccd1 _0860_.B _0856_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8228 vccd1 a_21575_3579# a_21491_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8229 vccd1 a_2842_2741# a_2776_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X8232 a_17857_15529# _0932_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8234 a_8021_18793# _0459_.X a_8105_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8237 vccd1 a_2752_1897# a_2762_1801# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8239 _0882_.A2 _0880_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8240 a_21150_3423# a_20982_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8241 a_13771_10383# a_12907_10389# a_13514_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8242 a_20598_22325# a_20430_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8243 a_5537_6575# _0686_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8245 vccd1 a_2639_4765# a_2807_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8246 vssd1 a_24554_2741# a_24512_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8248 vccd1 _0466_.A _0794_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8249 a_26417_20719# _0966_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8250 vssd1 _0491_.X a_15196_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X8251 a_25582_3677# a_25309_3311# a_25497_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8253 a_14920_1135# _0954_.D _0642_.D_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.19175 ps=1.24 w=0.65 l=0.15
X8254 a_23005_11791# _0505_.A1 a_22659_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8255 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8257 vssd1 _0664_.A2 a_20981_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8258 a_17612_17455# a_17213_17455# a_17486_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8259 a_12525_27791# a_12348_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8261 vccd1 _0809_.B2 a_4769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8262 a_2962_14735# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8263 a_15611_14735# a_14747_14741# a_15354_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8264 a_13441_10383# a_12907_10389# a_13346_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8265 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8267 vssd1 a_25842_4917# a_25800_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8268 vccd1 a_27847_8029# a_28015_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8269 vssd1 _0745_.A1 a_6600_11587# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8270 vccd1 _0764_.A1 a_5626_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X8271 vccd1 _0689_.X a_6749_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8273 a_21647_7663# _0516_.B1 a_21825_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X8274 a_21169_23983# a_21003_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8275 a_15630_16479# a_15462_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8277 vccd1 a_9834_7775# a_9761_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8278 a_6368_29423# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8280 fanout10.A a_11619_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8281 vccd1 temp1.capload\[12\].cap_42.LO temp1.capload\[12\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8283 a_24591_11177# _0664_.A2 a_24673_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8284 vssd1 ANTENNA_7.DIODE a_25707_25321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X8285 vccd1 a_12575_6031# a_12743_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8286 vssd1 a_15887_16733# a_16055_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8287 _0893_.D a_26267_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8288 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8289 a_17796_22895# a_17397_22895# a_17670_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8290 a_15281_14735# a_14747_14741# a_15186_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8291 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X8292 vccd1 _0964_.CLK a_25235_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8294 vccd1 _0521_.A a_13367_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8296 _1014_.Q a_28015_12283# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8300 a_10083_5853# a_9301_5487# a_9999_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8301 vssd1 a_20195_26677# a_20153_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8302 vccd1 _1078_.Q a_14563_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8303 a_22737_3311# _0632_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8304 a_15483_11177# _0614_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X8305 a_21361_6825# _1006_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8306 a_19659_13647# a_18961_13653# a_19402_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8307 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11244_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8309 vccd1 a_26099_15823# a_26267_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8310 a_19234_13647# a_18795_13653# a_19149_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8311 a_25539_16733# a_24757_16367# a_25455_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8312 vssd1 _0975_.CLK a_22107_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8313 a_22291_12559# _0563_.B1 a_22469_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X8314 vccd1 a_14342_19061# a_14269_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8316 vccd1 a_9503_19087# _0471_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8317 vssd1 _0798_.A2 a_7939_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8318 vccd1 _0579_.C a_17909_16395# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8319 _0783_.A1 _0778_.Y a_5813_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8320 _0788_.C _0809_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8321 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8322 a_17302_2767# a_17029_2773# a_17217_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8323 a_10386_4917# a_10218_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8324 _0746_.A2 _0678_.Y a_8033_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8325 vccd1 a_26175_12283# a_26091_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8326 a_23377_21269# a_23211_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8327 a_3057_17705# a_2869_17501# a_2975_17461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8328 a_12885_4233# a_11895_3861# a_12759_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8329 vccd1 a_8270_21237# a_8197_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8330 _0771_.C1 a_10147_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X8331 vssd1 _0594_.C a_18427_2473# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8332 a_16523_4765# a_15741_4399# a_16439_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8333 a_7277_3855# a_6743_3861# a_7182_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8334 _0814_.A2 a_3891_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8335 a_7832_10927# a_7801_11079# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X8336 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8767_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8337 _1019_.CLK a_15667_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8338 _0545_.B2 a_14011_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X8339 vssd1 a_11803_23439# _0444_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8340 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9319_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8341 a_27847_3677# a_26983_3311# a_27590_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8342 a_25405_7663# _0621_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8346 a_9573_4233# a_8583_3861# a_9447_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8347 a_1766_29423# temp1.inv1_1.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8348 a_23005_22729# a_22015_22357# a_22879_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8349 vssd1 a_2547_3855# a_2715_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8350 a_25769_10383# a_25235_10389# a_25674_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8351 _0975_.CLK a_22015_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8352 a_15281_3677# a_14747_3311# a_15186_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8353 a_17903_1679# a_17121_1685# a_17819_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8354 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8356 a_5060_31055# a_4811_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8357 a_20349_6575# _0548_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8358 vccd1 _0643_.B1 a_27249_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8359 a_7544_30761# a_7295_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8361 a_7461_6037# a_7295_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8362 a_25497_6031# _0506_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8363 _1046_.D a_23599_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8365 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8366 a_23975_26703# a_23193_26709# a_23891_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8367 vssd1 a_10183_9295# a_10351_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8368 a_2616_28335# a_2217_28335# a_2490_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8369 a_22185_26159# _1019_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8371 a_1775_31375# _0444_.A _0444_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8372 _0725_.A a_3983_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8373 _0565_.B1 _0474_.X a_14655_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8374 vssd1 a_25455_16733# a_25623_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8376 vssd1 _0917_.CLK a_14287_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8377 vssd1 a_12999_31055# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8378 vccd1 a_9919_6740# _1084_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8379 a_21258_19997# a_20819_19631# a_21173_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8381 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8382 a_8944_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8383 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9016_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8384 vssd1 io_in[0] a_2962_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8385 a_3559_4943# a_2695_4949# a_3302_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8386 vccd1 a_23637_12533# _0576_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8387 a_17209_26159# a_16219_26159# a_17083_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8389 a_25490_8029# a_25051_7663# a_25405_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8391 a_16347_21085# a_15649_20719# a_16090_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8392 a_14821_12381# a_14287_12015# a_14726_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8393 vssd1 _0959_.CLK a_9871_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8394 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8395 vssd1 a_4403_25589# _0840_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8396 a_4324_14197# _0456_.B a_4252_14197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X8397 a_15759_9001# _0595_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X8398 _0506_.A2 a_20761_9633# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X8399 a_22914_21085# a_22641_20719# a_22829_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8400 a_21257_1135# _1034_.Q a_20911_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8401 a_23373_1135# a_22383_1135# a_23247_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8403 a_9761_8029# a_9227_7663# a_9666_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8404 a_27337_23983# _0928_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8405 vccd1 a_13514_10357# a_13441_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8406 vssd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_2686_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8408 vccd1 _1015_.CLK a_26983_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8409 vccd1 a_12207_21085# a_12375_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8410 vccd1 a_18447_3579# a_18363_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8411 a_5399_4765# a_4701_4399# a_5142_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8412 vccd1 temp1.capload\[8\].cap.A temp1.capload\[8\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8414 a_26099_15823# a_25235_15829# a_25842_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8415 vccd1 _0725_.A a_3891_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X8416 vssd1 a_26099_4943# a_26267_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8417 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8418 a_15078_17973# a_14910_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8419 vssd1 a_5015_28603# a_4973_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8420 _0865_.Y a_12356_19203# a_12557_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8421 a_18022_3423# a_17854_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8423 a_9853_6037# a_9687_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8424 a_17125_19631# _1050_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8425 vccd1 a_15354_14709# a_15281_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8426 vssd1 _1015_.CLK a_25235_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8427 _0494_.X a_14637_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X8428 _1078_.D _0840_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8429 _0833_.Y _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8430 a_19517_26703# _1018_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8431 vssd1 a_5199_1653# a_5157_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8432 a_8393_12015# _0654_.Y a_8175_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X8433 a_20939_22351# a_20157_22357# a_20855_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8435 _0680_.Y _0685_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8436 vssd1 _0443_.A a_11803_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X8437 vccd1 a_13939_22325# a_13855_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8438 vssd1 a_25842_3829# a_25800_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8441 a_26091_6031# a_25309_6037# a_26007_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8442 a_18505_20175# _1049_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8443 a_20897_3311# _1040_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8444 a_7469_28585# _0821_.B _0821_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8446 _0922_.CLK a_4259_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8447 a_15937_9001# _0589_.X a_15841_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X8448 vssd1 _0511_.D a_10667_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X8449 vccd1 a_24462_22325# a_24389_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8452 _0618_.B2 a_23415_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8455 vccd1 a_22162_21919# a_22089_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8456 vccd1 temp1.inv1_1.Y a_1766_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8457 a_26225_19631# a_25235_19631# a_26099_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8458 vccd1 _0893_.CLK a_25235_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8459 a_12061_3861# a_11895_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8461 vssd1 a_26175_3579# a_26133_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8462 a_2309_4765# a_1775_4399# a_2214_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8463 vssd1 _0797_.A1 a_14644_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8464 a_12801_2767# _0946_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8465 vccd1 a_4590_1247# a_4517_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8466 a_15661_32463# temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8467 vccd1 a_19827_13621# a_19743_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8468 a_20153_27081# a_19163_26709# a_20027_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8469 a_22369_15823# _0925_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8470 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8473 a_22162_21919# a_21994_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8474 _0678_.Y _0546_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8475 a_18961_13653# a_18795_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8476 vssd1 a_2639_4765# a_2807_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8477 vccd1 _1028_.CLK a_14287_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8478 a_25143_9295# _0506_.A2 a_25321_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X8479 a_2405_12015# a_2228_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8480 vccd1 _0644_.A2 a_15833_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8481 _0727_.A1 a_7939_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X8482 _0575_.B a_25623_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8483 a_11505_14191# _0860_.A a_11067_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8484 vssd1 _0845_.A2 a_7385_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8485 vccd1 _0504_.A a_18059_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8486 a_14637_18005# a_14471_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8488 a_10819_2589# a_10037_2223# a_10735_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8489 vccd1 a_5015_26427# a_4931_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8490 vccd1 _0471_.X a_14559_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8491 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5060_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8493 vssd1 a_27847_8029# a_28015_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8495 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8496 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_7544_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8497 a_14188_27023# _0815_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8501 vccd1 a_27590_7775# a_27517_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8502 vssd1 _0494_.X a_20111_10955# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8504 a_27249_10383# _0893_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8506 vccd1 _0825_.S temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8507 a_20893_27247# a_20727_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8508 a_14341_15797# _0798_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X8509 vccd1 _0710_.A2 a_5445_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X8510 a_9911_12061# _0836_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8511 _0549_.B2 a_8971_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8512 vccd1 a_19770_6005# a_19697_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8513 a_9495_11249# _0597_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.335 w=0.64 l=0.15
X8514 vssd1 _0583_.C a_19281_18337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8515 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_13912_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8516 vssd1 a_8325_11769# a_8259_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X8517 a_12207_18909# a_11509_18543# a_11950_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8518 _1063_.Q a_23047_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8519 a_11877_6037# a_11711_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8521 a_27847_22173# a_27149_21807# a_27590_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8523 a_14483_15279# _1076_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X8524 a_6937_27497# _0845_.C1 _0837_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8525 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8526 a_12805_3561# _0586_.B2 a_12723_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8527 a_10275_4765# a_9411_4399# a_10018_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8528 a_25121_14025# a_24131_13653# a_24995_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8529 vccd1 _0964_.CLK a_22015_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8531 a_18597_21263# _1060_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8532 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8534 a_18025_7809# _0633_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X8535 vssd1 a_15319_10107# a_15277_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8536 a_3394_26677# a_3226_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8537 vssd1 _0475_.X a_10325_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X8538 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8539 a_4993_11471# _0708_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X8540 vccd1 _0602_.A a_14287_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8541 vssd1 a_14729_16911# _0582_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X8542 a_11149_14441# _0717_.A2 a_11067_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8544 vssd1 _0662_.X a_23579_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8545 a_6704_13077# _0768_.A1 a_6833_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8546 _0752_.Y _0444_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8547 a_22365_12265# _0939_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8548 vccd1 a_14894_12127# a_14821_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8549 vccd1 a_25455_22173# a_25623_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8550 vccd1 a_22879_16911# a_23047_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8551 a_15975_10721# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8552 a_2205_15101# _0456_.B a_2133_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8554 a_7928_15055# _0445_.A a_7625_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X8555 vssd1 _0512_.X a_18497_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X8556 a_27337_17455# _0927_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8557 a_23385_16367# _0929_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8558 vccd1 a_9003_15797# _0636_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X8559 a_4333_1685# a_4167_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8560 a_5177_27023# _0845_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8561 vssd1 _0845_.C1 _0845_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8563 _0551_.C1 a_20911_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X8564 a_25217_8751# a_25051_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8565 a_15193_2223# _0945_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8566 a_20157_22357# a_19991_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8567 a_14967_20175# a_14103_20181# a_14710_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8568 a_9761_13653# a_9595_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8569 a_25616_7663# a_25217_7663# a_25490_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8571 _1069_.Q a_26175_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8572 a_12242_27791# a_12065_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8573 vssd1 a_15812_6005# _0675_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8576 a_1591_21807# _0753_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8577 vccd1 _0491_.X a_17489_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8578 a_16940_11177# _0616_.B1 a_16685_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X8580 a_18141_17277# _0504_.A a_18059_17024# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8581 vccd1 _1030_.CLK a_20543_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8582 vccd1 a_13459_8751# _0521_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8583 a_17394_1679# a_16955_1685# a_17309_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8584 vccd1 a_13551_8215# _0582_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8585 a_27973_25071# a_26983_25071# a_27847_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8587 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8588 a_18088_13647# _0522_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X8589 a_19199_25615# a_18501_25621# a_18942_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8590 a_22622_1653# a_22454_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8591 a_20180_9615# _0533_.X a_19689_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X8593 a_22817_18517# _0662_.A1 a_23070_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X8595 a_14637_20175# a_14103_20181# a_14542_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8596 vccd1 a_17909_16395# _0648_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X8597 vccd1 a_25750_3423# a_25677_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8598 a_23201_9839# _0488_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8599 vssd1 _0532_.A2 a_11965_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X8601 a_15005_2223# a_14839_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8602 a_16826_26271# a_16658_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8604 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8605 a_25401_21269# a_25235_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8606 a_9636_20969# _0761_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8607 a_12333_20719# a_11343_20719# a_12207_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8608 vssd1 _0694_.A2 a_5510_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X8609 a_17086_17999# _0920_.D a_16929_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8610 vccd1 a_3270_2741# _0850_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X8611 a_6072_25077# _0445_.A a_6000_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X8612 vccd1 _0471_.X a_10791_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8613 a_2581_5487# a_1591_5487# a_2455_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8614 a_17861_10927# _0565_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8616 vssd1 a_21345_15253# _0542_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8617 vssd1 a_26267_14709# a_26225_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8619 a_7331_6941# a_6467_6575# a_7074_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8620 _0845_.C1 a_4811_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8621 a_9326_25398# _0816_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8622 a_24301_2767# _1034_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8623 vssd1 _0959_.CLK a_14839_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8624 a_26007_6031# a_25309_6037# a_25750_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8625 a_17041_7439# _0897_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X8626 a_19878_17821# a_19439_17455# a_19793_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8627 vccd1 a_7073_20149# _0789_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8629 a_6600_26409# _0819_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8630 a_2585_25621# a_2419_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8631 fanout9.A fanout11.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8632 a_21775_18909# a_21077_18543# a_21518_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8633 a_10125_1135# a_9135_1135# a_9999_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8635 vssd1 _0491_.X a_12333_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8636 vssd1 _0670_.A2 a_13437_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X8637 vssd1 _0483_.X a_20847_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8638 a_17213_17455# a_17047_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8639 a_22737_14191# _0939_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8640 a_25589_4943# _0531_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8641 a_25401_25621# a_25235_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8642 vssd1 _0917_.CLK a_11711_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8643 vssd1 a_11435_8751# _0842_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8644 _1077_.Q a_3083_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8645 a_10089_10089# _0545_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8646 a_23487_6825# _0619_.B1 a_23569_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8648 a_22990_1247# a_22822_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8649 vssd1 a_2455_6031# a_2623_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8650 a_17769_3311# _1041_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8651 vssd1 _0847_.B1 a_1735_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X8652 _0917_.D a_12743_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8653 a_18148_10089# _0624_.C a_18053_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X8655 a_17811_3855# a_17029_3861# a_17727_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8656 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8657 a_6463_7913# _0681_.X a_6376_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8659 vccd1 a_17470_2741# a_17397_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8660 vccd1 _0444_.A a_2787_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8664 a_21831_10089# _0666_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X8665 a_24462_20149# a_24294_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8667 vssd1 a_2991_2491# _0837_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8668 a_19970_2767# a_19531_2773# a_19885_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8669 a_7192_27497# _0837_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8671 a_12575_8207# a_11711_8213# a_12318_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8672 _0758_.A2 _0713_.A1 a_5639_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8674 a_12425_9839# a_11435_9839# a_12299_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8676 _0761_.X a_9636_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8677 _1024_.Q a_21851_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8678 a_7260_14441# _0778_.B1 a_6795_14343# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8679 vccd1 _0487_.X a_18409_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8680 vccd1 _1019_.CLK a_18243_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8681 vssd1 _0583_.C a_20237_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8683 a_25842_19743# a_25674_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8685 vssd1 a_18001_12043# _0667_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X8686 vccd1 _0845_.A1 a_7326_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X8687 a_24294_20175# a_24021_20181# a_24209_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8688 a_8116_10383# _0679_.A2 _0746_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X8689 _0582_.A a_13551_8215# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8690 vccd1 _0445_.A a_9811_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8691 a_17783_12672# _1026_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8692 vssd1 a_26099_19997# a_26267_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8693 _0740_.X a_6600_26409# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8694 a_27590_3423# a_27422_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8695 vccd1 _0614_.X a_18221_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8696 a_10988_10927# a_10589_10927# a_10862_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8697 vccd1 clkbuf_1_1__f__0390_.A a_2686_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8698 vccd1 a_19107_21263# a_19275_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8699 a_2539_6031# a_1757_6037# a_2455_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8700 vssd1 _0523_.B1 a_20521_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8701 a_16305_31599# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8702 vccd1 _0827_.A a_7469_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8704 vssd1 _0722_.B a_3028_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8705 _0905_.Q a_5383_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8707 vssd1 a_17928_8181# _0587_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8709 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8710 vssd1 a_19107_21263# a_19275_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8711 vssd1 a_27590_16479# a_27548_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8712 a_9945_4949# a_9779_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8713 a_15151_8029# a_14287_7663# a_14894_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8714 _0861_.B1 a_3799_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8715 a_2882_24527# a_2833_24759# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X8716 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8717 a_25674_1501# a_25401_1135# a_25589_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8718 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X8719 a_9574_1501# a_9301_1135# a_9489_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8722 a_21683_9117# a_20819_8751# a_21426_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8723 _0639_.B a_13479_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8724 a_6612_8181# _0686_.A a_7004_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X8726 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8727 a_22751_17455# _0994_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8730 _0583_.C a_14603_18589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X8731 a_22963_22351# a_22181_22357# a_22879_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8732 a_18354_7913# _0634_.C1 a_18274_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8734 vccd1 _0529_.Y a_22015_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8735 a_6611_25589# _0789_.B1 a_6809_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8736 _0483_.X a_15115_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X8737 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8739 vccd1 a_3727_4917# a_3643_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8740 a_24811_2767# a_24113_2773# a_24554_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8742 a_25030_22173# a_24591_21807# a_24945_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8744 _0584_.A2 a_15607_15307# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X8745 a_13629_4943# _0670_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8746 a_7649_6031# _0611_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8747 vssd1 a_25658_7775# a_25616_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8748 _0472_.X a_8859_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8749 a_25582_12381# a_25143_12015# a_25497_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8750 a_23966_12559# _0574_.X a_23886_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8751 a_17635_19997# a_16937_19631# a_17378_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8752 vssd1 a_17725_15073# _0487_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X8753 a_17520_2057# a_17121_1685# a_17394_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8754 a_2217_28335# a_2051_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8755 a_7810_4511# a_7642_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8756 a_3132_2045# a_2885_2057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.1493 ps=1.22 w=0.42 l=0.15
X8757 vssd1 _0651_.X _0684_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8758 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10791_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8759 a_24075_21263# a_23377_21269# a_23818_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8760 a_12532_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8761 a_6779_2589# a_6081_2223# a_6522_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8762 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_7387_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8763 vssd1 _0564_.C a_20819_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8766 a_27167_11471# _0619_.B1 a_27249_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8769 a_26233_22895# _0996_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8770 vccd1 _0734_.A2 _0696_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8771 vssd1 a_3523_13655# _0768_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8772 a_12299_10205# a_11435_9839# a_12042_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8773 vccd1 a_20303_17821# a_20471_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8774 vccd1 _0574_.C a_22751_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8775 vccd1 _0972_.CLK a_17415_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8776 a_18501_25621# a_18335_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8777 a_9184_25223# _0825_.A0 a_9326_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8778 a_17762_6031# a_17323_6037# a_17677_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8779 a_22914_21085# a_22475_20719# a_22829_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8780 a_4847_26525# a_4149_26159# a_4590_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8782 vccd1 a_25639_23439# a_25807_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8784 a_27590_17567# a_27422_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8785 a_7902_6005# a_7734_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8786 a_24294_20175# a_23855_20181# a_24209_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8787 vssd1 a_19770_6005# a_19728_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8789 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8790 a_22549_19093# a_22383_19093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8791 vccd1 _0934_.Q a_20204_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8792 _0666_.B a_20635_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X8793 a_16109_4765# a_15575_4399# a_16014_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8794 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9568_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8795 vssd1 a_11764_20149# _0858_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X8796 vssd1 a_25639_23439# a_25807_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8797 a_19697_16617# _0920_.Q a_19613_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8798 a_24757_4399# a_24591_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8799 vccd1 _0972_.CLK a_16863_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8800 vssd1 _0460_.C a_4137_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8802 a_14917_3855# _0954_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8803 vssd1 _1028_.CLK a_9227_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8804 a_2039_9295# a_1757_9301# a_1945_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X8805 _0583_.X a_20083_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8806 vssd1 a_9983_16885# a_9941_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8807 vssd1 a_9411_8751# _0917_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8808 a_19107_21263# a_18243_21269# a_18850_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8809 a_27847_16733# a_26983_16367# a_27590_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8810 a_12161_7119# _0636_.X a_12079_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8811 a_19517_3855# _0969_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8812 a_20614_5853# a_20175_5487# a_20529_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8813 a_4439_24233# _0774_.A2 io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8816 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8817 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8818 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8819 vccd1 _0850_.A _0850_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8820 _1053_.D a_17251_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8822 a_17489_1679# a_16955_1685# a_17394_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8823 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8825 a_21426_8863# a_21258_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8827 a_25658_8863# a_25490_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8828 a_4441_29423# _0845_.A1 _0845_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8830 a_6559_16911# _0472_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8831 vssd1 a_15611_14735# a_15779_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8832 a_4772_13621# _0768_.A1 a_4901_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8833 a_25589_3855# _1072_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8834 a_6809_25615# _0809_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X8835 a_23634_26677# a_23466_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8836 vssd1 a_19183_20149# a_19141_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8837 vssd1 a_20471_15547# a_20429_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8838 _1008_.Q a_28015_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8839 a_5796_31849# a_5547_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8840 a_18125_18517# _0662_.A1 a_18378_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X8841 vccd1 _0893_.CLK a_24131_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8842 vccd1 a_10147_15529# _0474_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X8843 a_19877_4399# _0497_.A1 a_19439_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8845 a_15369_9295# _0644_.X a_15115_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8848 _0659_.X a_22199_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X8849 vssd1 fanout10.A a_12355_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8850 a_10331_17999# _0749_.B1 a_10509_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X8851 a_19785_2057# a_18795_1685# a_19659_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8853 a_23097_10927# _0506_.A1 a_22659_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8854 _0737_.X a_8256_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8855 a_14603_18589# _1076_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8857 a_8355_11510# _0567_.A1 a_7896_11703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8858 vccd1 a_10091_8029# a_10259_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8859 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8860 a_6087_10927# _0707_.A1 _0708_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X8861 a_2198_5599# a_2030_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8862 vccd1 a_7499_6843# a_7415_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8863 a_7477_17999# _0737_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X8864 a_7515_5853# a_6817_5487# a_7258_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8865 a_2686_28879# clkbuf_1_1__f__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8866 a_22181_22357# a_22015_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8867 a_13261_22351# _1054_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8868 a_2398_3677# a_2125_3311# a_2313_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8869 a_8545_14709# _0546_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X8870 a_11877_13653# a_11711_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8872 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8873 _1035_.Q a_24979_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8877 vssd1 _0585_.X a_15759_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8878 a_14641_12015# _0897_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8881 _0808_.A a_6559_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8882 vccd1 _0845_.C1 a_9305_16672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X8884 vccd1 a_8859_17999# _0472_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8885 a_15841_1135# _1042_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8886 _0833_.Y _0845_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8887 a_13254_9295# a_12981_9301# a_13169_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8888 vccd1 _0523_.B1 a_19605_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8889 a_25582_12381# a_25309_12015# a_25497_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8890 vccd1 _0768_.A1 a_9497_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X8891 vccd1 a_10443_4667# a_10359_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8892 a_11913_13336# _0511_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X8893 a_6645_18543# _0795_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X8894 a_27149_14191# a_26983_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8895 vccd1 a_18539_1403# a_18455_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8896 a_3226_26703# a_2953_26709# a_3141_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8898 vssd1 a_10351_9269# a_10309_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8899 a_5621_3311# a_5455_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8900 a_26467_26525# a_25769_26159# a_26210_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8901 vssd1 a_15905_25589# _0861_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X8902 vccd1 a_4035_25045# _0843_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X8903 a_23910_9269# a_23742_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8904 a_27422_16733# a_27149_16367# a_27337_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8905 a_12042_9951# a_11874_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8906 vssd1 a_23615_8207# a_23783_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8907 a_19878_17821# a_19605_17455# a_19793_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8908 _0679_.A2 _0466_.A a_7663_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8909 vssd1 a_12207_15645# a_12375_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8910 vssd1 a_22325_6603# _0619_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X8911 a_20717_10383# _0531_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8912 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8915 vssd1 a_25842_16885# a_25800_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8916 vssd1 a_20977_10901# _0496_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8917 _0654_.Y _0662_.A1 a_8485_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8918 a_15369_11791# _0588_.A1 a_15023_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8919 _0856_.Y _0860_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8920 a_10218_2767# a_9945_2773# a_10133_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8921 a_7369_4399# a_7203_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8923 a_10103_26486# _0825_.A1 a_9644_26311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8924 vccd1 _1028_.CLK a_9687_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8925 _0535_.X a_12355_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X8926 a_12557_19407# _0866_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8929 a_22825_8751# a_22659_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8930 a_24738_13621# a_24570_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8931 vssd1 a_2455_9295# a_2626_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8932 vssd1 _0512_.A _0565_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8933 a_2823_27613# a_2125_27247# a_2566_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8934 a_27422_2589# a_26983_2223# a_27337_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8935 a_26965_4765# a_26431_4399# a_26870_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8936 a_11609_6825# _0522_.B1 a_11693_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8937 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8938 vccd1 _0546_.A2 a_8205_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8939 vccd1 a_9135_6575# _1028_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8940 a_10084_9839# _0475_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8941 a_25616_17455# a_25217_17455# a_25490_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8944 a_26601_18543# _1067_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8945 a_19329_3861# a_19163_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8946 a_17888_6409# a_17489_6037# a_17762_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8947 a_10876_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8948 a_20102_18793# _0584_.C1 a_20022_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8949 vccd1 a_21279_22895# _0994_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8950 _0794_.A3 _0768_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8951 vssd1 a_4847_2589# a_5015_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8952 _0631_.B a_22311_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8953 vccd1 a_5599_6263# _0694_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X8954 _0666_.D a_25143_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X8956 a_3183_2767# a_2401_2773# a_3099_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X8957 a_23699_8207# a_22917_8213# a_23615_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8958 io_out[1] a_4403_22869# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8960 a_2684_17231# _0873_.Y a_2381_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X8961 a_7258_5599# a_7090_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8962 a_14524_6549# _0901_.Q a_14744_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8964 a_8017_21263# _0935_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8967 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8969 a_24021_20181# a_23855_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8970 vssd1 _0797_.A1 a_8377_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X8971 a_14775_18589# a_14483_18543# a_14689_18589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X8972 vssd1 a_10073_26133# a_10007_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X8973 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8974 temp1.capload\[14\].cap.Y temp1.capload\[14\].cap_44.LO a_11797_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8975 vssd1 a_23415_19061# a_23373_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8976 a_2780_15285# a_2593_15325# a_2693_15543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X8979 vccd1 _0504_.A a_18059_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8980 vssd1 _0496_.X a_19439_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8981 vssd1 _0695_.A2 a_4524_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8982 a_25707_25321# _0854_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8983 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5796_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8984 vssd1 a_26099_15823# a_26267_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8985 a_20740_5487# a_20341_5487# a_20614_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8986 a_23469_9301# a_23303_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8987 a_4989_12879# _0758_.A1 a_4771_12791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X8988 a_9485_9301# a_9319_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8989 vssd1 _0685_.B a_6416_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8990 a_27590_12127# a_27422_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8993 a_7037_29177# _0825_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8994 _0579_.C a_13257_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X8995 _0444_.A a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8996 a_8228_21641# a_7829_21269# a_8102_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8997 vssd1 _0972_.CLK a_19531_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8998 a_15097_27797# a_14931_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8999 vssd1 a_27847_12381# a_28015_12283# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9000 a_27387_13469# a_26689_13103# a_27130_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9001 vssd1 a_28015_17723# a_27973_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9002 a_20893_27247# a_20727_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9003 a_25589_14735# _0966_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9004 _0873_.A a_2623_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9005 a_6833_13353# _0745_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X9008 vccd1 a_12743_8181# a_12659_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9014 vccd1 _0975_.CLK a_22659_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9015 _1053_.Q a_15963_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9016 vssd1 _0836_.A a_10147_15529# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X9017 a_23331_14557# a_22549_14191# a_23247_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9018 a_15945_21263# _0863_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9019 vccd1 a_18723_11445# a_18639_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9020 vccd1 _1053_.Q a_16258_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X9021 vssd1 _0722_.C a_5704_17461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
X9022 _0524_.X a_11582_13077# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9026 a_1766_29423# temp1.inv1_1.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9027 vssd1 a_8914_7093# a_8872_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9028 _0894_.Q a_26175_12283# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9030 vccd1 a_15595_23413# a_15511_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9031 a_26413_18543# a_26247_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9033 a_12889_4765# a_12355_4399# a_12794_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9035 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_6736_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9036 temp1.capload\[3\].cap.Y temp1.capload\[3\].cap.A a_15661_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9037 a_2686_27791# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9038 vccd1 _0508_.Y a_13735_12925# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9040 a_1941_4399# a_1775_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9041 _0708_.A3 a_4451_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X9042 a_22825_11177# _0926_.D a_22741_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9043 a_2773_25615# _1078_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9044 _0553_.X a_18243_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X9045 a_11041_17705# _0472_.X a_10791_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9046 a_20372_15113# a_19973_14741# a_20246_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9048 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X9049 a_5455_15279# _0778_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9050 vccd1 _0835_.A1 a_12342_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9051 a_6151_21781# _0764_.A1 a_6582_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X9052 vssd1 a_27038_4511# a_26996_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9053 _0845_.C1 a_4811_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9054 vssd1 _0812_.A2 a_10769_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9055 vccd1 a_25842_1247# a_25769_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9057 vccd1 a_9742_1247# a_9669_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9058 _0497_.B2 a_23047_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9059 a_21625_6575# _1006_.D a_21279_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9060 a_27517_10205# a_26983_9839# a_27422_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9061 a_23174_7093# a_23006_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9062 vccd1 a_21851_9019# a_21767_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9063 vccd1 _0888_.CLK a_6467_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9065 a_11888_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9066 a_24025_11471# _1014_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9067 _0963_.Q a_23507_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9070 a_20985_19631# a_20819_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9072 a_20556_20553# a_20157_20181# a_20430_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9073 vccd1 a_28015_15547# a_27931_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9075 vccd1 _0491_.X a_12245_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9076 fanout23.X a_27202_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9077 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_12999_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X9078 vssd1 _0460_.C a_2205_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9079 a_18590_4943# a_18151_4949# a_18505_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9081 a_21039_5853# a_20341_5487# a_20782_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9082 a_20027_6031# a_19329_6037# a_19770_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9083 vssd1 _1033_.CLK a_22567_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9084 vssd1 a_26099_1501# a_26267_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9085 vssd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_2686_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9086 a_10567_19061# _0771_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X9087 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9088 a_27149_3311# a_26983_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9089 _0626_.B1 a_17971_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X9090 vccd1 _0908_.CLK a_4351_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9091 _0787_.X a_6600_27907# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X9092 a_27548_2223# a_27149_2223# a_27422_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9093 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9094 a_1775_31375# _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9095 io_out[2] _0444_.A a_1591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9096 a_21909_21807# _1021_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9097 a_18616_18543# _0584_.A2 a_18125_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X9098 vssd1 a_1591_16367# _0722_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9099 vssd1 a_10167_1403# a_10125_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9100 a_25405_7663# _0621_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9101 a_5141_30199# _0809_.B2 a_5443_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X9103 a_17213_17455# a_17047_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9105 _0580_.C1 a_16127_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9106 a_17397_3855# a_16863_3861# a_17302_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9107 a_14011_7235# _0544_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9111 a_12355_22901# _0847_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X9112 _0816_.S _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9113 vccd1 _0847_.A2 a_1975_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X9114 vssd1 _0994_.CLK a_21555_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9116 vccd1 _0931_.CLK a_19439_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9117 _0543_.B2 a_17895_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9118 a_10643_4943# a_9945_4949# a_10386_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9120 a_8392_31599# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9121 a_4548_28335# a_4149_28335# a_4422_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9122 a_15078_17973# a_14910_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9123 _0630_.A1 a_17895_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9124 a_13360_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9125 a_17397_22895# a_17231_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9126 a_9669_21269# a_9503_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9128 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9129 a_26502_21085# a_26063_20719# a_26417_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9130 a_25309_9295# _0665_.B2 a_25225_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9131 vssd1 a_12467_10107# a_12425_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9133 vccd1 _0994_.CLK a_25879_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9134 _0999_.CLK a_22659_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X9137 _0584_.C1 a_22015_18112# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
R23 vssd1 temp1.capload\[7\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9140 a_2051_14848# _0456_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9142 _0937_.Q a_14767_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9143 a_6704_13077# _0745_.A1 a_6927_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9144 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13544_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9145 a_19517_6031# _0941_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9147 a_27149_23983# a_26983_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9148 a_10667_18543# _1078_.Q a_10576_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X9149 a_20267_6825# _0630_.A2 a_20349_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9150 a_10225_2223# _0637_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9151 a_26042_26525# a_25769_26159# a_25957_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9152 a_15370_1679# a_15097_1685# a_15285_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9153 a_17691_15279# _0523_.B1 a_17869_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9154 a_6733_12925# _0768_.A2 a_6651_12672# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9156 a_7005_5487# _0545_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9157 vccd1 _0829_.A1 a_9497_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X9158 vssd1 _0483_.X a_20145_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9160 vccd1 temp1.capload\[7\].cap.A temp1.capload\[7\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9161 vssd1 _1075_.Q a_15005_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X9162 a_23742_9295# a_23303_9301# a_23657_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9163 temp1.capload\[15\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9164 vccd1 a_15887_16733# a_16055_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9165 a_6319_3677# a_5455_3311# a_6062_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9166 vssd1 _0502_.X a_18673_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9167 a_9758_9295# a_9319_9301# a_9673_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9168 vssd1 fanout27.A a_18795_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9169 vccd1 _0445_.B a_14651_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X9170 vssd1 _0647_.X a_22199_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9171 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9172 vssd1 _0652_.A _0684_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9173 a_10147_15823# _0471_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9174 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15088_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9175 vssd1 a_2991_3579# a_2949_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9176 vccd1 _0513_.X a_13309_5515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X9178 vssd1 _0558_.X a_20819_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9179 _0630_.A2 _0842_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9180 vccd1 a_2566_3423# a_2493_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9181 a_26410_11293# a_25971_10927# a_26325_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9184 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_13544_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9185 a_11251_24233# _0444_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9186 vccd1 _0825_.S temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9187 _0761_.B a_5642_19637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9188 vccd1 a_17803_19899# a_17719_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9189 vccd1 _0845_.A1 a_7260_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9190 a_26225_19465# a_25235_19093# a_26099_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9191 vccd1 _0460_.C a_2051_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9192 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9193 a_4934_5737# _0694_.A2 a_4852_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9194 a_2405_25071# _0839_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9195 a_25769_21263# a_25235_21269# a_25674_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9196 a_6749_8207# _0681_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9197 vssd1 a_4802_27247# clkbuf_1_1__f__0390_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9198 a_8546_4917# a_8378_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9199 a_16853_8751# _0985_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X9200 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9201 vccd1 a_13422_9269# a_13349_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9202 a_15285_13103# _0511_.D a_15197_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X9203 vccd1 _1019_.CLK a_20727_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9204 _1079_.Q a_5015_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9205 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9206 vccd1 _0515_.B1 a_12069_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X9207 a_19770_6005# a_19602_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9208 vssd1 a_15793_6603# _0645_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X9209 vccd1 _0972_.CLK a_14931_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9210 vssd1 fanout37.A a_16495_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9211 vssd1 a_22879_16911# a_23047_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9212 a_2217_28335# a_2051_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9213 vssd1 a_19045_15797# _0658_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X9214 vssd1 _0850_.Y a_12428_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X9215 vccd1 _1019_.CLK a_19163_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9216 a_25842_14709# a_25674_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9217 a_7244_22057# _0866_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9218 a_21173_19631# _1023_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9219 a_13073_10389# a_12907_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9221 a_22465_9295# _0623_.D _0624_.D_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X9223 vccd1 _0471_.X _0840_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9224 a_25037_13103# _1011_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9226 a_9853_22357# a_9687_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9227 vssd1 a_10551_22351# a_10719_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9228 _0713_.A1 _0745_.A1 a_5731_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9229 a_18716_5321# a_18317_4949# a_18590_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9231 vccd1 _0893_.CLK a_25143_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9232 a_2842_2741# a_2683_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X9234 _0985_.D a_13939_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9235 vssd1 _0527_.X a_16061_10721# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9237 vccd1 a_10386_2741# a_10313_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9239 vccd1 _0821_.B a_11067_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9240 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9243 vccd1 _0922_.CLK a_9595_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9245 _0874_.X a_4300_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X9246 a_22270_26525# a_21831_26159# a_22185_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9248 vssd1 a_27590_2335# a_27548_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9249 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9251 a_21633_2223# _0575_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9253 a_23303_10383# _0558_.A2 a_23385_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X9254 vssd1 _0686_.X a_5812_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9255 _0925_.D a_15779_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9256 vssd1 _0795_.A1_N a_5904_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9257 vssd1 _0515_.X a_21647_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9258 vccd1 a_25455_16733# a_25623_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9259 vccd1 a_19183_4917# a_19099_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9260 vssd1 _1015_.CLK a_26983_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9261 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13735_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9262 a_21127_17249# _0504_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9263 vccd1 a_2823_2589# a_2991_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9264 vccd1 a_23431_7119# a_23599_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9265 vssd1 _0702_.B1_N a_5128_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9266 vccd1 a_25547_13469# a_25715_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9267 a_3983_18543# _0722_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9270 _0868_.A2 a_7244_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9272 vssd1 _0999_.CLK a_25235_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9273 a_14644_17455# _0662_.A1 a_14341_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X9275 a_10041_6031# _0901_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9276 vssd1 _0847_.A2 a_6876_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9278 a_10493_11849# a_9503_11477# a_10367_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9280 a_11793_15823# _0833_.A _0508_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9281 a_23579_14735# _0648_.A2 a_23757_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9282 a_27422_24349# a_26983_23983# a_27337_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9283 vccd1 a_23247_1501# a_23415_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9284 _0619_.B1 a_22325_6603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X9285 vccd1 _0809_.A1 a_5639_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9286 _0929_.Q a_24887_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9288 _1012_.Q a_28015_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9289 a_25033_6575# a_24867_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9292 vccd1 _0994_.CLK a_21555_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9294 a_22822_1501# a_22549_1135# a_22737_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9295 a_14651_24527# _0850_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9296 _0632_.B a_24887_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9298 a_25217_17455# a_25051_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9299 a_26091_3677# a_25309_3311# a_26007_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9300 vssd1 a_17895_2741# a_17853_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9301 a_6858_12015# _0745_.A3 a_6563_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X9302 _0847_.A2 a_11435_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9303 _0929_.Q a_24887_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9305 a_5601_18517# _0782_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X9306 vssd1 a_22015_8215# _1033_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9307 vssd1 _0558_.A2 a_25213_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X9308 a_16105_1135# _0946_.Q a_15759_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9309 a_11704_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9310 vccd1 a_2122_12015# a_2228_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X9311 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9312 a_9687_19881# _0751_.B1 a_9769_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X9314 _0854_.X a_25707_25321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X9315 a_24945_21807# _0929_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9316 vccd1 _0931_.CLK a_17047_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9317 a_2493_3677# a_1959_3311# a_2398_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9318 a_14829_6031# _0916_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X9320 vccd1 _0994_.CLK a_25235_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9321 vssd1 a_19439_13103# _0512_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X9323 a_12610_21807# a_12433_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9324 a_14441_13103# _1056_.Q a_14369_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
R24 vssd1 temp1.capload\[4\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9325 vccd1 _0722_.C a_3983_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9327 a_13912_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9328 _0715_.X a_2693_15543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9329 vccd1 _0523_.B1 a_22457_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9330 a_23637_12533# _0576_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9332 a_10551_22351# a_9687_22357# a_10294_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9333 vccd1 a_5047_21781# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9334 a_14405_20747# _0829_.A1 a_14319_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9335 _0807_.C a_5639_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9336 a_27847_15645# a_27149_15279# a_27590_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9337 a_24485_13647# _1046_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9338 vssd1 _0812_.A2 a_7663_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9339 vccd1 _0558_.A2 a_23745_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9340 a_12334_3855# a_12061_3861# a_12249_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9341 a_23868_9673# a_23469_9301# a_23742_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9342 a_15741_4399# a_15575_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9343 vssd1 a_17819_1679# a_17987_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9344 a_9884_9673# a_9485_9301# a_9758_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9346 a_22580_20553# a_22181_20181# a_22454_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9347 vssd1 _0563_.B1 a_27513_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X9349 a_5600_14165# _0734_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X9350 vssd1 _1030_.CLK a_19807_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9351 a_19605_10089# _0983_.D a_19521_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9352 vccd1 _0545_.A1 a_10356_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9353 a_24205_11471# a_23671_11477# a_24110_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9355 _0847_.A3 a_10055_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9356 vccd1 _0505_.A2 a_25777_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X9357 a_8116_10383# _0679_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9358 a_5639_12879# _0756_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9359 _0629_.X a_18059_17024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9360 a_7515_5853# a_6651_5487# a_7258_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9362 vssd1 a_20563_2741# a_20521_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9363 a_7902_6005# a_7734_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9364 a_5171_14851# _0722_.C a_5089_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9365 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9366 a_21993_13103# a_21003_13103# a_21867_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9367 vssd1 a_4985_12061# a_5091_12021# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9368 vccd1 clkbuf_1_1__f__0390_.A a_2686_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9369 a_26007_6031# a_25143_6037# a_25750_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9370 vssd1 a_3891_21263# _0814_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X9372 vccd1 a_27095_20987# a_27011_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9373 a_6081_2223# a_5915_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9375 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9376 a_3041_25071# a_2051_25071# a_2915_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9378 a_15795_27791# a_15097_27797# a_15538_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9379 a_2313_27247# _0837_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9380 a_10140_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9381 a_9811_22923# _0850_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9385 _0935_.CLK a_10791_16919# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9386 a_5905_15823# _0807_.C _0880_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9387 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9389 vccd1 _1076_.Q a_8031_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X9390 vssd1 a_26007_3677# a_26175_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9391 a_7653_9001# _0778_.A2 _0686_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9392 vssd1 fanout13.A a_15667_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9393 a_14729_14191# _1075_.Q a_14629_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X9394 a_25582_6031# a_25143_6037# a_25497_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9395 a_7745_8207# _0677_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9396 a_20947_21263# a_20083_21269# a_20690_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9397 vssd1 _0994_.D a_23308_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X9399 a_10229_15529# _0833_.A a_10147_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9400 a_10313_2767# a_9779_2773# a_10218_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9401 vccd1 _0959_.CLK a_11895_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9402 a_8661_7119# _0653_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9403 vccd1 a_11929_9633# _0491_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X9404 vssd1 a_3983_31849# io_out[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9405 vssd1 a_21334_27359# a_21292_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9406 clkbuf_1_0__f_net57.X a_1674_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9408 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9410 a_3333_19407# a_3141_19148# _0872_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X9411 vccd1 _0722_.A a_3983_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9412 a_11747_3677# a_11049_3311# a_11490_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9414 a_12069_4943# _0673_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X9415 _0684_.A1 _0651_.X a_15563_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9416 vssd1 _0917_.CLK a_9503_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9417 a_12694_23983# _0860_.A a_12316_24135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X9418 vccd1 a_28015_2491# a_27931_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9419 a_20529_5487# _0669_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9420 _0516_.B1 a_18645_7457# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X9422 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9424 a_2401_2773# a_2235_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9425 a_27337_5487# _0650_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9426 _0873_.A a_2623_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9427 vssd1 a_2623_6843# a_2581_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9428 vssd1 a_9919_6740# _1084_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9429 vssd1 _0664_.A2 a_23189_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9430 a_8205_13647# _0626_.B2 a_8123_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9432 vccd1 _0908_.CLK a_8583_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9433 a_22622_1653# a_22454_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9434 vccd1 fanout10.A a_12355_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X9437 _0908_.CLK a_1959_4951# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9438 a_22879_22351# a_22015_22357# a_22622_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9439 _0966_.Q a_27095_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9440 vssd1 a_3799_11471# _0861_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X9443 a_6319_3677# a_5621_3311# a_6062_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9444 vccd1 a_27003_11195# a_26919_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9445 _0662_.B1 a_21127_17249# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9447 a_25842_25589# a_25674_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9448 vssd1 _0726_.X a_5047_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X9449 a_25455_2589# a_24591_2223# a_25198_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9450 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_7387_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9451 vssd1 a_12575_6031# a_12743_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9452 _0489_.X a_19531_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X9453 a_23745_14735# _0999_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9454 vccd1 a_10073_26133# a_10103_26486# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9456 vssd1 a_21242_20831# a_21200_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9457 _0619_.B2 a_27923_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9459 vccd1 a_27555_13371# a_27471_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9460 vssd1 _0825_.S temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X9461 vssd1 _0619_.X _0624_.D_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9462 vccd1 a_22990_19061# a_22917_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9464 a_22549_22351# a_22015_22357# a_22454_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9465 a_9003_15797# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X9467 a_25401_19093# a_25235_19093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9468 vssd1 a_15151_10205# a_15319_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9469 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9470 vccd1 a_19439_13103# _0512_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X9471 _0641_.D1 a_11711_1792# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9472 a_19521_10749# _0521_.A a_19439_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9474 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9476 a_22963_16911# a_22181_16917# a_22879_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9477 _0735_.Y _0717_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X9478 _0680_.Y _0655_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X9480 vccd1 a_12355_8751# _0535_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X9482 a_20303_17821# a_19605_17455# a_20046_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9483 vccd1 a_13479_2741# a_13395_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9484 a_25842_7093# a_25674_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9485 a_19015_4943# a_18317_4949# a_18758_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9486 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9487 vssd1 _1019_.CLK a_18335_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9490 a_27755_9117# a_27057_8751# a_27498_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9492 vssd1 _0835_.A1 a_11344_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X9493 vssd1 fanout23.X a_26431_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9494 a_13432_26409# a_13183_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9495 _0594_.C a_15759_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9496 a_22879_1679# a_22181_1685# a_22622_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9497 a_22622_15797# a_22454_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9498 a_19041_17277# _1020_.Q a_18969_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9499 _0590_.B2 a_20839_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9500 a_20522_21263# a_20249_21269# a_20437_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9501 a_9865_28335# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9502 a_4439_24233# _0814_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9503 a_12659_6031# a_11877_6037# a_12575_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9504 a_2852_15285# _0722_.A a_2780_15285# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X9505 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9507 _0574_.X a_22751_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9510 a_6336_15253# _0758_.A1 a_6556_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9511 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9513 a_1639_7338# io_in[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9514 vssd1 a_24887_1653# a_24845_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9515 vssd1 _0664_.X a_25143_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9516 a_21591_27613# a_20727_27247# a_21334_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9517 a_27111_18909# a_26413_18543# a_26854_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9518 vssd1 _0533_.X a_13989_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9519 a_13069_3311# _0910_.Q a_12723_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9520 vssd1 _1015_.CLK a_23303_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9521 vccd1 a_24278_11445# a_24205_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9522 a_7285_9661# _0655_.X a_7203_9408# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9523 vssd1 _0917_.CLK a_9319_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9524 vssd1 a_23763_10927# _1015_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9525 a_4149_28335# a_3983_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9526 vccd1 a_15319_10107# a_15235_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9527 vssd1 _0931_.CLK a_20083_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9528 vccd1 _0836_.A a_12995_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X9529 a_27337_9839# _0572_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9530 a_27379_4765# a_26597_4399# a_27295_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9532 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9533 vccd1 a_6487_3579# a_6403_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9535 vccd1 a_9999_1501# a_10167_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9537 a_25639_12559# a_24775_12565# a_25382_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9538 a_2686_28879# clkbuf_1_1__f__0390_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9539 a_21261_27613# a_20727_27247# a_21166_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9540 a_15922_21085# a_15649_20719# a_15837_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9541 a_25030_22173# a_24757_21807# a_24945_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9542 a_22822_14557# a_22383_14191# a_22737_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9543 a_22659_11471# _0662_.B1 a_22741_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9544 _0847_.X a_1735_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9546 a_27847_14557# a_27149_14191# a_27590_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9547 vssd1 a_5142_4511# a_5100_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9548 a_4981_4943# _0677_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9549 a_4262_25393# a_4213_25223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X9550 vssd1 _0645_.B2 a_17236_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X9551 vssd1 _0888_.CLK a_6467_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9552 a_23431_7119# a_22567_7125# a_23174_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9553 a_6062_3423# a_5894_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9556 a_4040_10901# a_4251_11249# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X9557 vssd1 _0994_.CLK a_22015_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9558 a_23247_3677# a_22549_3311# a_22990_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9559 a_10589_10927# a_10423_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9561 a_25030_15645# a_24591_15279# a_24945_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9562 a_19557_6603# _0512_.A a_19471_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9563 a_6831_22351# _0868_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9564 a_16013_16367# a_15023_16367# a_15887_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9565 a_13529_2057# a_12539_1685# a_13403_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9566 a_14913_3311# a_14747_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9569 a_19991_5056# _0632_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9570 a_25708_6409# a_25309_6037# a_25582_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9571 _0614_.X a_15483_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X9573 vccd1 a_3028_14165# _0758_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X9574 a_21069_16617# _0559_.X a_20997_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9575 _0576_.D1 a_22015_6144# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9576 a_6000_25077# a_5813_25117# a_5913_25335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X9577 vssd1 a_14894_12127# a_14852_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9578 _0920_.D a_15135_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9579 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9580 a_15002_23439# a_14729_23445# a_14917_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9581 a_15576_21379# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9582 a_4864_15797# _0456_.A a_5256_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X9583 vssd1 _0959_.CLK a_12447_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9584 _0986_.D a_10535_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9586 _0602_.X a_18887_17024# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9587 vccd1 a_24243_21237# a_24159_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9589 a_13081_27791# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE _0824_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9590 vssd1 a_10811_1653# a_10769_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9591 vccd1 a_8159_6031# a_8327_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9592 vccd1 io_in[4] a_1591_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X9593 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9594 vssd1 _0931_.CLK a_19439_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9595 vssd1 _0803_.X a_4929_19659# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9596 _0620_.X a_25143_14441# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9597 a_4847_1501# a_4149_1135# a_4590_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9598 vssd1 _0922_.CLK a_2787_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9600 vccd1 a_24887_20149# a_24803_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9601 a_25214_12559# a_24941_12565# a_25129_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9602 vssd1 _0858_.A2 a_12068_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9603 vccd1 a_21775_18909# a_21943_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9604 a_4729_26703# _0833_.Y a_4984_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9606 a_9573_14191# _0835_.A1 _0717_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X9607 a_27973_9839# a_26983_9839# a_27847_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9609 _0564_.C a_19531_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X9610 a_9588_16617# _0880_.A2 _0880_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X9611 vccd1 _0584_.A2 a_17857_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9612 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X9613 a_21265_18543# _0991_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9614 _0711_.B _0710_.B1 a_5445_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9615 clkbuf_1_0__f_io_in[0].X a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9616 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13432_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9617 a_22162_21919# a_21994_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9619 vssd1 a_26267_19061# a_26225_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9620 vssd1 _0932_.Q a_18616_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X9623 a_20310_17231# _1022_.Q a_20220_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X9624 vssd1 a_15667_21807# _1019_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9625 a_27337_2223# _0665_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9626 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9627 _0994_.CLK a_21279_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X9628 a_10125_5487# a_9135_5487# a_9999_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9629 vccd1 a_4403_22869# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9630 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9631 vccd1 a_22990_1247# a_22917_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9632 _0670_.A2 a_16895_5281# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X9634 vccd1 _0847_.A2 a_5445_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9635 a_7477_17999# _0813_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9636 a_26318_23261# a_25879_22895# a_26233_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9637 vccd1 _0666_.X a_16209_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9639 vccd1 a_5141_30199# io_out[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X9640 a_11797_29199# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9641 a_25589_16911# _0999_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9642 vssd1 a_11458_17429# _0574_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9643 a_22181_15829# a_22015_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9644 a_17117_8751# _0615_.A1 a_16771_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9645 vccd1 _0850_.A a_8338_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9646 a_27422_3677# a_27149_3311# a_27337_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9647 a_15575_19200# _0860_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9648 _0840_.A0 _0471_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X9649 vssd1 _0722_.A a_4324_14197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X9652 vccd1 a_21334_27359# a_21261_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9653 _0877_.A2 _0439_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X9654 vccd1 clkbuf_1_0__f_io_in[0].X a_1591_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9655 a_25999_9117# a_25217_8751# a_25915_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9656 a_26225_10761# a_25235_10389# a_26099_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9657 a_20046_17567# a_19878_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9658 vccd1 a_16745_6549# _0646_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X9659 a_8175_11989# _0654_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X9660 vccd1 a_6467_16367# _0717_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X9661 vssd1 _0824_.Y a_13183_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9662 vccd1 a_25658_7775# a_25585_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9663 vssd1 a_16829_12161# _0565_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X9664 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9665 vccd1 a_12502_3829# a_12429_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9666 _0607_.B a_21575_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9667 a_10451_11471# a_9669_11477# a_10367_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9668 _0854_.B a_11895_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9669 _0669_.B2 a_23691_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9670 a_2382_4511# a_2214_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9671 a_8803_4943# a_7939_4949# a_8546_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9672 vssd1 _1019_.CLK a_20727_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9674 vssd1 a_12743_13621# a_12701_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9675 fanout24.A a_16495_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X9677 vssd1 _0609_.X a_15483_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X9678 a_27548_17455# a_27149_17455# a_27422_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9679 vccd1 a_7683_5755# a_7599_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9680 vssd1 a_14341_15797# _0763_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9681 a_24167_9295# a_23303_9301# a_23910_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9683 a_23247_14557# a_22383_14191# a_22990_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9684 a_27590_7775# a_27422_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9685 a_2686_27791# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9687 a_24941_8213# a_24775_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9688 vccd1 _0722_.A a_3129_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X9690 a_12429_3855# a_11895_3861# a_12334_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9691 vccd1 _0840_.A0 a_13735_12925# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X9693 vccd1 a_9791_12015# a_9911_12061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X9694 vssd1 a_14433_24501# _0852_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9695 vccd1 _0908_.CLK a_7939_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9696 vssd1 _0643_.B1 a_23833_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X9697 _0590_.B2 a_20839_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9698 vssd1 _0893_.CLK a_25143_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9699 a_9016_31055# a_8767_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9700 vccd1 _1062_.CLK a_26247_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9701 a_9574_5853# a_9301_5487# a_9489_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9702 a_10589_10927# a_10423_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9703 vccd1 a_17635_19997# a_17803_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9707 a_1945_8751# _0875_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9708 vssd1 _0479_.Y a_13551_8215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9711 a_5992_14441# _0735_.A2 a_5737_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9712 a_9117_3855# a_8583_3861# a_9022_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9713 a_16829_12161# _0564_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9715 a_20671_8029# a_19973_7663# a_20414_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9716 a_6645_12265# _0745_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X9717 a_4984_26703# _0845_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9718 a_7565_22671# _0866_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9719 a_5809_3311# _0566_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9721 a_21134_11177# _0662_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9722 vccd1 a_23339_21085# a_23507_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9723 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X9724 vccd1 fanout23.X a_26983_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9725 temp1.capload\[11\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9726 vccd1 a_23599_7093# a_23515_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9727 a_1766_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9730 vssd1 _0861_.X a_3326_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9731 vccd1 a_17267_22173# a_17435_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9732 _1022_.Q a_22587_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9733 a_6808_29967# a_6559_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9734 vccd1 a_25623_2491# a_25539_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9736 vccd1 a_12777_24501# fanout13.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9740 a_26183_1501# a_25401_1135# a_26099_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9741 a_24945_5487# _1031_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9742 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X9743 a_6559_19631# _0807_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9745 _0893_.Q a_28015_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9746 vssd1 _1075_.Q a_14471_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9747 a_9949_13647# _0921_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9748 a_25198_2335# a_25030_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9749 a_25033_6575# a_24867_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9750 vccd1 _0798_.A1 a_4342_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9751 vssd1 a_2655_24501# _0839_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X9752 a_12525_21263# _0934_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9753 a_25731_6941# a_24867_6575# a_25474_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9754 a_25217_17455# a_25051_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9755 a_4847_2589# a_3983_2223# a_4590_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9757 a_19770_6005# a_19602_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9758 a_1775_28879# _0836_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9759 a_24591_11177# _0664_.A2 a_24673_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9761 _0491_.X a_11929_9633# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X9762 _0722_.A a_1591_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9763 vssd1 _0444_.B a_1775_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9764 vccd1 a_12207_15645# a_12375_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9765 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8392_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9766 vssd1 _0931_.CLK a_17047_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9768 a_23592_18377# a_23193_18005# a_23466_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9769 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13360_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9770 vssd1 a_23855_15831# _0964_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9771 a_4337_31599# _0814_.A1 a_3983_31849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9772 a_22714_2741# a_22546_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9773 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9776 a_25585_8029# a_25051_7663# a_25490_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9777 vccd1 _0836_.A a_11793_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9778 vccd1 temp1.capload\[5\].cap_50.LO temp1.capload\[5\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9779 vccd1 a_1757_26703# _0832_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X9781 a_20111_26703# a_19329_26709# a_20027_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9782 a_4342_30761# _0798_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X9783 a_26686_18909# a_26247_18543# a_26601_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9784 vssd1 a_6423_8903# _0698_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X9785 vccd1 a_21023_22325# a_20939_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9786 _0576_.B1 a_24315_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9788 _0959_.D a_10811_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9789 a_23569_6825# _0552_.B2 a_23487_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9790 a_24209_22351# _0928_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9791 vssd1 a_7896_11703# _0734_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X9793 a_27590_9951# a_27422_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9794 a_11697_20719# _0987_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9795 a_12532_28335# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9796 a_18317_4949# a_18151_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9797 _0504_.A a_18703_12567# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X9798 vssd1 a_1585_24135# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.209625 pd=1.295 as=0.08775 ps=0.92 w=0.65 l=0.15
X9799 _0685_.X a_6651_12672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9800 _0619_.B2 a_27923_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9801 a_4356_23983# _0774_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9802 a_14833_17277# a_14563_16911# a_14729_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9803 a_19234_1679# a_18961_1685# a_19149_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9804 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_10699_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9807 _0591_.X a_14655_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X9808 a_22990_14303# a_22822_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9809 vssd1 a_6522_2335# a_6480_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9811 vccd1 _1078_.Q a_14637_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X9812 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9814 _1041_.Q a_21575_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9815 vssd1 _0788_.C a_6072_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X9817 a_26225_4233# a_25235_3861# a_26099_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9818 a_20430_22351# a_19991_22357# a_20345_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9819 vssd1 clkbuf_0__0390_.A a_4802_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9820 a_11152_30511# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9821 a_7203_9408# _0685_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9822 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].vref.TE a_18059_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9824 vccd1 _0471_.X a_10147_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9825 a_11238_19631# _0441_.B a_11149_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X9826 vssd1 a_2686_27791# _0798_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9827 a_5243_14851# _0722_.B a_5171_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9828 vssd1 a_18611_14191# _0931_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9829 vssd1 a_6608_29111# _0825_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X9830 vccd1 a_7900_14165# _0770_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X9831 vssd1 _0735_.A2 a_11505_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9832 a_5273_29687# _0445_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9833 _0444_.A a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9834 vssd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_1766_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9835 vssd1 _0565_.B1 a_14524_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X9836 vccd1 _0832_.A a_4075_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9837 _0778_.Y _0778_.A2 a_5537_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X9839 a_10110_21237# a_9942_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9840 vssd1 a_4958_2741# a_4916_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9841 a_10218_4943# a_9779_4949# a_10133_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9842 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9843 vccd1 _0807_.A a_5905_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9844 a_2581_6409# a_1591_6037# a_2455_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9846 vccd1 _0972_.CLK a_18795_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9848 a_15335_17999# a_14637_18005# a_15078_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9849 vccd1 _0471_.X _0840_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9850 vccd1 a_2823_27613# a_2991_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9851 vccd1 _0935_.CLK a_11343_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9853 a_23005_16201# a_22015_15829# a_22879_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9854 a_23385_10383# _0621_.B2 a_23303_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9859 a_15093_20553# a_14103_20181# a_14967_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9860 vssd1 _1076_.Q a_13091_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9861 vssd1 a_25623_4667# a_25581_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9862 vssd1 a_20671_14735# a_20839_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9863 _0533_.X a_16897_12897# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X9864 _0669_.B2 a_23691_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9866 a_25769_15823# a_25235_15829# a_25674_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9867 vccd1 _0502_.X a_22015_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9868 a_4167_17999# _0722_.B a_4589_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9869 a_17470_2741# a_17302_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9870 a_26502_21085# a_26229_20719# a_26417_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9871 a_6336_15253# _0735_.A2 a_6728_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X9872 _0513_.X a_9911_12061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X9874 vccd1 fanout24.A a_22015_8215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X9875 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9876 a_9815_16911# a_8951_16917# a_9558_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9877 a_5817_6351# _0681_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9878 a_5721_12559# _0791_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9879 a_5731_10703# _0745_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9880 vccd1 _1053_.CLK a_9687_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9881 vccd1 a_20855_20175# a_21023_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9882 a_11609_6825# _0674_.C1 a_11527_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9883 vccd1 a_11685_25045# fanout11.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X9884 a_14729_23445# a_14563_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9885 a_11711_1792# _0905_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9886 vssd1 _0605_.C1 a_17289_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X9887 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_4811_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9888 _0925_.D a_15779_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9889 a_5031_1679# a_4333_1685# a_4774_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9890 a_2949_1135# a_1959_1135# a_2823_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9891 vccd1 _0523_.B1 a_22365_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9893 vssd1 _1028_.CLK a_13275_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9894 vccd1 a_13771_10383# a_13939_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9895 vssd1 a_11030_11039# a_10988_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9896 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_5547_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9897 _0809_.B2 a_3155_21271# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X9898 vssd1 a_20855_20175# a_21023_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9899 vccd1 _0835_.A1 _0749_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9901 vssd1 a_4772_13621# _0794_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X9902 a_12042_9951# a_11874_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9903 vssd1 _0888_.CLK a_4535_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9904 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9905 vssd1 a_6613_22325# _0868_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9906 a_25589_7119# _0573_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9907 a_9485_16911# a_8951_16917# a_9390_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9908 a_6287_21807# _0797_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X9909 vssd1 a_3270_2741# a_3228_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9910 vccd1 _0460_.C a_1945_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X9911 a_13432_26703# a_13183_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9914 _1013_.Q a_28015_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9916 a_6835_15055# _0794_.A2 a_6741_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X9917 vssd1 _0614_.X a_17971_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9918 a_18716_20553# a_18317_20181# a_18590_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9919 vssd1 a_18371_11293# a_18539_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9920 a_17811_15073# _0521_.A a_17725_15073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9921 a_25455_16733# a_24757_16367# a_25198_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9922 a_20138_2741# a_19970_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9923 vccd1 a_1591_9839# _0466_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X9924 a_19593_10749# _0607_.B a_19521_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9925 vccd1 a_21150_4511# a_21077_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9927 _0946_.D a_15871_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9928 _0645_.B2 a_15963_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9929 a_4149_28335# a_3983_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9930 a_1775_27791# _0845_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9931 _0653_.A1 a_7499_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9934 a_4589_17999# _0722_.C _0798_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9935 a_26099_14735# a_25401_14741# a_25842_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9936 a_27590_16479# a_27422_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9937 _0847_.A2 a_11435_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X9938 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11704_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9940 vccd1 _0579_.C a_18059_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9941 a_16182_4511# a_16014_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9943 a_24945_2223# _1035_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9944 a_26962_13469# a_26689_13103# a_26877_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9945 _0988_.Q a_10535_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9946 a_24462_1653# a_24294_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9947 vssd1 _0710_.B1 a_4259_7669# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X9948 a_6556_8751# _0656_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X9951 vccd1 a_24719_22351# a_24887_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9954 vssd1 a_27847_16733# a_28015_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9955 vccd1 a_27590_3423# a_27517_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9956 a_16140_14191# a_15741_14191# a_16014_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9957 a_17470_2741# a_17302_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9958 a_15829_2223# a_14839_2223# a_15703_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9959 a_25589_19087# _1067_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9960 vssd1 a_19439_13103# _0512_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9961 a_7457_10089# _0778_.A2 _0680_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9962 a_27111_18909# a_26247_18543# a_26854_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9963 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9964 vssd1 a_24719_22351# a_24887_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9965 vccd1 _0931_.CLK a_20911_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9967 vssd1 _1028_.CLK a_14563_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9969 vccd1 _0861_.B1 a_4429_16672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X9970 a_27167_11471# _0619_.B1 a_27249_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9971 vccd1 _0513_.X a_13367_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9972 vccd1 a_25899_6843# a_25815_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9973 a_16127_13103# _0917_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9974 a_12849_12879# a_12447_12559# a_12763_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X9975 _0610_.X a_13551_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9976 vccd1 a_8971_4917# a_8887_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9980 a_21813_7913# _1003_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9982 _0565_.A1 a_15319_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9983 a_23040_20719# a_22641_20719# a_22914_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9984 vccd1 io_in[0] a_2962_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9985 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9986 vssd1 _1078_.Q a_14913_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X9987 a_3283_25615# a_2585_25621# a_3026_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9988 io_out[0] a_5047_21781# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9989 vccd1 a_14483_18543# a_14603_18589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X9991 vccd1 a_24335_9269# a_24251_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9993 vssd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_1674_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9994 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9995 vssd1 a_8235_4667# a_8193_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9996 a_13633_6031# _0538_.C1 a_13551_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9997 a_13422_9269# a_13254_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
R25 vccd1 temp1.capload\[11\].cap_41.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9998 a_9313_10703# _0466_.A a_9095_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X9999 a_9781_10927# a_9495_11249# a_9284_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10000 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10001 vccd1 a_18611_14735# _0662_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10002 _0570_.X a_23303_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10003 vssd1 _0848_.X a_12114_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10004 a_20138_2741# a_19970_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10005 a_1945_9295# _1084_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X10006 vssd1 a_1674_31599# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10007 vssd1 _0466_.A _0546_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10008 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10009 a_3026_25589# a_2858_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10010 vccd1 a_9742_5599# a_9669_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10011 a_27517_14557# a_26983_14191# a_27422_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10012 a_10551_22351# a_9853_22357# a_10294_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10013 a_25593_11791# _1013_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X10014 vssd1 a_6704_13077# _0747_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X10016 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8767_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10017 vssd1 _0812_.A2 a_5720_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10020 a_25129_8207# _0621_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10021 a_27149_17455# a_26983_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10022 a_10344_5321# a_9945_4949# a_10218_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10024 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10025 a_2687_2045# a_2114_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1197 ps=1.41 w=0.42 l=0.15
X10026 _0962_.D a_15319_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10027 a_18774_25615# a_18335_25621# a_18689_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10028 vccd1 a_2455_6941# a_2623_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10029 vccd1 a_4590_26271# a_4517_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10030 a_11068_16617# _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10031 a_14524_6549# _0531_.X a_14916_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X10032 _0609_.C1 a_19439_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10033 a_21813_7913# _0967_.Q a_21729_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10034 a_20548_17231# _0512_.X a_20057_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X10035 vssd1 a_2114_1653# _0860_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X10037 vccd1 a_15503_17973# a_15419_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10038 a_2639_4765# a_1775_4399# a_2382_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10039 a_15023_11471# _0667_.B1 a_15105_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X10041 io_out[7] a_3983_31849# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X10044 vssd1 a_2823_3677# a_2991_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10045 a_6559_10383# _0778_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10046 vccd1 a_26635_26427# a_26551_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10047 vssd1 a_6611_25589# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10048 vccd1 _0809_.B2 a_5245_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10050 vssd1 a_3799_11471# _0861_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10052 vccd1 _0752_.Y io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10053 _0836_.A a_8031_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10054 vssd1 _0609_.C1 a_17657_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X10055 a_27149_7663# a_26983_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10056 vccd1 a_26083_9019# a_25999_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10059 vccd1 a_11803_23439# _0444_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10060 vccd1 a_9558_16885# a_9485_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10061 a_17928_8181# _0587_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X10062 vccd1 _0827_.A a_13081_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X10063 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_13432_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10064 _1068_.Q a_27279_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10065 a_4789_4233# a_3799_3861# a_4663_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10066 _0831_.D a_9811_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X10067 a_23818_21237# a_23650_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10068 vssd1 a_10167_5755# a_10125_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10070 vccd1 _0975_.CLK a_24591_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10071 vccd1 _0931_.CLK a_16771_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10072 vccd1 _0513_.X a_13735_3968# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10073 a_9850_4765# a_9411_4399# a_9765_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10074 a_20257_7119# _0941_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X10075 a_25122_13469# a_24683_13103# a_25037_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10076 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X10077 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9016_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10078 a_23523_9117# a_22659_8751# a_23266_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10079 vccd1 a_19439_13103# _0512_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10080 vssd1 a_1766_29423# clkbuf_1_1__f_net57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10081 vssd1 _0735_.A2 a_8479_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X10082 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_4811_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10083 _0965_.D a_24059_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10084 a_4153_3855# _0908_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10085 a_2037_3855# _0882_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10087 a_15793_6603# _0504_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10088 vccd1 a_22035_13371# a_21951_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10089 a_23650_21263# a_23377_21269# a_23565_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10090 a_24945_15279# _0891_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10091 vccd1 _1062_.CLK a_25235_19093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10092 a_4590_2335# a_4422_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10093 a_22879_22351# a_22181_22357# a_22622_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10094 a_22879_16911# a_22015_16917# a_22622_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10097 a_26325_10927# _1063_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10098 vssd1 _0824_.Y a_13183_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10100 vssd1 a_4771_12791# _0734_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10101 vccd1 a_11760_26935# _0823_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X10102 a_22454_22351# a_22015_22357# a_22369_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10103 vccd1 _1076_.Q a_10055_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X10104 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10105 vssd1 a_10535_21237# a_10493_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10106 _0813_.A2 a_4132_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X10108 vssd1 a_21610_24095# a_21568_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10109 vssd1 a_18645_7457# _0516_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X10111 _0801_.X a_14319_20747# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X10112 a_20027_6031# a_19163_6037# a_19770_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10113 a_23119_10089# _0487_.X a_23201_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X10114 a_7602_23555# _0441_.B a_7520_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10115 vccd1 a_26267_14709# a_26183_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10116 vccd1 _0460_.C a_2879_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X10117 a_25674_4943# a_25401_4949# a_25589_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10118 a_15565_7235# _0642_.D_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10119 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A a_7932_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10120 vccd1 a_27847_22173# a_28015_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10121 a_25401_14741# a_25235_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10122 vssd1 _1015_.CLK a_25971_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10123 a_22549_16911# a_22015_16917# a_22454_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10124 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10125 a_11322_3677# a_10883_3311# a_11237_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10127 a_7256_17429# _0812_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X10128 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10129 vssd1 _0511_.D a_13533_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X10130 a_17906_13647# _0608_.X a_17657_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10131 vssd1 a_1867_15831# _0722_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X10132 a_27245_8751# _0647_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10133 a_19602_6031# a_19163_6037# a_19517_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10134 _0845_.A2 a_2686_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10136 a_25639_8207# a_24941_8213# a_25382_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10137 a_15023_11471# _0667_.B1 a_15105_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10138 vccd1 a_15779_3579# a_15695_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10139 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_14188_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10140 a_9687_19881# _0751_.B1 a_9769_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10142 a_20897_3311# _1040_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10143 a_17029_7119# _1029_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X10144 a_4252_20291# _0722_.C a_4170_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10145 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10146 vccd1 a_19402_1653# a_19329_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10148 vssd1 a_10107_10615# _0626_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10152 a_15354_3423# a_15186_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10153 vssd1 a_20025_10955# _0643_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X10155 a_5626_28879# _0825_.S a_5323_29111# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X10156 vccd1 a_20395_2767# a_20563_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10157 a_26597_4399# a_26431_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10158 _0721_.A a_2975_17461# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X10160 vccd1 a_8079_28500# _0821_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10161 vssd1 a_23818_21237# a_23776_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10162 a_21426_19743# a_21258_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10163 vssd1 a_3727_4917# a_3685_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10165 a_15277_5487# _0543_.A1 a_14839_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10166 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11960_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10167 vccd1 _0698_.A2_N a_4251_11249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X10168 vssd1 _0824_.Y a_12355_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10169 vssd1 _0959_.CLK a_9779_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10170 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10171 vccd1 a_4132_17429# _0813_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10172 _1033_.CLK a_22015_8215# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10173 vccd1 a_9963_17455# _0511_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10174 vccd1 _1033_.CLK a_24867_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10175 a_19793_17455# _0937_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10176 a_19329_1679# a_18795_1685# a_19234_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10177 _0653_.A1 a_7499_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10178 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10179 a_23266_8863# a_23098_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10180 vssd1 a_13422_9269# a_13380_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10181 a_26007_3677# a_25143_3311# a_25750_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10182 vssd1 _0506_.A2 a_23097_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X10183 vccd1 a_21242_20831# a_21169_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10184 a_5234_4917# a_5066_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10185 a_13360_28335# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10186 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10187 a_6269_2223# _0910_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10188 _0710_.A2 _0689_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10189 a_27330_9117# a_26891_8751# a_27245_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10190 _0583_.A a_20635_13655# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10191 vssd1 a_23487_15279# _0893_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10193 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10194 a_6582_21807# _0797_.B1 a_6287_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X10195 a_2686_23439# clkbuf_1_1__f__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10196 _0605_.D1 a_13367_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10198 vccd1 a_1639_7828# input3.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10199 _0805_.A a_4843_19659# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X10200 a_4065_18543# _0456_.A a_3983_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10201 a_25030_16733# a_24757_16367# a_24945_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10203 _0622_.A1 a_18539_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10204 a_7004_8207# _0685_.X a_6749_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X10205 vssd1 _1053_.CLK a_14931_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10207 _0840_.X a_4403_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10208 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X10209 a_25455_5853# a_24757_5487# a_25198_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10210 a_27973_12015# a_26983_12015# a_27847_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10211 a_27931_12381# a_27149_12015# a_27847_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10213 _0758_.A1 a_3028_14165# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X10214 vccd1 a_10367_11471# a_10535_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10215 a_26045_22895# a_25879_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10216 a_13714_4943# a_13441_4949# a_13629_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10218 temp1.capload\[8\].cap.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10219 vccd1 _0489_.X a_19689_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10220 a_2589_2767# _0852_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X10221 _0565_.A1 a_15319_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10223 vccd1 _0816_.S temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10224 a_4705_2767# _0586_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10225 a_11969_10205# a_11435_9839# a_11874_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10226 vssd1 a_10367_11471# a_10535_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10227 _0872_.A1 a_4386_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10228 a_9669_11477# a_9503_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10229 a_26099_19997# a_25401_19631# a_25842_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10230 vccd1 a_6336_15253# _0760_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X10232 vccd1 _0994_.CLK a_26983_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10233 a_9407_18793# _0812_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10234 vccd1 a_7625_14709# _0793_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X10235 a_25842_1247# a_25674_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10238 vssd1 _0994_.CLK a_26983_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10239 vssd1 a_7111_13655# _0735_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X10240 a_19697_3855# a_19163_3861# a_19602_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10241 a_9742_1247# a_9574_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10242 a_20027_26703# a_19329_26709# a_19770_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10245 a_26927_21085# a_26229_20719# a_26670_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10246 a_16208_25935# _0861_.A1 a_15905_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X10247 vssd1 _0908_.CLK a_5915_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10248 a_9976_4399# a_9577_4399# a_9850_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10249 _0839_.Y _0839_.B a_5547_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10250 _0522_.B1 a_16897_16395# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X10251 vssd1 _0656_.Y a_7032_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17875 ps=1.2 w=0.65 l=0.15
X10252 a_21468_10927# _0643_.B1 a_20977_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X10253 vccd1 _0856_.Y a_11983_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X10254 a_17727_2767# a_16863_2773# a_17470_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10255 vssd1 a_2686_31055# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10256 _0847_.B1 a_10515_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X10257 a_18095_23261# a_17231_22895# a_17838_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10258 a_17971_10089# a_17865_9845# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X10260 a_4929_19659# _0440_.A a_4843_19659# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10261 a_15193_2223# _0945_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10262 a_15641_8323# _0675_.B a_15569_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10263 _0840_.A1 a_2991_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10266 a_17625_16161# _0602_.A a_17539_16161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10267 a_18256_11849# a_17857_11477# a_18130_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10268 vccd1 _0849_.X a_12433_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X10269 a_18777_21263# a_18243_21269# a_18682_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10270 vccd1 _1015_.CLK a_25051_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10271 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10272 vccd1 a_5642_19637# _0761_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X10273 a_12065_11471# _0580_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10274 a_14655_2767# _0670_.A2 a_14737_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X10275 vssd1 a_2455_6941# a_2623_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10276 vssd1 _1033_.CLK a_25051_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10279 temp1.capload\[13\].cap.Y temp1.capload\[13\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10280 a_2861_4949# a_2695_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10281 a_12893_21807# a_12716_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X10282 a_2198_9269# a_2039_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X10284 a_9313_20495# _0813_.A2 a_9095_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X10285 vssd1 a_17470_2741# a_17428_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10286 _0549_.B2 a_8971_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10287 vssd1 _0643_.X a_15667_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10288 _0555_.C1 a_11987_2473# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X10289 a_7571_18319# _0739_.A2 a_7477_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X10290 vccd1 a_8175_9527# _0689_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X10291 vssd1 a_4036_30663# _0798_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X10292 a_10493_21641# a_9503_21269# a_10367_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10293 _0461_.A a_3983_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10294 a_14260_26703# a_14011_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10295 _0543_.A1 a_13571_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10296 a_11448_3311# a_11049_3311# a_11322_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10297 a_24673_10927# _1011_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X10298 a_10037_2223# a_9871_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10300 a_19728_6409# a_19329_6037# a_19602_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10301 _1056_.Q a_10719_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10303 vssd1 io_in[5] a_1626_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10304 _0574_.C a_11458_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10305 vssd1 _0964_.CLK a_22015_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10306 vccd1 _1015_.CLK a_25971_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10308 _0595_.D a_18427_2473# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X10309 _0768_.B1 a_4165_14455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10310 vccd1 _0840_.A1 a_15575_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10312 _0812_.A2 a_1775_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10313 _1041_.Q a_21575_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10314 a_1863_24233# _0765_.B1 a_1585_24135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10315 _1056_.Q a_10719_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10316 a_20598_22325# a_20430_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10317 vssd1 _1030_.CLK a_19163_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10318 vssd1 a_14524_6549# _0544_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X10319 vccd1 _0602_.A a_20635_13655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X10320 vccd1 _0831_.D a_1757_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
D4 vssd1 _0861_.X sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X10322 a_9095_10615# _0466_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X10323 _0619_.X a_27167_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X10324 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5888_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10325 vccd1 _0893_.CLK a_26523_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10326 vccd1 _0837_.A1 a_8393_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X10327 vssd1 a_21683_9117# a_21851_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10328 a_25639_23439# a_24775_23445# a_25382_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10329 a_13395_5515# _0582_.A a_13309_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10330 a_10367_11471# a_9503_11477# a_10110_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10331 a_4422_1501# a_3983_1135# a_4337_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10334 vccd1 a_10183_9295# a_10351_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10335 a_10183_9295# a_9485_9301# a_9926_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10336 a_17769_3311# _1041_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10337 vssd1 _0888_.CLK a_6651_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10338 a_27847_25437# a_27149_25071# a_27590_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10339 _1019_.D a_20195_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10340 a_20249_21269# a_20083_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10341 vssd1 _0445_.A a_10948_21813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X10342 a_20430_22351# a_20157_22357# a_20345_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10343 a_12257_7439# _0899_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X10344 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_14740_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10345 vssd1 a_9284_10901# _0685_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10346 _0776_.A2 a_7623_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10350 a_16439_4765# a_15575_4399# a_16182_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10351 a_14265_5321# a_13275_4949# a_14139_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10352 a_6651_12672# _0685_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10354 a_10037_11471# a_9503_11477# a_9942_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10356 vccd1 _0441_.B a_11067_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X10357 vccd1 _0472_.X a_12447_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X10358 _0932_.D a_21115_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10359 a_27456_8751# a_27057_8751# a_27330_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10360 a_11711_24527# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10361 vssd1 _1019_.CLK a_18243_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10362 a_19877_9839# _0940_.Q a_19439_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10363 vccd1 a_4863_23413# _0814_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X10364 vccd1 _0734_.A2 a_5737_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10365 _1012_.D a_25715_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10366 vccd1 a_23047_15797# a_22963_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10367 vccd1 a_27847_3677# a_28015_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10368 a_4984_26703# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10369 _0847_.A1 clkbuf_1_0__f_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X10370 a_4589_17999# _0722_.C _0798_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10372 a_20813_1999# _1041_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X10373 _0506_.X a_22659_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10374 a_2962_14735# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X10375 a_2949_27247# a_1959_27247# a_2823_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10377 a_27931_5853# a_27149_5487# a_27847_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10378 vssd1 a_2626_9269# _0835_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X10379 a_22365_12265# _0892_.D a_22281_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10380 vccd1 a_2807_4667# a_2723_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10382 a_14747_6031# _0516_.B1 a_14829_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10383 _0698_.A2_N _0696_.A1 a_2689_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
D5 vssd1 ANTENNA_7.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X10384 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10968_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10385 vccd1 _0925_.D a_18088_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10386 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12355_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10387 a_15657_19453# _0840_.A1 a_15575_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10388 a_1766_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X10389 vssd1 a_5031_1679# a_5199_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10392 vccd1 _0778_.A2 a_6651_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10393 a_18232_13967# _0925_.D a_17657_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X10394 a_10202_13621# a_10034_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10395 vccd1 a_23047_1653# a_22963_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10396 vssd1 _0614_.A a_15483_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X10397 vccd1 a_25707_25321# _0854_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10398 vccd1 a_25623_22075# a_25539_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10399 a_21279_6825# _0630_.A2 a_21361_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10400 vssd1 a_20598_22325# a_20556_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10401 _0758_.A2 _0756_.A2 a_5721_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X10402 a_13521_6575# _0604_.B a_13449_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10403 a_20161_7663# _1029_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10404 vccd1 _0860_.A a_12622_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X10405 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10406 vssd1 a_22419_22173# a_22587_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10408 vccd1 fanout13.A _0828_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10409 vssd1 _0845_.C1 _0835_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10410 a_10313_24847# _0837_.A1 _0819_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X10411 _0632_.B a_24887_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10412 a_7271_7663# _0656_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112125 ps=0.995 w=0.65 l=0.15
X10414 vccd1 a_23691_9019# a_23607_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10415 a_25214_23439# a_24941_23445# a_25129_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10416 vssd1 _0590_.B2 a_20180_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X10417 a_8914_7093# a_8746_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10418 vccd1 a_3298_17143# _0812_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X10419 _0512_.X a_19195_18337# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X10421 _0938_.Q a_20471_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10426 vssd1 temp1.dcdc.Z a_5078_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10427 a_10140_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10428 vssd1 a_15871_2491# a_15829_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10429 a_7850_11249# a_7801_11079# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X10430 _0582_.C a_14729_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X10431 a_14875_15325# _1075_.Q a_14775_15325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10432 _0586_.B2 a_8971_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10433 a_1591_21807# _0814_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10434 vssd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10436 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI a_14260_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10437 vssd1 a_22622_20149# a_22580_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10438 a_12207_15645# a_11509_15279# a_11950_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10440 vssd1 _0735_.A2 a_9583_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X10445 vssd1 _0888_.CLK a_8307_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10446 vssd1 _0494_.X a_19593_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10447 a_1945_8751# _0875_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10448 a_15236_10383# _0487_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10450 a_12622_24233# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10451 vccd1 a_25842_4917# a_25769_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10453 vccd1 a_25842_16885# a_25769_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10454 vssd1 _0893_.CLK a_22383_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10456 vssd1 fanout10.A a_9871_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10457 a_14651_24527# _0861_.B1 a_14433_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X10458 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_5639_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10459 a_2823_2589# a_1959_2223# a_2566_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10460 a_13069_7663# _0646_.A1 a_12631_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10461 vssd1 a_11490_3423# a_11448_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10462 _0905_.Q a_5383_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10463 a_22143_2589# a_21445_2223# a_21886_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10464 a_25217_13469# a_24683_13103# a_25122_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10465 a_2524_27247# a_2125_27247# a_2398_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10468 a_25213_18319# _0998_.Q a_24867_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X10469 a_20246_8029# a_19807_7663# a_20161_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10470 vccd1 a_25163_13621# a_25079_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10471 temp1.capload\[5\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10472 a_8392_26159# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10473 vssd1 a_9503_19087# _0471_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10474 a_22549_19093# a_22383_19093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10478 a_27337_14191# _1012_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10482 a_10386_2741# a_10218_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10483 a_16981_5281# _0582_.A a_16895_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10484 a_26225_21641# a_25235_21269# a_26099_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10485 _0888_.CLK a_2787_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X10486 vssd1 _0815_.Y a_14011_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10487 a_20997_16617# _0564_.C a_20901_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10488 a_12716_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10489 a_4356_23983# _0774_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10490 a_13054_15797# a_12886_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10491 a_14829_6351# _0671_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X10493 _0606_.X a_16863_14848# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10494 vccd1 _0959_.CLK a_14747_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10496 a_16757_21807# _0933_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10497 vccd1 _0483_.X a_20761_9633# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10498 a_4149_2223# a_3983_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10499 a_27513_10703# _0893_.Q a_27167_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X10500 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10501 a_27149_17455# a_26983_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10502 a_4548_1135# a_4149_1135# a_4422_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10503 a_6741_15055# _0794_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X10504 _1042_.Q a_18447_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10505 a_3028_14165# _0456_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10506 _0674_.C1 a_11987_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X10507 vssd1 _0588_.X a_19439_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10509 a_25198_21919# a_25030_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10510 a_4167_17999# _0722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10511 a_2114_1653# a_2464_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X10512 vccd1 _0995_.CLK a_15667_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X10513 vssd1 a_21115_21237# a_21073_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10514 a_25750_12127# a_25582_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10515 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15016_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10516 _0638_.X a_18059_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10518 vssd1 _0768_.A1 a_5692_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X10519 vssd1 _0975_.CLK a_22015_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10520 a_16032_6351# _0670_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X10521 a_7642_4765# a_7369_4399# a_7557_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10522 _0694_.A2 _0680_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X10523 _0714_.B1 _0735_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10524 vccd1 _0583_.A a_22751_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10525 vssd1 a_27498_8863# a_27456_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10526 a_10504_18543# a_10055_18543# a_10202_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10527 _0961_.D a_10903_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10528 a_9945_23759# _0835_.A1 _0816_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X10529 vccd1 a_2686_23439# _0844_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10530 _0931_.CLK a_18611_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10531 a_10872_25935# _0847_.A2 _0847_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X10532 vccd1 _0511_.D a_14729_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X10533 a_16293_7913# _1059_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X10534 a_16904_24643# _0860_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10535 a_25750_3423# a_25582_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10536 a_14629_14191# _1076_.Q a_14557_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X10539 vccd1 a_25455_4765# a_25623_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10541 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10542 a_14011_7235# _0544_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10543 vssd1 _0824_.Y a_13183_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10544 a_17405_2473# _0516_.B1 a_17489_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10545 a_13169_9295# _1026_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10546 vccd1 _0444_.A a_2051_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10547 a_17029_10389# a_16863_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10548 a_15879_27791# a_15097_27797# a_15795_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10549 a_2125_3311# a_1959_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10550 vccd1 a_13882_4917# a_13809_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10552 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10553 a_15054_10383# _0612_.X a_14805_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10554 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R26 vssd1 temp1.capload\[12\].cap_42.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10555 vccd1 a_9227_17455# _0995_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10556 vssd1 fanout24.A a_25235_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10558 a_10689_21853# _0850_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10562 vssd1 _1030_.CLK a_20175_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10564 a_4589_17999# _0722_.B a_4167_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10565 a_4403_25589# _0840_.A0 a_4612_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X10566 a_2405_25071# _0839_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10567 a_7197_20969# _0869_.B1 _0869_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10571 a_22971_2767# a_22273_2773# a_22714_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10572 a_23119_10089# _0487_.X a_23201_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10575 a_10533_18776# _1075_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X10576 vssd1 a_2752_1897# a_2762_1801# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10577 a_18221_10089# _0616_.X a_18148_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X10578 vccd1 a_17895_2741# a_17811_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10579 vccd1 _0860_.A a_16029_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X10580 vssd1 _0582_.C a_20237_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10583 _0910_.Q a_3727_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10584 _0749_.A1 _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10585 vccd1 a_27590_15391# a_27517_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10586 vssd1 _0725_.A a_3891_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X10588 a_4132_17429# a_3983_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X10589 io_out[4] _0752_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X10590 a_2464_1653# a_2762_1801# a_2710_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09135 ps=0.855 w=0.42 l=0.15
X10591 a_5510_8207# _0694_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X10592 _0521_.A a_13459_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10595 vssd1 a_22990_3423# a_22948_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10596 vssd1 _0917_.CLK a_12815_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10597 _0936_.Q a_8695_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10599 _0758_.B1 _0685_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10600 vccd1 a_3270_2741# _0850_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10601 _0573_.B a_26267_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10602 vssd1 _0456_.A a_5089_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X10603 vssd1 _0602_.A a_18703_12567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10604 vccd1 a_2991_27515# _1076_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10606 vccd1 a_20471_17723# a_20387_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10607 _0466_.A a_1591_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10608 a_2030_5853# a_1757_5487# a_1945_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10610 vccd1 _0472_.X a_6559_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10612 vccd1 fanout27.A a_22659_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10613 a_6549_9001# _0656_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X10614 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10616 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10617 a_14342_19061# a_14174_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10618 a_20372_7663# a_19973_7663# a_20246_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10621 vccd1 _0850_.A a_7602_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10623 a_25125_15645# a_24591_15279# a_25030_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10624 a_9999_1501# a_9135_1135# a_9742_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10625 a_11597_5487# _0907_.Q a_11251_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X10626 a_12701_6409# a_11711_6037# a_12575_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10627 a_21442_13469# a_21169_13103# a_21357_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10629 a_25842_14709# a_25674_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10632 a_18325_9001# _0667_.B1 a_18409_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10633 vssd1 a_18125_18517# _0559_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X10634 vccd1 a_9171_7119# a_9339_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10636 a_7376_20495# _0784_.A1 a_7073_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X10637 vssd1 _1033_.CLK a_24867_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10638 a_17217_2767# _0622_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10640 a_18148_8527# _0648_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X10641 a_27249_11471# _0619_.B2 a_27167_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10642 _0563_.B1 a_20299_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X10643 vccd1 a_5078_30511# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10644 vccd1 a_8067_4765# a_8235_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10646 a_2217_25071# a_2051_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10647 a_10861_2223# a_9871_2223# a_10735_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10648 _0807_.A a_2623_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10650 a_10212_31055# a_9963_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10651 _0745_.A2 a_4040_10901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X10652 vccd1 _0521_.A a_16127_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10653 vssd1 clkbuf_1_0__f_temp1.i_precharge_n.A a_1674_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10654 vccd1 a_22449_15253# _0561_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X10655 vssd1 a_4590_1247# a_4548_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10656 a_20982_4765# a_20543_4399# a_20897_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10657 a_25674_14735# a_25401_14741# a_25589_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10659 a_4255_12265# _0776_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10661 vccd1 a_6612_8181# _0710_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X10662 a_17289_13249# _0602_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X10663 a_14457_20175# _0919_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10664 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10665 vccd1 a_26267_19899# a_26183_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10666 a_6559_16911# _0836_.A a_6809_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10668 a_19521_4649# _0630_.A2 a_19605_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10669 vssd1 ANTENNA_7.DIODE a_4811_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10670 vccd1 a_16607_4667# a_16523_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10671 a_7841_15279# _0760_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X10672 vccd1 a_11030_11039# a_10957_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10674 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8767_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10675 a_11782_21085# a_11343_20719# a_11697_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10676 vssd1 a_20195_6005# a_20153_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10677 vssd1 a_8159_6031# a_8327_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10678 vccd1 _0506_.A2 a_20349_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10679 _0546_.B1 a_9895_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X10681 a_6831_22351# _0861_.B1 a_6613_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X10682 a_21073_21641# a_20083_21269# a_20947_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10683 a_14683_19087# a_13901_19093# a_14599_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10684 vssd1 _0722_.B a_2852_15285# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X10685 vssd1 a_8327_6005# a_8285_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10686 a_12629_23145# a_12355_22901# a_12547_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10687 vssd1 a_18611_14735# _0662_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X10688 vccd1 a_1674_32143# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10690 vssd1 a_24059_26677# a_24017_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10691 a_8611_21263# a_7829_21269# a_8527_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10692 a_18308_27497# a_18059_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10693 a_2823_2589# a_2125_2223# a_2566_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10695 vccd1 _1033_.CLK a_25235_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10696 _1021_.Q a_22035_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10697 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10698 vccd1 a_15151_10205# a_15319_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10699 a_24021_22357# a_23855_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10700 a_4137_18543# _0722_.B a_4065_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10701 a_4712_16617# _0877_.A2 _0877_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X10702 vccd1 _0502_.X a_18519_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
R27 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10703 vssd1 a_26175_12283# a_26133_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10705 _0565_.B1 _0512_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10706 vccd1 _0752_.Y io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10707 _0836_.A a_8031_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X10708 vssd1 io_in[6] a_1591_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10709 vccd1 clkbuf_1_0__f_io_in[0].X a_1775_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10711 vssd1 a_16607_14459# a_16565_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10712 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10714 a_10325_15529# _0836_.A a_10229_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10715 vssd1 a_20046_15391# a_20004_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10716 vccd1 _0549_.X a_15365_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10717 vssd1 _1053_.CLK a_14471_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10718 _0798_.A2 _0722_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10719 vccd1 a_21683_9117# a_21851_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10720 vccd1 _0685_.B a_6559_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10721 a_12610_21263# a_12171_21269# a_12525_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10722 _0864_.Y _0863_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10725 a_16101_18517# _0667_.B1 a_16258_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X10726 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10727 a_16573_26159# _1052_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10729 _0994_.Q a_26635_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10730 a_6423_8903# _0657_.X a_6663_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X10732 vccd1 a_27111_18909# a_27279_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10733 a_24849_13103# a_24683_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10735 vssd1 a_23507_20987# a_23465_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10738 _0531_.X a_20635_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X10739 a_14825_17999# _1056_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10740 a_17727_2767# a_17029_2773# a_17470_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10741 vccd1 a_26099_7119# a_26267_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10743 a_10968_30287# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10744 _0998_.Q a_28015_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10748 a_19885_2767# _0970_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10749 a_10073_26133# _0819_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X10750 a_16264_18543# _0577_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X10751 vssd1 a_25455_4765# a_25623_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10752 a_9765_4399# _0959_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10753 vccd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10754 vccd1 a_19015_20175# a_19183_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10755 a_23385_14013# _0583_.A a_23303_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10757 a_9189_18517# _0797_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X10758 vssd1 _0456_.B a_4864_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X10759 vssd1 _0474_.X _0565_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10761 a_2686_31055# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10762 vccd1 a_25198_15391# a_25125_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10763 a_5353_10089# _0776_.A2 _0756_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X10764 a_15553_23817# a_14563_23445# a_15427_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10765 a_13054_15797# a_12886_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10766 vccd1 _0505_.A2 a_22741_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10768 vssd1 a_19015_20175# a_19183_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10769 vssd1 _0807_.B _0882_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10770 a_13855_10383# a_13073_10389# a_13771_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10771 a_20671_14735# a_19807_14741# a_20414_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10772 vccd1 a_2991_2491# a_2907_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10773 a_11764_20149# _0850_.A a_11987_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X10774 vssd1 _0931_.CLK a_20819_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10776 vccd1 _0710_.A1 a_5325_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X10777 a_13679_9295# a_12815_9301# a_13422_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10778 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X10779 vccd1 a_26175_10107# a_26091_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10780 a_5173_20719# a_4981_21024# _0870_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X10781 vssd1 a_20414_7775# a_20372_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10782 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10783 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10784 vssd1 a_24167_9295# a_24335_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10785 a_20395_2767# a_19697_2773# a_20138_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10786 a_22185_26159# _1019_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10787 vssd1 _0893_.CLK a_25235_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10788 a_12061_3861# a_11895_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10789 a_15115_5059# _0556_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X10790 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10212_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10793 a_20989_20719# _1048_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10794 a_22833_7913# _0618_.C1 a_22751_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10795 vccd1 a_16347_21085# a_16515_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10796 vccd1 _0935_.CLK a_14103_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10798 a_15695_14735# a_14913_14741# a_15611_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10799 vssd1 a_15151_12381# a_15319_12283# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10800 a_20341_14735# a_19807_14741# a_20246_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10801 a_10073_26133# _0819_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X10803 vccd1 a_8176_19061# _0765_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X10804 _0621_.X a_23303_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X10807 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10808 a_17121_1685# a_16955_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10809 vccd1 _0880_.A1 a_9588_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X10810 a_4015_5515# _0695_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10812 a_9769_19881# _0751_.B2 a_9687_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10813 a_20303_15645# a_19439_15279# a_20046_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10814 a_11237_3311# _0543_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10815 a_25658_7775# a_25490_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10816 a_22741_11177# _0505_.X a_22659_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10817 a_2125_27247# a_1959_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10819 vssd1 _0667_.X a_18059_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10821 vccd1 _0922_.CLK a_9135_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X10823 vssd1 a_13939_10357# a_13897_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10825 vccd1 a_27847_16733# a_28015_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10826 a_10225_2223# _0637_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10827 vccd1 a_2198_5599# a_2125_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10830 a_24803_22351# a_24021_22357# a_24719_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10832 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10833 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_13360_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10834 a_22503_22173# a_21721_21807# a_22419_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10835 _0585_.X a_19439_12675# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X10836 a_11897_12265# _0474_.X a_11815_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10837 vssd1 _0444_.A a_2419_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10838 vccd1 a_13367_17999# _0866_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10839 vccd1 a_7810_4511# a_7737_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10840 vccd1 a_13146_1653# a_13073_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10841 vccd1 a_12631_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10843 vccd1 a_9815_16911# a_9983_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10844 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10845 a_27517_25437# a_26983_25071# a_27422_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10846 a_2686_23439# clkbuf_1_1__f__0390_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X10847 vssd1 _0471_.X a_10147_15529# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X10848 vssd1 a_22990_19061# a_22948_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10849 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_11980_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10850 vssd1 _0832_.A a_4075_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10851 a_27931_24349# a_27149_23983# a_27847_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10852 a_9117_16917# a_8951_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10856 a_19602_26703# a_19329_26709# a_19517_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10857 a_11987_2473# _0532_.A2 a_12069_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10858 vssd1 _0801_.X a_13367_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X10860 _0751_.B2 _0798_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10861 vccd1 _0511_.D a_14603_15325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X10862 a_14821_10205# a_14287_9839# a_14726_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10863 a_20981_10703# _0531_.A1 a_20635_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X10866 vssd1 _0959_.CLK a_10883_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10867 _0517_.D a_21647_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10868 a_2198_8863# a_2030_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10870 a_23469_6037# a_23303_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10872 a_11987_20495# _0847_.A2 a_11893_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X10874 a_22622_15797# a_22454_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10875 vccd1 fanout23.X a_25235_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10876 a_10478_2335# a_10310_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10877 _0674_.A1 a_9615_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10878 a_9171_7119# a_8307_7125# a_8914_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10879 a_27245_8751# _0647_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10880 a_27337_21807# _0998_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10881 a_4333_1685# a_4167_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10882 vssd1 a_8067_4765# a_8235_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10884 a_27847_12381# a_26983_12015# a_27590_12127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10886 a_20429_17455# a_19439_17455# a_20303_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10887 a_9761_13653# a_9595_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10888 _0807_.A a_2623_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10889 vssd1 a_14621_8897# _0614_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X10890 a_9942_21263# a_9669_21269# a_9857_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10891 a_16983_16395# _0521_.A a_16897_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10892 _0803_.X a_6283_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10894 vccd1 a_1639_7338# input2.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10895 vssd1 _0908_.CLK a_5455_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10896 a_19697_2773# a_19531_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10897 a_8832_27791# a_8583_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10898 vccd1 _0558_.X a_21069_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10899 vccd1 a_9613_25045# a_9643_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10902 a_13073_10389# a_12907_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10903 a_14710_20149# a_14542_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10904 a_25401_19631# a_25235_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10905 a_22454_15823# a_22181_15829# a_22369_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10906 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10908 a_25037_13103# _1011_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10909 vssd1 _0680_.Y _0694_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.105625 ps=0.975 w=0.65 l=0.15
X10911 a_9853_22357# a_9687_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10912 vccd1 a_12375_20987# a_12291_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10913 a_4065_14237# _0460_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10914 _0648_.X a_23303_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X10915 _0735_.A2 a_7111_13655# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10916 vssd1 _0440_.C _0445_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10917 vssd1 _0847_.A3 a_10313_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X10918 a_25309_3311# a_25143_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10920 vccd1 a_17727_10383# a_17895_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10921 a_5547_25615# _0845_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10922 _0939_.Q a_25623_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10923 _0860_.A a_2114_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X10924 vccd1 a_1674_26159# clkbuf_1_0__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10926 a_12701_11849# a_11711_11477# a_12575_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10927 a_24462_20149# a_24294_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10929 vccd1 a_22035_24251# a_21951_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10930 a_27237_18543# a_26247_18543# a_27111_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10931 a_10876_32463# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10932 vccd1 a_4663_3855# a_4831_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10933 vccd1 a_12207_18909# a_12375_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10934 a_26099_19087# a_25401_19093# a_25842_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10935 vssd1 a_17654_17567# a_17612_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10938 vccd1 _0722_.A a_2051_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10940 vssd1 _1015_.CLK a_26891_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10942 a_10643_2767# a_9779_2773# a_10386_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10943 a_1591_26703# _1081_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10944 a_4338_10089# _0699_.A0 a_4035_9813# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X10947 a_11697_18543# _0918_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10948 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10948_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10950 vccd1 _0502_.X a_19471_6603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10951 a_14641_7663# _1027_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10952 a_12777_16885# _0798_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X10953 a_12318_8181# a_12150_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10954 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_12065_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X10955 _0749_.B2 _0812_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10956 vccd1 a_22971_2767# a_23139_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10957 a_26578_11039# a_26410_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10959 vssd1 _0570_.X a_23361_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X10960 vccd1 a_26267_25589# a_26183_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10961 vccd1 a_20414_14709# a_20341_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10962 a_27149_9839# a_26983_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10964 _0988_.D a_12375_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10965 vssd1 a_17838_23007# a_17796_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10966 a_14483_15279# _1076_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X10967 a_25030_5853# a_24591_5487# a_24945_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10971 vssd1 a_10386_2741# a_10344_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10972 a_10386_1653# a_10218_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10973 a_2125_5853# a_1591_5487# a_2030_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10975 a_11842_25321# _0829_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X10976 a_7348_17973# _0739_.B1 a_7477_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X10977 vssd1 _0768_.B1 a_7900_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X10978 a_5491_4943# a_4793_4949# a_5234_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10979 a_27422_12381# a_27149_12015# a_27337_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10981 a_12613_15829# a_12447_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10982 a_24738_13621# a_24570_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10983 a_21265_18543# _0991_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10984 a_14453_9839# a_14287_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10985 a_19360_14025# a_18961_13653# a_19234_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10986 a_26053_13647# _0928_.D a_25971_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10987 _0976_.Q a_28015_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10988 a_17946_1501# a_17507_1135# a_17861_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10991 a_22549_3311# a_22383_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10992 a_13073_1679# a_12539_1685# a_12978_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10993 vssd1 a_8859_17999# _0472_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X10995 vccd1 a_20046_15391# a_19973_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10996 vssd1 _0922_.CLK a_9135_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10997 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10998 a_13345_4399# a_12355_4399# a_13219_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10999 a_10948_28879# a_10699_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11000 vccd1 _0808_.A a_8123_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11001 a_12150_13647# a_11711_13653# a_12065_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11003 a_14726_8029# a_14287_7663# a_14641_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11004 vccd1 fanout27.A a_21003_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11005 vssd1 _0577_.C a_12015_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11006 a_6682_11587# _0745_.A3 a_6600_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11007 a_24570_13647# a_24297_13653# a_24485_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11008 a_13261_22351# _1054_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11009 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11010 vssd1 _0513_.X a_15879_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11011 vssd1 _0444_.A a_2051_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11012 a_18125_18517# _0584_.A2 a_18282_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X11013 vssd1 _0975_.CLK a_22383_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11014 a_4988_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11015 vssd1 _0814_.A2 a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11016 a_11950_20831# a_11782_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11017 vccd1 a_16055_16635# a_15971_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11019 vccd1 _0758_.A2 a_6473_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11020 a_6516_18695# a_6646_18865# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X11022 a_15101_14735# _0924_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11025 vccd1 a_3891_21263# _0814_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11026 _0594_.D a_19899_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X11027 vccd1 a_14894_9951# a_14821_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11028 a_22377_10499# _0651_.C a_22281_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11029 a_4337_1135# _0849_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11030 vccd1 _0972_.CLK a_15575_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11031 _0558_.A2 a_21127_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11032 temp1.capload\[4\].cap.Y temp1.capload\[4\].cap.A a_15661_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11033 a_22438_26271# a_22270_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11034 _1027_.Q a_13847_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11035 a_22469_12879# _0891_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11036 a_10643_1679# a_9945_1685# a_10386_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11037 vccd1 _0472_.X _0678_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11039 a_10576_18543# a_10533_18776# a_10504_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X11040 a_15093_6351# _0916_.D a_14747_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X11041 a_17911_17821# a_17047_17455# a_17654_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11042 a_10147_15823# _0472_.X a_10397_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11043 a_2398_1501# a_1959_1135# a_2313_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11044 a_11877_8213# a_11711_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11045 _0675_.C a_16863_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11046 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X11048 a_10367_11471# a_9669_11477# a_10110_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11049 a_1591_25615# _0845_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11051 a_18371_11293# a_17507_10927# a_18114_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11052 a_23523_4765# a_22825_4399# a_23266_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11053 a_4340_12015# _0745_.A2 a_4037_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X11055 _0848_.X a_12547_23145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X11056 a_10217_7663# a_9227_7663# a_10091_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11057 vssd1 a_2658_28447# a_2616_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11058 a_26225_1135# a_25235_1135# a_26099_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11060 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A a_8832_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11061 a_2776_2767# a_2235_2773# a_2683_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X11062 a_4422_2589# a_4149_2223# a_4337_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11063 a_20214_16911# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11064 vccd1 _0572_.A2 a_22097_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X11065 vccd1 _0572_.A2 a_24673_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X11067 vccd1 _0888_.CLK a_4627_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11068 _0863_.A1 a_15575_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11069 vccd1 _0583_.A a_17231_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11070 _0544_.D a_14839_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X11071 a_17581_17821# a_17047_17455# a_17486_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11072 a_21384_19631# a_20985_19631# a_21258_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11074 a_27590_24095# a_27422_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11075 a_18041_11293# a_17507_10927# a_17946_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11077 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_8215_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11079 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11080 a_21077_18543# a_20911_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11081 vssd1 _0735_.A2 a_12711_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11082 _0645_.B2 a_15963_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11084 a_4238_3855# a_3965_3861# a_4153_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11085 vccd1 a_3799_11471# _0861_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11087 a_22369_20175# _1022_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11088 vccd1 a_5601_18517# _0784_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11090 vssd1 a_28015_10107# a_27973_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11091 vccd1 _1046_.D a_21134_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X11092 a_10055_24527# _0837_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11094 a_15795_1679# a_14931_1685# a_15538_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11097 a_12532_29199# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11098 a_2631_3855# a_1849_3861# a_2547_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11099 vssd1 temp1.dcdc.Z a_5078_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11100 _0828_.Y fanout13.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11101 _0930_.Q a_25623_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11104 vccd1 _0527_.X a_15975_10721# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X11105 vssd1 a_4811_10383# _0845_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11107 vccd1 _0964_.CLK a_25051_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11109 a_8546_1653# a_8378_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11110 a_21867_13469# a_21169_13103# a_21610_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11111 vssd1 _1015_.CLK a_25143_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11115 a_16553_15425# _0577_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11116 a_8017_21263# _0935_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11117 vccd1 a_25623_16635# a_25539_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11118 vssd1 a_15538_1653# a_15496_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11119 a_25401_19093# a_25235_19093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11120 vssd1 _0972_.CLK a_16863_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11121 a_2566_3423# a_2398_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11122 a_12333_18543# a_11343_18543# a_12207_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11123 a_20782_5599# a_20614_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11124 a_8392_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11125 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A a_8392_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11126 vccd1 a_13847_9269# a_13763_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11127 vccd1 fanout10.A a_10791_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11128 _0952_.Q a_14307_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11131 vccd1 _0613_.A1 a_15236_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X11132 a_15844_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11133 a_4337_26159# _0843_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11134 a_25156_5487# a_24757_5487# a_25030_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11135 vccd1 _0577_.C a_14287_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11136 a_17313_19453# _0583_.A a_17231_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11137 a_27571_6941# a_26707_6575# a_27314_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11140 vssd1 a_12318_8181# a_12276_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
R28 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11141 vssd1 _0819_.S temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11142 vssd1 _0994_.CLK a_24591_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R29 temp1.capload\[14\].cap_44.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11144 vssd1 _0814_.A2 a_4337_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X11145 vccd1 _0472_.X _0838_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11146 vccd1 _0835_.A1 a_11067_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X11147 a_4356_23983# _0814_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11148 a_18427_2473# _0594_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11149 a_2915_28701# a_2051_28335# a_2658_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11150 a_21150_4511# a_20982_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11151 vccd1 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_1766_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11152 vccd1 a_15170_3829# a_15097_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11153 vssd1 _0893_.CLK a_24131_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11155 a_10791_17705# _0471_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11156 vssd1 a_6795_14343# _0779_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X11157 _0558_.X a_24867_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X11158 a_17725_15073# _0521_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11159 a_20161_7663# _1029_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11160 _0676_.B a_15391_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X11161 _0546_.B1 a_9895_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11162 vssd1 a_27003_11195# a_26961_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11163 a_26183_4943# a_25401_4949# a_26099_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11164 a_19439_9001# _0517_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11165 vccd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11166 vssd1 _0764_.A1 a_6600_26409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11167 a_11895_1385# _0850_.Y a_11895_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X11168 a_2585_28701# a_2051_28335# a_2490_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11170 a_14852_7663# a_14453_7663# a_14726_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11171 a_9791_12015# _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X11172 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X11173 vccd1 _0814_.A2 a_4439_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X11174 vssd1 a_8079_28500# _0821_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11175 vssd1 a_5015_2491# _0829_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11177 vssd1 _0619_.B1 a_23465_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X11178 vssd1 a_13771_22351# a_13939_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11179 vccd1 a_10202_18517# _0577_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X11180 _0642_.D_N _0638_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.24 as=0.12025 ps=1.02 w=0.65 l=0.15
X11181 a_11877_13653# a_11711_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11182 vssd1 _0546_.X a_10779_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11183 _0660_.X a_25695_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X11185 a_18505_4943# _0543_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11187 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11188 a_4581_25847# _0844_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X11189 _1053_.CLK a_8307_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11190 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11192 vccd1 _0995_.CLK a_21831_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11193 a_6713_19631# _0807_.B a_6641_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11194 _0797_.B1 a_6876_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X11195 a_20993_1135# _1040_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11196 a_7182_3855# a_6909_3861# a_7097_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11197 a_9687_23439# _0835_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11198 vccd1 _0791_.A3 a_4035_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X11199 a_2125_2223# a_1959_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11202 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A a_5078_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11203 a_2524_1135# a_2125_1135# a_2398_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11204 a_5417_20149# _0812_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X11205 a_27973_16367# a_26983_16367# a_27847_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11207 a_16581_23983# _0860_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11208 vccd1 a_17654_17567# a_17581_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11210 vccd1 a_26927_21085# a_27095_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11211 vssd1 _0835_.A1 a_11895_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11212 vccd1 clkbuf_1_0__f_io_in[0].X a_1591_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11213 a_4931_28701# a_4149_28335# a_4847_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11215 a_22822_14557# a_22549_14191# a_22737_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11217 a_19617_9001# _0506_.X a_19521_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11219 vssd1 a_1639_7828# input3.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11220 vccd1 a_18114_11039# a_18041_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11221 a_22921_7119# _1045_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11222 vssd1 _0711_.A a_5091_12021# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11223 a_18409_21269# a_18243_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11224 vssd1 _0680_.Y a_6423_8903# vssd1 sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X11225 a_25674_19997# a_25401_19631# a_25589_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11226 vccd1 _0655_.X _0707_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11227 a_23792_13353# _0569_.X a_23690_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11228 a_12962_4511# a_12794_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11231 vssd1 a_7939_19631# _0833_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X11232 a_9742_5599# a_9574_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11233 vssd1 _0860_.B a_16115_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11234 _1061_.D a_19275_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11235 a_15278_2589# a_15005_2223# a_15193_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11237 a_15088_29967# a_14839_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11238 temp1.capload\[0\].cap.Y temp1.capload\[0\].cap.A a_16305_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11239 a_10397_15529# _0472_.X a_10325_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11240 vssd1 a_15963_27765# a_15921_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11242 vccd1 _0908_.CLK a_6743_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11243 _0726_.X a_6559_23552# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11244 a_3028_14165# a_2879_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11245 a_15473_8323# _0675_.D a_15391_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11248 a_11041_17705# _0833_.A a_11238_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11249 a_12759_3855# a_11895_3861# a_12502_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11250 _0710_.B1 a_4015_5515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
R30 vccd1 temp1.capload\[1\].cap_46.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11252 a_10275_4765# a_9577_4399# a_10018_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11253 a_25401_16917# a_25235_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11254 a_14603_15325# a_14287_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11255 a_14223_4943# a_13441_4949# a_14139_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11256 a_3302_4917# a_3134_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11257 vssd1 a_7037_29177# a_6971_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X11258 vccd1 a_14599_19087# a_14767_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11259 a_13705_14013# _0936_.Q a_13633_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11260 a_19329_3861# a_19163_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11261 vssd1 _0843_.B _0843_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11262 vssd1 a_27463_4667# a_27421_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11263 _0621_.B2 a_26083_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11268 vccd1 temp1.capload\[1\].cap_46.LO temp1.capload\[1\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11269 vssd1 a_28015_24251# a_27973_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11270 vssd1 _0639_.X _0642_.D_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.125125 ps=1.035 w=0.65 l=0.15
X11271 vccd1 a_10811_2741# a_10727_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11272 a_24068_12559# _0576_.B1 a_23966_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11273 _1000_.Q a_26267_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11274 a_23105_8207# _0590_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11276 a_9447_3855# a_8583_3861# a_9190_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11278 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11279 a_25842_3829# a_25674_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11280 a_17854_3677# a_17415_3311# a_17769_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11281 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11282 a_15151_12381# a_14287_12015# a_14894_12127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11283 a_7900_14165# _0768_.C1 a_8292_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X11285 a_15887_16733# a_15189_16367# a_15630_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11286 a_23457_14013# _1012_.Q a_23385_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11287 a_6612_14709# _0778_.B1 a_6835_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X11288 _1015_.CLK a_23763_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X11289 vssd1 a_12502_3829# a_12460_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11290 _0506_.A1 a_24335_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11291 vccd1 _0658_.B1 a_19697_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X11293 a_20004_17455# a_19605_17455# a_19878_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11294 vssd1 a_24335_9269# a_24293_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11296 a_2125_27247# a_1959_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11297 _0487_.X a_17725_15073# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X11299 vssd1 a_25198_5599# a_25156_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11300 a_12713_7913# _0522_.B1 a_12797_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11301 a_25198_15391# a_25030_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11302 a_10777_10927# _0588_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11304 vssd1 _0833_.A _0518_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11305 a_27337_2223# _0665_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11306 _0938_.Q a_20471_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11307 a_22741_11471# _0992_.D a_22659_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11309 a_5541_29199# _0809_.B2 a_5323_29111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X11310 a_27337_25071# _0998_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11311 a_15097_27797# a_14931_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11312 vccd1 _0840_.A1 a_12625_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X11313 vssd1 a_9190_3829# a_9148_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11315 _0713_.A3 a_6600_11587# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X11316 vccd1 _0994_.CLK a_24591_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11318 a_7357_9661# _0685_.B a_7285_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11319 a_21242_20831# a_21074_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11320 vssd1 a_3983_3311# ANTENNA_7.DIODE vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11321 vccd1 a_2658_28447# a_2585_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11322 _0569_.X a_22383_14848# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
R31 temp1.capload\[2\].cap_47.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11324 vssd1 fanout37.A a_4259_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X11325 _0546_.A2 _0466_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11326 a_14641_9839# _0961_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11327 vssd1 a_11619_29423# fanout10.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11328 a_22546_2767# a_22107_2773# a_22461_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11329 a_16305_7663# _0549_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11330 a_3302_4917# a_3134_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11332 _0505_.A2 a_19471_6603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X11333 vssd1 a_14894_7775# a_14852_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11334 a_25582_10205# a_25309_9839# a_25497_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11336 _0845_.A2 a_2686_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11337 a_7331_6941# a_6633_6575# a_7074_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11338 vssd1 _1053_.CLK a_10791_16919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11339 a_10133_2767# _0673_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11340 a_20479_2767# a_19697_2773# a_20395_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11341 vccd1 a_3523_6039# fanout37.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11342 _0575_.B a_25623_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11343 a_2214_4765# a_1941_4399# a_2129_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11344 vccd1 _0917_.CLK a_12907_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11346 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_18236_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11348 _0652_.C a_12631_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X11349 vccd1 a_7939_19631# _0833_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11351 vssd1 a_16553_15425# _0580_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X11352 a_25842_3829# a_25674_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11353 vssd1 clkbuf_1_1__f_net57.A a_1674_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11354 a_6809_16911# _0836_.A a_6559_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11355 a_20897_4399# _0649_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11356 vccd1 _0662_.A1 a_11897_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X11357 _0768_.A1 a_3523_13655# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X11358 a_23013_4399# _0548_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11359 vssd1 _1033_.CLK a_26983_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11360 a_16842_22173# a_16403_21807# a_16757_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11361 a_24845_20553# a_23855_20181# a_24719_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11362 a_12479_5515# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11363 a_21407_3677# a_20709_3311# a_21150_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11364 a_24297_13653# a_24131_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11366 vccd1 a_22817_18517# _0662_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X11367 a_25769_7119# a_25235_7125# a_25674_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11368 vssd1 a_1674_26159# clkbuf_1_0__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11369 a_3424_19087# _0872_.A2 _0872_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X11370 vssd1 a_2566_1247# a_2524_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11371 a_14599_19087# a_13735_19093# a_14342_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11372 a_1757_6575# a_1591_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11373 a_18731_7457# _0582_.A a_18645_7457# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11374 a_18689_25615# _1061_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11375 a_8527_21263# a_7663_21269# a_8270_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11376 vssd1 a_13054_15797# a_13012_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11377 vccd1 a_4590_2335# a_4517_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11378 a_19981_1135# _0970_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11379 vssd1 a_21867_24349# a_22035_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11380 vccd1 a_15611_14735# a_15779_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11382 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11383 a_26413_23261# a_25879_22895# a_26318_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11384 a_26183_16911# a_25401_16917# a_26099_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11385 a_3333_9839# _0745_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11386 _0564_.X a_20819_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X11387 vccd1 a_27387_13469# a_27555_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11388 a_9016_29967# a_8767_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11389 a_7256_17429# _0869_.B1 a_7476_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11390 a_20246_8029# a_19973_7663# a_20161_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11391 vssd1 a_19275_21237# a_19233_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11393 a_14805_10357# _0610_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11394 a_14269_19087# a_13735_19093# a_14174_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11395 vssd1 _1033_.CLK a_23303_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11397 a_10613_7119# _0475_.X a_10198_7351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11401 a_8197_21263# a_7663_21269# a_8102_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11402 a_25156_21807# a_24757_21807# a_25030_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11403 a_9301_5487# a_9135_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11404 vssd1 _0756_.A2 a_4989_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X11405 a_6876_21379# _0813_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11406 vccd1 a_4406_3829# a_4333_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11407 a_7469_26703# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11408 a_1757_26703# _0847_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X11409 a_26486_23007# a_26318_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11410 a_25674_14735# a_25235_14741# a_25589_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11411 a_26099_10383# a_25401_10389# a_25842_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11412 a_25708_12015# a_25309_12015# a_25582_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11413 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE a_7111_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11415 vccd1 a_1775_15279# _0812_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11416 a_21836_15279# _0558_.A2 a_21345_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X11417 a_5809_3311# _0566_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11418 vssd1 _0908_.CLK a_4351_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11419 vccd1 a_15963_1653# a_15879_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11420 vccd1 a_25639_8207# a_25807_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11421 vccd1 _0678_.Y _0746_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11422 vssd1 a_11067_19631# _0860_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X11423 a_18887_17024# _1020_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11424 _1019_.CLK a_15667_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11426 vssd1 a_7348_17973# _0742_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X11427 a_9384_32143# a_9135_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11428 a_5245_22057# _0727_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X11429 _0549_.X a_16127_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11430 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11433 _0543_.A1 a_13571_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11434 io_out[1] a_4403_22869# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11435 vccd1 a_9189_18517# _0782_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11438 a_16281_13103# _0917_.D a_16209_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11439 vccd1 _0583_.A a_22015_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11442 a_15812_6005# _0670_.A1 a_16032_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11443 a_2490_25437# a_2051_25071# a_2405_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11444 a_2686_31055# clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11445 a_26781_18909# a_26247_18543# a_26686_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11446 a_5084_16143# _0722_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X11447 a_17980_3311# a_17581_3311# a_17854_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11449 temp1.capload\[15\].cap.B a_2686_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11450 a_13437_2223# _0951_.D a_12999_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11451 vccd1 clkbuf_0__0390_.A a_4802_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11452 a_24420_20553# a_24021_20181# a_24294_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11453 vccd1 a_11435_22895# _0847_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11454 a_8117_18543# _0719_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11455 _1049_.Q a_21667_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11456 a_11782_21085# a_11509_20719# a_11697_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11457 a_11893_20495# _0835_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X11458 _0717_.A2 a_6467_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X11459 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10968_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11461 a_3409_25993# a_2419_25621# a_3283_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11462 a_20855_20175# a_19991_20181# a_20598_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11463 _0565_.B1 _0474_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11465 vccd1 _0964_.CLK a_24591_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11466 _1028_.CLK a_9135_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11467 vssd1 a_13387_4667# a_13345_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11469 a_26225_25993# a_25235_25621# a_26099_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11471 a_2073_30287# _0847_.A2 a_1975_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X11472 _0976_.Q a_28015_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11473 a_10585_14025# a_9595_13653# a_10459_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11474 a_11960_31055# a_11711_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11475 vssd1 _0995_.CLK a_19439_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X11476 a_22822_1501# a_22383_1135# a_22737_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11477 a_21442_24349# a_21169_23983# a_21357_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11478 a_25842_25589# a_25674_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11479 a_15285_1679# _1042_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11481 vssd1 a_13479_2741# a_13437_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11486 vccd1 a_4403_22869# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11487 vccd1 a_3559_4943# a_3727_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11488 a_18371_11293# a_17673_10927# a_18114_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11489 _0880_.Y a_9305_16672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X11490 vccd1 _0959_.CLK a_9779_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11492 a_17539_16161# _0602_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11493 vssd1 a_23415_14459# a_23373_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11495 a_12705_21263# a_12171_21269# a_12610_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11496 a_10677_22729# a_9687_22357# a_10551_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11497 a_22672_3145# a_22273_2773# a_22546_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11498 vssd1 a_18025_7809# _0634_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X11499 a_2858_25615# a_2585_25621# a_2773_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11500 a_12065_8207# _0916_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11503 vssd1 _0827_.A _0821_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11504 a_25674_25615# a_25401_25621# a_25589_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11505 a_25842_21237# a_25674_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11506 clkbuf_1_1__f_net57.A a_1766_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11507 a_4249_19881# _0803_.X _0872_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11508 vssd1 _1076_.Q a_10055_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11511 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15088_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11513 a_22097_6397# _0583_.A a_22015_6144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11514 a_10267_9295# a_9485_9301# a_10183_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11515 vssd1 a_9815_16911# a_9983_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11516 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_13544_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11517 vccd1 a_8123_13647# _0778_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X11518 vssd1 a_10259_7931# a_10217_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11519 a_5325_8181# _0710_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11520 vssd1 a_26267_15797# a_26225_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11521 a_21495_14219# _0842_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11522 vssd1 a_26267_1403# a_26225_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11523 a_5575_4943# a_4793_4949# a_5491_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11524 vssd1 _0793_.X a_6612_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X11525 vccd1 _0745_.A1 a_6682_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X11526 _0798_.A1 a_2686_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11527 a_24719_22351# a_23855_22357# a_24462_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11528 _1017_.D a_23415_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11529 a_12318_8181# a_12150_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11530 vccd1 a_7350_3829# a_7277_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11532 a_22419_22173# a_21555_21807# a_22162_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11534 _0472_.X a_8859_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X11537 vccd1 a_26486_23007# a_26413_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11538 vssd1 _0972_.CLK a_14931_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11539 a_17405_2473# _0551_.C1 a_17323_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11540 a_22449_10499# _0648_.X a_22377_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11541 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_12631_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X11543 a_23891_17999# a_23027_18005# a_23634_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11544 a_10509_18319# _0749_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11545 vccd1 a_5015_1403# a_4931_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11546 a_4333_3855# a_3799_3861# a_4238_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11547 a_10147_15529# _0472_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11548 a_19973_14741# a_19807_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11549 a_23523_4765# a_22659_4399# a_23266_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11550 a_21407_4765# a_20543_4399# a_21150_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11551 a_24389_22351# a_23855_22357# a_24294_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11552 a_15905_25589# _0861_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X11553 a_22089_22173# a_21555_21807# a_21994_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11554 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11556 a_27847_24349# a_26983_23983# a_27590_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11557 vssd1 _0917_.CLK a_11711_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11558 a_6001_11177# _0778_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X11559 vccd1 _0807_.A a_6559_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11560 a_18279_3677# a_17581_3311# a_18022_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11561 vccd1 _1049_.Q a_16902_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X11562 vssd1 a_11582_13077# _0524_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11563 a_4403_22869# _0847_.A3 a_4769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11564 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11566 vssd1 _0658_.X a_22199_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11567 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X11568 a_1674_31599# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11569 a_8151_4765# a_7369_4399# a_8067_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11570 vccd1 clkbuf_1_0__f_io_in[0].X a_1591_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11571 a_23561_17999# a_23027_18005# a_23466_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11572 a_15462_16733# a_15189_16367# a_15377_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11573 _0586_.B2 a_8971_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11574 vccd1 _1015_.CLK a_26707_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11575 a_5812_7439# _0698_.B1 a_5509_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X11576 a_12065_13647# _0917_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11577 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9384_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11578 vssd1 _0964_.CLK a_25051_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11579 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_11746_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11580 vccd1 a_15446_2335# a_15373_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11581 _0600_.X a_15943_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11582 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X11583 a_22741_11177# _0648_.B1 a_22825_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11585 vccd1 a_28015_7931# a_27931_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11586 a_11601_9839# a_11435_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11587 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11588 a_18059_17999# _0584_.A2 a_18237_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X11589 _0959_.D a_10811_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11590 a_8803_1679# a_7939_1685# a_8546_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11591 vssd1 a_12318_13621# a_12276_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11592 a_7472_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11593 vssd1 _0922_.CLK a_9595_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11594 a_24937_3145# a_23947_2773# a_24811_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11595 _0677_.A1 a_6487_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11596 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11597 vccd1 _0999_.CLK a_25235_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11598 _0964_.CLK a_23855_15831# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11599 vccd1 a_12927_3829# a_12843_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11600 a_10142_24847# _0847_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X11601 _0827_.A a_8123_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11602 a_7005_5487# _0545_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11603 vssd1 _0717_.A2 a_6997_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X11605 vccd1 a_17435_22075# a_17351_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11606 vccd1 a_26854_18655# a_26781_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11608 vssd1 _0555_.C1 a_12999_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11609 a_24167_6031# a_23469_6037# a_23910_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11612 vssd1 _1053_.CLK a_9687_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11614 a_22373_12559# _0563_.C1 a_22291_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11615 vssd1 _0836_.Y _0837_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X11616 vssd1 _0483_.X a_24469_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11618 a_14729_23445# a_14563_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11619 _0445_.A _0440_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11620 vssd1 a_25658_17567# a_25616_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11621 a_23190_8207# a_22751_8213# a_23105_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11623 a_14775_15325# a_14483_15279# a_14689_15325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X11624 a_15777_21583# _0863_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11626 vssd1 a_8546_1653# a_8504_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11627 vccd1 _0710_.B2 a_4533_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11628 a_4065_31599# _0814_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11629 vccd1 a_9615_3829# a_9531_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11630 a_6376_7913# _0681_.X a_6635_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X11631 a_16658_26525# a_16219_26159# a_16573_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11635 vssd1 a_24979_2741# a_24937_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11636 a_17415_5737# _0535_.X a_17497_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11637 _0897_.D a_23691_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11638 a_5632_17461# _0456_.A a_5549_17719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11641 _0588_.X a_15023_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X11642 a_27249_10703# _0647_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11643 vccd1 _0842_.A0 a_13735_3968# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11644 vccd1 a_12375_15547# a_12291_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11645 a_25695_1679# _0619_.B1 a_25777_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11646 a_9999_5853# a_9135_5487# a_9742_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11647 _0658_.B1 a_17539_16161# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11648 a_4232_32143# a_3983_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11650 a_18325_9001# _0553_.C1 a_18243_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11651 vssd1 _0860_.A a_16904_24643# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11652 a_14894_9951# a_14726_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11654 vssd1 _0527_.X a_17017_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11655 vccd1 _0959_.CLK a_9411_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11656 vccd1 a_12778_21237# a_12705_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11657 vccd1 _0717_.A2 a_7829_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X11658 a_27422_24349# a_27149_23983# a_27337_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11659 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X11661 a_22948_1135# a_22549_1135# a_22822_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11662 a_17385_19453# _1061_.D a_17313_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11663 a_22879_15823# a_22181_15829# a_22622_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11664 a_8120_14191# _0768_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X11665 a_19329_13647# a_18795_13653# a_19234_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11666 vssd1 _0935_.CLK a_11343_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11667 a_25750_6005# a_25582_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11668 a_15052_9001# _0491_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X11670 a_22454_15823# a_22015_15829# a_22369_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11671 _0549_.C1 a_20267_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X11672 a_15845_12879# _0990_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11673 vssd1 _0995_.CLK a_21831_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11674 vssd1 a_8859_17999# _0472_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11675 a_12249_3855# _0956_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11676 a_4521_1679# _0905_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11678 a_17489_6037# a_17323_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11679 a_6821_6575# _0596_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11680 vssd1 _0616_.B1 a_16548_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X11681 vssd1 _0444_.B _0816_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X11682 a_24945_2223# _1035_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11683 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_9963_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11685 _0847_.A3 a_10055_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11687 a_19605_17455# a_19439_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11688 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11689 vssd1 _0935_.CLK a_12447_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11690 a_22606_15529# _0662_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X11691 a_11980_30511# fanout10.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11692 a_11437_16617# _0882_.A2 _0882_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11694 a_25750_9951# a_25582_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11695 a_10294_22325# a_10126_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11696 vccd1 a_1591_14191# _0456_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11698 a_19195_18337# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11699 vccd1 _0524_.X a_13183_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11700 a_17394_1679# a_17121_1685# a_17309_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11701 _0621_.B2 a_26083_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11702 vccd1 a_16548_10901# _0616_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X11703 vccd1 a_2382_4511# a_2309_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11706 a_17928_8181# _0965_.D a_18148_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11707 a_6997_16143# _0440_.A a_6559_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11708 _0763_.A2 a_7663_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11710 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_12532_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11711 a_17861_1135# _0631_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11712 _0832_.A a_1757_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11713 a_27337_15279# _0893_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11716 a_27973_5487# a_26983_5487# a_27847_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11717 a_25674_19997# a_25235_19631# a_25589_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11719 vccd1 _0813_.A2 a_10567_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X11721 a_17864_13103# _1062_.Q a_17289_13249# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X11722 a_17010_21919# a_16842_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11723 vccd1 _1062_.CLK a_18611_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11724 vssd1 _0533_.X a_17301_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X11725 a_25915_17821# a_25051_17455# a_25658_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11726 a_14641_7663# _1027_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11727 vssd1 _0821_.B a_10239_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11728 vssd1 _0807_.C a_6713_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11729 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_15667_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11731 a_15373_2589# a_14839_2223# a_15278_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11732 a_16895_5281# _0582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11733 a_18141_4399# _0504_.A a_18059_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11734 a_19617_12675# _0580_.X a_19521_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11735 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11738 vssd1 _0959_.CLK a_11895_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11739 vccd1 _0494_.X a_18645_7457# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X11740 _0827_.A a_8123_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11741 _0642_.D_N _0641_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.481 ps=2.78 w=0.65 l=0.15
X11743 a_9494_10927# _0597_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X11744 a_4630_25615# a_4581_25847# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X11746 vccd1 a_23634_17973# a_23561_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11747 _0991_.D a_16055_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11748 _0778_.B1 a_5089_14851# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X11750 vssd1 _1033_.CLK a_24591_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11751 a_20690_21237# a_20522_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11753 vccd1 _1053_.CLK a_14563_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11754 a_10397_15823# _0472_.X a_10147_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11755 vccd1 _0779_.X _0783_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X11756 a_15293_5059# _0553_.X a_15197_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11757 a_2539_9117# a_1757_8751# a_2455_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11758 vssd1 _0842_.A0 _0630_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11759 vccd1 _0845_.C1 a_1591_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11760 vccd1 a_13479_15797# a_13395_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11761 vccd1 a_20414_7775# a_20341_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11763 _0825_.A0 _0825_.A1 a_11251_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11764 _0844_.B a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11765 a_25585_17821# a_25051_17455# a_25490_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11766 a_17654_17567# a_17486_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11767 a_20096_3145# a_19697_2773# a_19970_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11769 a_17765_23261# a_17231_22895# a_17670_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11770 vssd1 _0866_.B a_7283_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11771 vssd1 _0908_.CLK a_8583_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11772 a_2313_1135# _0863_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11773 vssd1 _0483_.X a_22411_6603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11774 vccd1 a_3799_11471# _0861_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11775 a_5066_4943# a_4627_4949# a_4981_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11776 vssd1 _0642_.C a_15671_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11779 vccd1 a_10791_16919# _0935_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11780 a_17470_10357# a_17302_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11781 a_24995_13647# a_24297_13653# a_24738_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11782 a_22622_22325# a_22454_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11783 vccd1 a_12575_8207# a_12743_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11784 _1016_.D a_24703_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11785 a_12604_28879# a_12355_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11786 a_12333_5263# _0673_.A1 a_11987_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X11788 a_22822_19087# a_22383_19093# a_22737_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11789 vccd1 _0527_.X a_16863_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11791 io_out[4] _0752_.Y a_4356_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11792 _0577_.X a_17139_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11793 _0445_.B a_7520_23555# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11794 vccd1 a_20057_16885# _0557_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X11796 a_25539_5853# a_24757_5487# a_25455_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11797 vssd1 a_13309_5515# _0515_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X11798 _0684_.A1 _0652_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11799 vccd1 a_26267_19061# a_26183_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11800 vssd1 a_23047_16885# a_23005_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11801 _1016_.D a_24703_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11802 _0644_.X a_15667_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11803 vssd1 _0845_.A1 a_7244_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11804 a_27422_22173# a_26983_21807# a_27337_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11805 a_19659_1679# a_18795_1685# a_19402_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11806 a_15812_6005# _0669_.X a_16204_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X11807 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE a_11711_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11809 vssd1 a_15503_17973# a_15461_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11810 _0798_.A2 _0722_.C a_4589_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11811 a_14729_16911# _1076_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X11812 a_27931_17821# a_27149_17455# a_27847_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11813 a_11842_25321# _0828_.Y a_11685_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11814 a_23316_8585# a_22917_8213# a_23190_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11815 _0972_.CLK a_15667_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X11816 vssd1 _0518_.Y a_13705_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11817 a_12428_1135# _0850_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X11818 a_25309_12015# a_25143_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11819 temp1.dcdc.Z temp1.dcdc.A a_4232_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11821 vccd1 a_11950_18655# a_11877_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11822 _0440_.A a_2623_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11823 _0680_.Y _0778_.A2 a_7457_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11824 _0644_.A2 a_15975_10721# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11825 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8392_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11826 a_1591_25615# _0840_.X _1078_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11828 _1025_.Q a_20839_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11829 a_17949_3677# a_17415_3311# a_17854_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11831 vssd1 a_24887_20149# a_24845_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11832 a_26870_4765# a_26597_4399# a_26785_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11834 vccd1 a_12242_27791# a_12348_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11836 vccd1 a_4847_2589# a_5015_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11837 a_10218_1679# a_9779_1685# a_10133_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11840 _0460_.C a_1626_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X11841 a_20153_4233# a_19163_3861# a_20027_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11842 a_21213_11809# _0512_.A a_21127_11809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11843 vssd1 a_4590_28447# a_4548_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11844 vssd1 a_19402_1653# a_19360_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11845 _0532_.A2 a_12479_5515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11847 vccd1 _0860_.A a_16986_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X11848 vssd1 a_15595_3829# a_15553_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11849 _0956_.Q a_16607_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11850 vssd1 _1062_.CLK a_25235_19093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11851 a_26628_20719# a_26229_20719# a_26502_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11852 a_12065_6031# _0954_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11858 _0939_.Q a_25623_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11859 _0648_.B1 a_21495_14219# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X11860 a_27847_3677# a_27149_3311# a_27590_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11862 vccd1 _0574_.C a_21127_17249# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X11863 a_20521_7439# _0941_.Q a_20175_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X11864 _0466_.A a_1591_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11865 a_11030_11039# a_10862_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11866 vccd1 a_2991_3579# _0845_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11868 vccd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11869 a_20529_5487# _0669_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11870 vssd1 a_21851_19899# a_21809_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11871 vssd1 a_2962_29967# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11872 vccd1 _0935_.CLK a_11343_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11873 a_2907_1501# a_2125_1135# a_2823_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11874 _0597_.A1_N a_15759_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X11875 _0668_.X a_18059_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X11876 a_22917_8213# a_22751_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11877 _0647_.X a_27167_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X11879 a_6600_27907# _0825_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11880 a_12893_1679# _0604_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11881 a_2686_27791# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11882 a_26233_22895# _0996_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11884 a_26225_16201# a_25235_15829# a_26099_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11885 a_1757_6575# a_1591_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11886 a_2658_28447# a_2490_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11887 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11888 _0556_.D a_12999_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11889 vssd1 a_4811_10383# _0845_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11890 a_4255_12265# _0745_.A1 a_4037_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X11892 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X11893 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11894 a_8123_13647# _0626_.B1 a_8205_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11895 a_5078_30511# temp1.dcdc.Z vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11896 a_7385_27247# _0845_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X11897 a_26536_10927# a_26137_10927# a_26410_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11898 a_13035_12879# _0833_.A a_12935_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X11900 vccd1 _0873_.A a_6553_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X11901 a_11848_25071# _0825_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X11902 a_24619_11471# a_23837_11477# a_24535_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11903 a_21350_18909# a_20911_18543# a_21265_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11905 a_20341_8029# a_19807_7663# a_20246_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11907 _0652_.A a_15671_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X11908 vccd1 _0922_.CLK a_11711_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11909 a_9568_30761# a_9319_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11910 _0847_.X a_1735_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11912 vssd1 a_20393_8545# _0523_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
R32 temp1.capload\[6\].cap_51.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11913 a_27337_14191# _1012_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11914 a_18371_1501# a_17507_1135# a_18114_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11915 vssd1 input2.X a_3523_6039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11917 io_out[5] a_6611_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11918 a_10635_22351# a_9853_22357# a_10551_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11919 a_11987_2473# _0532_.A2 a_12069_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11920 a_5245_22057# _0723_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11921 a_17869_15279# _0937_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11922 vssd1 _0863_.A1 a_14405_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11923 vccd1 a_25658_17567# a_25585_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11924 a_25290_13215# a_25122_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11925 vccd1 a_21575_4667# a_21491_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11926 vssd1 a_3819_26677# a_3777_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11927 vccd1 a_23691_4667# a_23607_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11928 a_18456_7913# _0634_.B1 a_18354_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X11929 vccd1 a_17838_23007# a_17765_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11930 a_19521_10089# _0630_.A2 a_19605_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11931 vccd1 a_12575_11471# a_12743_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11932 a_6713_23805# _0847_.A3 a_6641_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11933 vccd1 a_1959_4951# _0908_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11934 a_12245_7119# _0637_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X11935 vccd1 fanout37.A a_16863_11479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11937 a_16658_26525# a_16385_26159# a_16573_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11938 a_12794_4765# a_12521_4399# a_12709_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11939 a_14012_12925# _0472_.X a_13906_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X11941 vssd1 a_3451_25589# a_3409_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11942 a_19202_15823# _0512_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11944 a_9497_16367# _0880_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11946 a_25589_15823# _0892_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11947 vssd1 a_26099_7119# a_26267_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11948 a_22733_7125# a_22567_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11949 vssd1 a_12575_11471# a_12743_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11950 a_4959_22895# _0742_.A2 a_4769_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11951 a_4847_28701# a_3983_28335# a_4590_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11953 vssd1 a_26267_25589# a_26225_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11955 vssd1 a_7939_19631# _0833_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11956 a_6269_2223# _0910_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11957 vccd1 _0745_.A2 a_4632_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X11958 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_12604_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11959 vssd1 a_10627_13621# a_10585_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11960 a_5091_12021# _0711_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11962 _0707_.A1 _0685_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11963 a_5192_5321# a_4793_4949# a_5066_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11964 vccd1 a_8971_1653# a_8887_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11965 a_16745_6549# _0512_.A a_16998_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X11966 vccd1 a_22622_20149# a_22549_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11967 a_25777_1679# _1072_.D a_25695_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11968 vssd1 a_10719_22325# a_10677_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11969 a_27590_5599# a_27422_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11970 a_9305_16911# _0986_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11971 vccd1 a_27295_4765# a_27463_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11973 vccd1 _0664_.A2 a_26053_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X11974 a_22396_26159# a_21997_26159# a_22270_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11975 a_2655_24501# _0838_.A0 a_2864_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X11976 vccd1 a_2593_15325# a_2693_15543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X11977 vssd1 _0715_.X a_1775_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11978 a_23657_9295# _0894_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11979 a_21625_20719# a_20635_20719# a_21499_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11980 vccd1 a_26099_1501# a_26267_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11981 _0681_.X a_7203_9408# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11984 a_8285_6409# a_7295_6037# a_8159_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11986 a_9673_9295# _0899_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11987 a_3983_15279# _0722_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11988 a_4772_13621# _0791_.A1 a_4995_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X11989 a_6893_25935# _0789_.A2 a_6809_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11990 vssd1 a_2686_23439# _0844_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11991 a_9669_11477# a_9503_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11992 _1000_.Q a_26267_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11993 vccd1 _0583_.A a_20083_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11994 vssd1 a_18079_17723# a_18037_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11995 vssd1 _0964_.CLK a_24591_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11996 vssd1 a_20395_2767# a_20563_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11997 a_1945_6031# _0872_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12001 vccd1 _0964_.CLK a_25235_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12002 a_8123_13647# _0626_.B1 a_8205_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12003 clkbuf_1_0__f_temp1.i_precharge_n.A a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12005 a_21445_2223# a_21279_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12006 a_2833_24759# _0844_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X12007 vssd1 _0527_.X a_16281_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12008 a_10110_21237# a_9942_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12010 a_22097_5487# _1045_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X12011 a_7073_20149# _0798_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X12012 temp1.capload\[1\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12013 vccd1 _0807_.C a_4712_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X12014 _0722_.C a_1867_15831# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X12015 _0899_.Q a_11455_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R33 temp1.capload\[13\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12017 a_10344_2057# a_9945_1685# a_10218_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12018 vccd1 _0572_.A2 a_21361_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X12019 vccd1 a_26099_16911# a_26267_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12021 a_22990_1247# a_22822_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12022 a_27548_23983# a_27149_23983# a_27422_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12023 a_17210_19997# a_16771_19631# a_17125_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12024 a_7939_18543# _0459_.X a_8117_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X12025 a_17302_3855# a_17029_3861# a_17217_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12026 vssd1 _0975_.CLK a_21279_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12027 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12028 a_10533_18776# _1075_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12029 a_10769_5321# a_9779_4949# a_10643_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12030 vssd1 a_27847_10205# a_28015_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12031 a_12815_25071# _0847_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12032 a_4811_27791# _1080_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12033 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X12034 _1048_.D a_26267_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12035 vccd1 _0460_.C a_3983_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12036 a_8293_1679# _0674_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12037 a_17904_14441# _0627_.X a_17802_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X12038 a_13054_2741# a_12886_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12039 a_23569_6825# _1064_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12040 vccd1 a_16182_4511# a_16109_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12041 vccd1 a_7331_6941# a_7499_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12043 a_4422_28701# a_4149_28335# a_4337_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12044 vssd1 a_10567_19061# _0773_.A1_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12046 a_27847_12381# a_27149_12015# a_27590_12127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12048 a_3241_16617# _0872_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X12050 _0518_.Y _0833_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12051 vssd1 a_23174_7093# a_23132_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12052 a_12575_11471# a_11711_11477# a_12318_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12054 a_25405_8751# _1001_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12056 _0813_.A2 a_4132_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12057 a_10133_4943# _0952_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12058 vccd1 a_28015_22075# a_27931_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12059 _0538_.B2 a_7775_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12060 _0511_.D a_9963_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X12061 _0615_.A1 a_20195_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12062 vssd1 a_15170_23413# a_15128_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12063 vssd1 _0583_.C a_16983_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X12064 a_14921_5737# _0542_.X a_14839_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12065 _0656_.Y _0685_.B a_6646_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X12067 _0648_.A2 a_17909_16395# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X12068 a_5060_32143# a_4811_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12069 a_4422_26525# a_3983_26159# a_4337_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12070 vccd1 a_17562_1653# a_17489_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12073 fanout10.A a_11619_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X12074 temp1.capload\[12\].cap.Y temp1.capload\[12\].cap_42.LO a_9865_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12075 a_19536_16143# _0658_.B1 a_19045_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12076 a_11244_27247# _0821_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12077 a_20165_19453# _0583_.A a_20083_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12078 a_12245_11471# a_11711_11477# a_12150_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12080 vssd1 a_25807_8181# a_25765_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12081 vccd1 a_7939_19631# _0833_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12082 vccd1 a_13219_4765# a_13387_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12083 _0618_.C1 a_22015_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X12084 vssd1 _1075_.Q a_15391_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X12085 a_4995_13967# _0791_.A2 a_4901_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X12086 vssd1 clkbuf_1_1__f_net57.A a_1674_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12087 a_21610_24095# a_21442_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12088 a_21675_27613# a_20893_27247# a_21591_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12089 a_18221_22895# a_17231_22895# a_18095_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12090 vccd1 a_19015_4943# a_19183_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12092 vssd1 _0814_.A2 a_2229_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12093 vssd1 _0908_.CLK a_7939_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12094 _0897_.D a_23691_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12095 vccd1 a_26007_10205# a_26175_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12097 vssd1 _1015_.CLK a_26707_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12098 a_14369_13103# _0602_.A a_14287_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12100 vssd1 _0546_.A2 a_8848_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X12101 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12102 _0956_.Q a_16607_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R34 temp1.capload\[5\].cap_50.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12103 a_6815_7913# _0680_.Y a_6376_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X12104 vssd1 a_10110_21237# a_10068_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12105 a_5600_14165# _0768_.A1 a_5820_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12106 vccd1 _0491_.X a_19605_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X12107 vssd1 _0994_.CLK a_25879_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12108 a_20249_21269# a_20083_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12109 a_14921_5737# _0645_.B1 a_15005_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12110 a_10585_15055# _0807_.A a_10147_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12112 vssd1 a_3083_28603# a_3041_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12114 a_25490_9117# a_25051_8751# a_25405_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12115 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12118 a_4582_17705# _0722_.B a_4498_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12120 vccd1 a_1735_29941# _0847_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X12122 vccd1 _0833_.A a_8763_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X12124 _0686_.X a_6653_10933# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X12125 a_10367_21263# a_9669_21269# a_10110_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12126 _0646_.A1 a_6947_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12129 a_7810_4511# a_7642_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12130 a_26099_16911# a_25235_16917# a_25842_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12131 _0515_.B2 a_18355_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12132 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10948_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12133 vccd1 a_21867_13469# a_22035_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12135 a_1766_29423# temp1.inv1_1.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12136 vssd1 fanout27.A a_23487_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12138 a_4863_23413# _0813_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X12139 a_27149_5487# a_26983_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12140 clkbuf_1_1__f_net57.A a_1766_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X12141 a_14737_2767# _0959_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12142 vssd1 a_9411_15279# _0602_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12144 a_23308_18543# _0662_.B1 a_22817_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12145 a_14772_1385# _0670_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.1375 ps=1.275 w=1 l=0.15
X12146 vccd1 a_19827_1653# a_19743_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12147 vssd1 a_21591_27613# a_21759_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12148 clkbuf_1_1__f_net57.X a_1674_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12149 vssd1 _0512_.X a_22637_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X12150 vssd1 a_26083_7931# a_26041_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12152 a_19149_13647# _1025_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12153 vssd1 _0717_.A2 _0717_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X12155 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12156 a_14950_9001# _0599_.X a_14870_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12158 a_9393_7663# a_9227_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12159 vccd1 _1078_.Q a_9503_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X12160 vssd1 a_14453_14557# _0662_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X12161 vssd1 a_19402_13621# a_19360_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12162 a_26042_26525# a_25603_26159# a_25957_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12163 vccd1 _1019_.CLK a_16219_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12164 a_9945_1685# a_9779_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12165 vssd1 a_5491_4943# a_5659_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12166 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12167 vssd1 a_4864_15797# _0795_.A1_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X12169 vccd1 a_11435_22895# _0847_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12170 vssd1 a_1766_30511# temp1.capload\[13\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12173 vccd1 a_13735_12925# _0572_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X12175 _0836_.A a_8031_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12176 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_7288_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12178 vssd1 a_10423_3855# _0959_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12179 a_19605_17455# a_19439_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12180 a_4065_15279# _0722_.A a_3983_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12182 a_1585_24135# _0764_.X a_1863_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12183 a_22369_16911# _1062_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12184 a_3559_4943# a_2861_4949# a_3302_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12188 a_16842_22173# a_16569_21807# a_16757_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12189 vssd1 a_21499_21085# a_21667_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12190 a_6646_18865# _0795_.A2_N a_6645_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X12191 _0992_.D a_21943_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12192 a_13165_2473# _0908_.Q a_13081_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12193 _0849_.X a_12114_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12194 vssd1 a_2198_9269# a_2136_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X12195 vssd1 _0872_.A2 a_3333_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X12197 vccd1 a_10259_7931# a_10175_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12199 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_13367_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12201 a_16439_14557# a_15575_14191# a_16182_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12203 _0515_.B1 a_13309_5515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X12204 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_5060_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12206 vccd1 a_10478_2335# a_10405_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12207 vssd1 _0579_.C a_17385_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12208 a_13054_2741# a_12886_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12209 vssd1 a_27295_4765# a_27463_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12210 a_19149_1679# _0645_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12211 vssd1 a_7683_5755# a_7641_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12212 a_2198_5599# a_2030_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12213 vccd1 a_12318_11445# a_12245_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12214 a_27249_11471# _1068_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12215 _0768_.A2 _0654_.Y a_7663_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12218 vccd1 a_7256_17429# _0719_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X12220 vccd1 _0768_.A2 a_6651_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12222 vssd1 a_25623_22075# a_25581_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12224 a_11782_15645# a_11509_15279# a_11697_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12225 vssd1 _1030_.CLK a_17323_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12227 a_22737_1135# _0967_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12228 a_18225_11471# a_17691_11477# a_18130_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12231 vccd1 _0471_.X a_7226_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12232 a_22948_14191# a_22549_14191# a_22822_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12235 vssd1 a_25163_13621# a_25121_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12236 _0821_.Y _0821_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12237 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X12238 a_3326_2057# a_2762_1801# a_2956_1956# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.06615 ps=0.735 w=0.42 l=0.15
X12239 a_10198_7351# _0566_.B1 a_10335_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12241 _0778_.A2 a_8123_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X12245 a_25156_15279# a_24757_15279# a_25030_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12246 vccd1 a_13311_2767# a_13479_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12247 a_4447_9295# a_4259_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X12248 vssd1 temp1.inv1_1.Y a_1766_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12249 vssd1 a_23247_19087# a_23415_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12251 vssd1 a_17911_17821# a_18079_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12252 vccd1 a_18942_25589# a_18869_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12253 _0951_.D a_11915_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12254 vssd1 _0972_.CLK a_18795_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12255 a_25616_8751# a_25217_8751# a_25490_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12257 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12258 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE a_9871_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12259 vccd1 a_12962_4511# a_12889_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12260 a_21140_10927# _0662_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X12261 vccd1 _0511_.D a_9595_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X12262 a_15837_20719# _0920_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12263 a_20635_1679# _0645_.B1 a_20813_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X12264 a_23189_7663# _1014_.Q a_22751_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12265 a_15483_11177# _0605_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12266 a_2405_12015# a_2228_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X12267 vccd1 a_26007_3677# a_26175_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12268 vssd1 _0502_.X a_20479_8545# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X12269 a_19689_12675# _0576_.X a_19617_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12270 vssd1 a_3099_2767# a_3270_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X12271 a_25750_6005# a_25582_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12272 _0727_.A1 a_7939_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X12273 vccd1 _0972_.CLK a_20543_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12274 a_23193_26709# a_23027_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12275 vssd1 a_12355_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12276 _0863_.Y a_15576_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X12277 a_1674_31599# clkbuf_1_0__f_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12279 vccd1 fanout27.A a_19807_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12280 vssd1 a_11803_23439# _0444_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12281 vccd1 a_23507_20987# a_23423_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12282 vccd1 a_26267_10357# a_26183_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12283 vssd1 a_11765_22325# _0858_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12286 vssd1 a_18095_23261# a_18263_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12287 a_16945_7119# _0672_.C1 a_16863_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12288 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12289 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A a_7472_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12290 vssd1 _1077_.Q a_8859_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X12291 a_24294_22351# a_23855_22357# a_24209_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12292 a_25309_12015# a_25143_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12293 vccd1 _0829_.A1 a_12995_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X12294 vssd1 _0850_.A a_4999_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X12296 a_21508_15279# _0582_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X12298 a_17029_10389# a_16863_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12299 _0612_.X a_19439_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12301 a_26099_21263# a_25401_21269# a_25842_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12302 _0827_.A a_8123_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X12303 vccd1 _0847_.A2 a_9398_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X12304 a_15741_14191# a_15575_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12305 a_13633_6031# _0644_.A2 a_13717_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12306 a_15088_30761# a_14839_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12308 vssd1 _0513_.X a_13521_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12309 vssd1 a_13219_4765# a_13387_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12310 a_4985_12061# _0807_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12313 a_4252_14197# a_4065_14237# a_4165_14455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X12314 a_4974_4765# a_4701_4399# a_4889_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12315 a_15115_5059# _0556_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12316 a_2581_6575# a_1591_6575# a_2455_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12317 vccd1 _0698_.B1 _0695_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12318 vssd1 _0845_.C1 _0837_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12319 a_12805_3311# _0586_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X12320 a_7032_6575# a_6633_6575# a_6906_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12321 a_25589_25615# _0993_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12322 a_25309_6037# a_25143_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12323 vccd1 a_15667_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12324 a_12886_15823# a_12613_15829# a_12801_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12325 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12326 _0866_.Y _0845_.A1 a_7565_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12327 a_15607_15307# _0521_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12328 a_9613_25045# _0816_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X12330 vccd1 clkbuf_1_0__f_io_in[0].X a_1959_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12332 a_25765_12937# a_24775_12565# a_25639_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12333 vssd1 _0768_.A1 a_6704_13077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X12334 vccd1 _1048_.D a_22974_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X12335 a_22641_20719# a_22475_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12336 a_25842_19061# a_25674_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12337 a_22637_12015# _0939_.Q a_22199_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12338 vccd1 temp1.capload\[11\].cap_41.LO temp1.capload\[11\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12340 temp1.capload\[10\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12341 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].vref.TE a_18059_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12342 _0934_.Q a_17435_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12343 a_21108_3311# a_20709_3311# a_20982_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12345 a_4356_23983# _0814_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X12346 _0819_.S _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X12347 a_7648_17705# _0717_.B1 a_7393_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X12348 _0551_.C1 a_20911_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X12349 a_6608_29111# _0825_.A1 a_6750_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X12350 a_10405_2589# a_9871_2223# a_10310_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12351 a_12713_7913# _0646_.C1 a_12631_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12352 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12353 vccd1 _0999_.CLK a_23855_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12355 a_20175_7119# _0516_.B1 a_20257_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12357 vccd1 a_17470_3829# a_17397_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12358 vssd1 _0491_.X a_17761_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X12359 a_27931_2589# a_27149_2223# a_27847_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12360 vccd1 _1030_.CLK a_17507_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12363 vssd1 a_2991_3579# _0845_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12364 _0675_.D a_11527_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X12365 a_25674_19087# a_25401_19093# a_25589_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12366 a_16182_14303# a_16014_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12367 a_26444_22895# a_26045_22895# a_26318_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12368 vccd1 fanout24.A a_16035_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X12369 _0751_.B1 a_10331_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X12370 vccd1 clkbuf_1_0__f_io_in[0].X a_2235_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12372 a_14373_31599# temp1.capload\[13\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12373 _0479_.Y _1079_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12374 a_2658_28447# a_2490_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12377 vccd1 a_23082_20831# a_23009_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12378 a_25971_13647# _0648_.B1 a_26053_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X12379 vssd1 a_2915_28701# a_3083_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12380 a_4981_4943# _0677_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12381 vccd1 a_18298_11445# a_18225_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12383 _0990_.D a_12375_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12386 _0601_.B1 a_14655_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12387 vssd1 _1019_.CLK a_16403_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12388 vccd1 _1076_.Q a_13091_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12389 vccd1 a_2686_15823# _0444_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12390 vssd1 a_16863_11479# fanout27.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12391 a_22369_1679# _0618_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12393 a_23082_20831# a_22914_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12394 a_24167_6031# a_23303_6037# a_23910_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12395 vccd1 a_1766_30511# temp1.capload\[13\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R35 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12397 vccd1 _1028_.CLK a_11711_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12398 vccd1 a_24811_2767# a_24979_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12399 vccd1 a_6612_14709# _0795_.A2_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X12400 a_24757_4399# a_24591_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12402 a_19015_20175# a_18151_20181# a_18758_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12403 a_11697_18543# _0918_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12404 a_23013_8751# _0488_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12405 a_16209_10089# _0676_.B _0679_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12406 a_18114_11039# a_17946_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12408 a_17305_19997# a_16771_19631# a_17210_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12409 _0882_.Y _0882_.A2 a_11437_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12410 vssd1 a_10018_4511# a_9976_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12411 vssd1 a_27590_17567# a_27548_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12412 _0456_.B a_1591_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X12413 a_6001_11177# _0807_.B _0708_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12415 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_5547_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12416 a_15821_16189# _1055_.Q a_15749_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12419 a_23247_1501# a_22383_1135# a_22990_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12421 _0839_.B a_2655_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12422 _0910_.Q a_3727_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12423 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_15667_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12424 _0497_.A1 a_15595_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12425 a_5894_3677# a_5455_3311# a_5809_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12426 vccd1 _0504_.A a_20543_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12427 vccd1 fanout27.A a_16863_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12428 a_10212_29967# a_9963_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12429 a_18685_20175# a_18151_20181# a_18590_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12430 a_22974_18793# _0662_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X12431 vccd1 _0648_.A2 a_19697_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X12434 _0827_.A a_8123_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X12435 a_18187_6031# a_17489_6037# a_17930_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12436 vssd1 _0666_.X _0679_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12437 vccd1 a_18703_12567# _0504_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12438 vccd1 _0816_.S a_6498_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12440 a_1945_5487# _0880_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12441 a_15151_12381# a_14453_12015# a_14894_12127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12443 vssd1 a_25658_8863# a_25616_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12444 _0573_.B a_26267_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12445 _0657_.X a_6416_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12447 _1081_.Q a_5015_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12448 _0837_.Y _0837_.A1 a_7385_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12450 vccd1 a_5399_4765# a_5567_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12451 vssd1 _0814_.A2 a_6713_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12452 a_25658_17567# a_25490_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12454 a_15170_3829# a_15002_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12455 a_20257_7439# _0649_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X12456 a_25674_19087# a_25235_19093# a_25589_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12458 a_15197_13103# _0471_.X a_15115_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X12459 a_2133_15101# _0722_.A a_2051_14848# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12462 a_5727_7119# _0656_.Y a_5509_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X12463 vssd1 a_10091_8029# a_10259_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12464 vccd1 _1067_.D a_24068_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X12465 vssd1 a_5047_21781# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12467 _0835_.A1 a_2626_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X12468 vssd1 a_4221_8725# _0699_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12469 a_7623_10901# _0699_.A0 a_7832_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X12470 _0441_.B a_5015_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12471 a_24021_22357# a_23855_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12472 vccd1 _1033_.CLK a_22751_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12473 a_24212_12879# _1067_.D a_23637_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X12475 a_19439_12675# _0584_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X12476 a_11789_9839# _0625_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12478 vccd1 a_19439_14191# _1062_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12479 a_11413_10927# a_10423_10927# a_11287_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12481 a_22449_15253# _0512_.A a_22702_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X12482 vssd1 a_7074_6687# a_7032_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12483 a_4035_13077# _0791_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X12484 a_15538_27765# a_15370_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12485 a_11509_18543# a_11343_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12486 _0464_.X a_2051_14848# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12487 a_24757_5487# a_24591_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12488 a_23303_10383# _0558_.A2 a_23385_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12489 _0444_.Y _0444_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12491 _1025_.Q a_20839_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12493 a_15170_23413# a_15002_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12494 vccd1 fanout37.A a_9227_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X12495 vccd1 a_10551_22351# a_10719_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12496 a_13311_2767# a_12447_2773# a_13054_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12497 a_17501_2223# _0969_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X12499 vssd1 _0441_.B a_11435_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X12500 a_4589_17999# _0722_.B a_4167_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12501 a_27847_17821# a_26983_17455# a_27590_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12502 vccd1 _0521_.A a_19439_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12504 _0583_.C a_14603_18589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X12505 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8944_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12506 a_9899_16911# a_9117_16917# a_9815_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12507 a_15370_27791# a_15097_27797# a_15285_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12509 vssd1 a_21150_3423# a_21108_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12510 vccd1 clkbuf_1_0__f_io_in[0].X a_1959_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12511 _1062_.Q a_21023_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12513 a_22641_20719# a_22475_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12514 a_7369_4399# a_7203_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12515 _0935_.Q a_13203_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12516 _0628_.X a_15667_15936# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12517 _0671_.B2 a_20195_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12519 vccd1 _0667_.B1 a_16685_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12521 vccd1 a_20671_14735# a_20839_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12523 _1062_.Q a_21023_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12524 vssd1 _0565_.B1 a_15812_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X12525 a_4864_11445# _0708_.B1 a_4993_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X12527 _0935_.Q a_13203_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12528 vccd1 a_15135_20149# a_15051_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12529 a_15170_3829# a_15002_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12530 vccd1 _0444_.A a_2051_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12532 vccd1 fanout27.A a_20819_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12533 vssd1 a_13054_2741# a_13012_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12534 vssd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12535 a_10788_25615# _0847_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12536 a_26812_18543# a_26413_18543# a_26686_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12537 a_10202_13621# a_10034_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12538 _1029_.Q a_18539_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12539 vssd1 _0574_.C a_17811_15073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X12540 a_25731_6941# a_25033_6575# a_25474_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12541 a_2198_6687# a_2030_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12542 _0825_.S _0840_.A1 a_11798_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X12543 a_9326_25071# _0816_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X12544 a_24895_2767# a_24113_2773# a_24811_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12545 vssd1 _0668_.X a_15391_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X12546 _0702_.B1_N a_4852_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12547 vccd1 _0840_.A1 a_11711_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X12548 vccd1 a_17378_19743# a_17305_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12550 vccd1 a_18758_4917# a_18685_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12551 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_8116_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12552 a_2686_27791# clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X12553 a_26053_13647# _1012_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12554 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12555 vssd1 _0893_.CLK a_24683_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12556 vccd1 _0444_.A a_3983_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12557 vccd1 _1031_.Q a_18456_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X12558 vccd1 _1019_.CLK a_16403_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12560 a_22917_19087# a_22383_19093# a_22822_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12561 _0798_.A2 _0722_.C a_4589_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12563 vssd1 _0662_.B1 a_25489_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X12564 a_10034_13647# a_9761_13653# a_9949_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12566 vccd1 _1053_.D a_18282_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X12568 _1045_.D a_19827_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12569 vssd1 _0935_.CLK a_14103_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12570 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_9496_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12571 vccd1 a_2686_31055# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12572 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10212_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12573 vccd1 a_18758_20149# a_18685_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12574 temp1.capload\[3\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12575 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE a_14195_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12576 _0880_.A1 a_8155_16161# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X12578 clkbuf_1_1__f__0390_.A a_4802_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12580 vccd1 a_5813_25117# a_5913_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X12581 a_20556_22729# a_20157_22357# a_20430_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12582 a_20237_19453# _1019_.D a_20165_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12583 a_27195_18909# a_26413_18543# a_27111_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12585 a_24941_12565# a_24775_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12586 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE a_14839_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12587 vccd1 _1062_.CLK a_23855_15831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X12588 vccd1 a_10719_6005# a_10635_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12591 a_6020_3311# a_5621_3311# a_5894_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12592 a_11237_3311# _0543_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12593 a_14809_4399# _0954_.Q a_14737_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12595 vccd1 _0847_.A2 a_6958_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12596 _0965_.D a_24059_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12597 a_27422_17821# a_27149_17455# a_27337_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12599 clkbuf_1_1__f__0390_.A a_4802_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12600 vccd1 _0833_.A a_10814_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12601 _1066_.D a_28015_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12602 a_23910_9269# a_23742_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12603 a_24945_15279# _0891_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12604 a_11815_12265# _0474_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12605 _0710_.A2 _0680_.Y a_6645_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12606 vssd1 a_25639_8207# a_25807_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12607 a_8037_14441# _0768_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12609 a_4248_29673# _0845_.B1 a_3993_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12611 vssd1 _0975_.CLK a_22659_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12613 _0659_.X a_22199_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X12614 a_2455_5853# a_1591_5487# a_2198_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12615 a_15427_23439# a_14729_23445# a_15170_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12616 a_27422_15645# a_26983_15279# a_27337_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12617 vssd1 _1080_.Q a_11936_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12618 vssd1 _0466_.A a_9781_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12621 a_27422_3677# a_26983_3311# a_27337_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12623 vssd1 _0880_.A2 a_9497_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X12624 a_13119_21263# a_12337_21269# a_13035_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12626 a_4882_19087# a_4705_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12627 a_20797_7663# a_19807_7663# a_20671_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12628 a_2915_25437# a_2217_25071# a_2658_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12629 a_21583_21085# a_20801_20719# a_21499_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12630 vssd1 a_24462_20149# a_24420_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12631 a_8105_4949# a_7939_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12632 a_26133_9839# a_25143_9839# a_26007_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12634 a_12886_2767# a_12447_2773# a_12801_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12636 vssd1 _1019_.CLK a_16219_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12637 a_17302_10383# a_17029_10389# a_17217_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12638 a_17017_15101# _0919_.D a_16945_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12641 a_14894_12127# a_14726_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12642 vccd1 a_9644_26311# _0820_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X12643 a_14261_7235# _0544_.B a_14189_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12644 vccd1 a_23358_8181# a_23285_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12645 _0564_.D a_22291_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X12646 a_9583_13103# _0768_.A1 _0747_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X12647 a_15370_27791# a_14931_27797# a_15285_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12649 a_4901_13967# _0791_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X12652 a_18850_21237# a_18682_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12654 a_18427_2473# _0591_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12655 vssd1 a_26083_17723# a_26041_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12656 _0663_.X a_23579_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X12657 a_8546_4917# a_8378_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12658 vccd1 _0872_.A1 a_3424_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X12659 vccd1 _0471_.X a_10397_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X12662 _0656_.Y _0655_.X a_6559_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12663 a_6809_25935# _0787_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12665 vssd1 _0684_.A1 a_7663_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12666 a_17657_13621# _0606_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X12667 vssd1 a_26099_16911# a_26267_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12668 _0877_.Y a_4429_16672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X12669 _0517_.B a_19439_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X12670 a_19439_9001# _0517_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12671 a_24661_11849# a_23671_11477# a_24535_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12672 vccd1 _0824_.Y a_12355_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12673 a_19347_8207# _0515_.B1 a_19429_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X12675 a_2861_4949# a_2695_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12677 vccd1 a_15427_3855# a_15595_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12678 vccd1 a_22015_3855# _0975_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12679 _0614_.X a_15483_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X12680 a_18045_11471# _0897_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12681 vccd1 a_15667_2767# _0972_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12682 vssd1 a_5399_4765# a_5567_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12684 a_21993_23983# a_21003_23983# a_21867_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12685 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12686 temp1.capload\[15\].cap.B a_2686_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12687 a_15759_1385# _0645_.B1 a_15841_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12688 a_18685_4943# a_18151_4949# a_18590_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12689 vssd1 a_11287_11293# a_11455_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12691 a_26229_20719# a_26063_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12692 vccd1 a_4802_27247# clkbuf_1_1__f__0390_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12693 a_16937_19631# a_16771_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12694 vssd1 a_20761_9633# _0506_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X12695 a_4606_1679# a_4333_1685# a_4521_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12696 vccd1 a_11913_13336# a_11582_13077# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X12697 a_10126_22351# a_9853_22357# a_10041_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12698 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12700 a_17029_2773# a_16863_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12701 a_22659_11471# _0662_.B1 a_22741_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X12702 a_4137_15279# _0722_.B a_4065_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12703 vssd1 a_18022_3423# a_17980_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12706 _0873_.Y _0873_.A a_3057_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12707 a_19973_7663# a_19807_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12708 vssd1 a_17470_10357# a_17428_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12709 vccd1 a_10107_10615# _0626_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X12710 vssd1 _0582_.C a_17937_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12711 _0613_.A1 a_10351_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12712 vccd1 _0444_.A a_1959_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12714 _0613_.C1 a_13183_7232# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12715 vssd1 _0699_.A0 a_4253_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X12716 vssd1 _0847_.A2 a_12815_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12717 vccd1 a_26099_19997# a_26267_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12718 vccd1 _1080_.Q a_4811_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12719 a_17995_16395# _0842_.A0 a_17909_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12720 a_27698_4943# a_27521_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12721 a_25490_8029# a_25217_7663# a_25405_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12722 a_15017_5487# _0543_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X12723 _0843_.Y _0845_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12724 vssd1 _0584_.C1 a_19773_18689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X12726 a_2780_3145# a_2401_2773# a_2683_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X12727 vccd1 a_24335_6005# a_24251_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12728 a_20022_18793# _0583_.X a_19773_18689# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X12729 a_25581_9615# _1066_.D a_25143_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12730 _0866_.B a_13367_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X12731 vccd1 a_4132_17429# _0813_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12733 a_9834_7775# a_9666_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12734 a_19202_15823# _1060_.D a_19045_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12735 a_5100_4399# a_4701_4399# a_4974_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12736 _0548_.A1 a_26175_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12737 vssd1 _0505_.A2 a_17761_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X12738 vccd1 a_2686_28879# _0845_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12740 vssd1 a_12375_20987# a_12333_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12741 _0710_.B2 a_5128_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12742 a_10110_11445# a_9942_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12743 a_13311_15823# a_12613_15829# a_13054_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12744 a_1674_32143# clkbuf_1_1__f_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12746 _0999_.Q a_28015_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12747 vccd1 _0935_.CLK a_8951_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12748 a_9834_7775# a_9666_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12749 a_26137_10927# a_25971_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12750 vssd1 a_22863_26427# a_22821_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12751 _0850_.A a_3270_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X12752 vccd1 a_23415_1403# a_23331_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12753 a_25957_26159# _0994_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12754 vssd1 _0797_.A1 a_13080_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X12755 _0951_.D a_11915_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12756 clkbuf_1_1__f_net57.X a_1674_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X12757 vssd1 a_25807_12533# a_25765_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12758 a_27931_10205# a_27149_9839# a_27847_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12760 a_20111_3855# a_19329_3861# a_20027_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12761 a_12575_11471# a_11877_11477# a_12318_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12763 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE a_6191_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12764 vccd1 a_28015_16635# a_27931_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12765 vssd1 a_11915_3579# a_11873_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12767 a_2229_23983# _0444_.B a_2113_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X12768 a_2842_2741# a_2683_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12769 vccd1 fanout11.A a_11619_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X12770 a_27337_25071# _0998_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12772 vssd1 a_5509_7093# _0695_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12773 a_6815_7913# _0656_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12774 vssd1 a_4663_3855# a_4831_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12775 _0844_.B a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12776 a_12291_18909# a_11509_18543# a_12207_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12777 a_24386_2767# a_23947_2773# a_24301_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12778 a_6833_13103# _0745_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X12780 a_18900_25993# a_18501_25621# a_18774_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12781 a_14188_30287# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12782 vccd1 _1080_.Q a_12018_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12783 vssd1 _0999_.CLK a_26983_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12784 a_23285_8207# a_22751_8213# a_23190_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12786 a_13771_22351# a_12907_22357# a_13514_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12787 vssd1 a_10564_20407# _0774_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X12788 _1023_.Q a_23047_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12790 a_4498_17705# _0722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12791 a_27548_3311# a_27149_3311# a_27422_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12793 a_16354_18543# _1053_.Q a_16264_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X12794 a_19981_1385# _0976_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12795 a_1766_29423# temp1.inv1_1.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X12796 a_22015_5737# _0645_.B1 a_22097_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12797 a_16986_24643# _0860_.B a_16904_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12799 a_27422_14557# a_26983_14191# a_27337_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12801 _1023_.Q a_23047_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12802 vssd1 a_4882_19087# a_4988_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12803 a_13012_3145# a_12613_2773# a_12886_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12804 a_25405_8751# _1001_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12805 vccd1 a_4771_12791# _0734_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X12806 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_11527_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12807 vccd1 _0845_.C1 a_5547_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12809 a_6916_22671# _0866_.Y a_6613_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X12810 temp1.dcdc.A a_1674_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12812 vssd1 a_20635_13655# _0583_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12813 a_25842_10357# a_25674_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12814 a_13441_22351# a_12907_22357# a_13346_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12818 a_20214_16911# _0582_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X12819 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12820 a_11885_14735# _0880_.A1 _0882_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12821 a_15427_3855# a_14563_3861# a_15170_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12824 a_25581_4399# a_24591_4399# a_25455_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12825 vssd1 a_13514_10357# a_13472_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12826 _0505_.X a_22659_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X12827 a_12428_1135# _0835_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12829 a_2686_10383# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12830 _0970_.Q a_17895_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12831 vssd1 _1030_.CLK a_17507_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12832 vssd1 a_27923_9019# a_27881_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12833 vssd1 fanout10.A a_10147_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12834 a_5157_2057# a_4167_1685# a_5031_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12835 vccd1 a_24167_9295# a_24335_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12836 a_24167_9295# a_23469_9301# a_23910_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12837 _0602_.A a_9411_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X12838 a_25248_13103# a_24849_13103# a_25122_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12841 _1030_.CLK a_16035_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X12842 _0642_.C a_12079_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X12843 a_25674_10383# a_25401_10389# a_25589_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12844 a_16853_9001# _0615_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12845 clkbuf_1_0__f_io_in[0].X a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X12846 a_26099_3855# a_25235_3861# a_25842_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12847 _0986_.D a_10535_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12848 vssd1 _1033_.CLK a_25143_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12849 a_23523_9117# a_22825_8751# a_23266_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12851 a_2639_4765# a_1941_4399# a_2382_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12853 vssd1 _1028_.CLK a_14287_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12854 a_5047_21781# _0726_.X a_5245_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X12855 _0836_.A a_8031_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X12856 a_13771_10383# a_13073_10389# a_13514_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12857 a_27981_4943# a_27804_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X12858 a_23005_17289# a_22015_16917# a_22879_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12859 vssd1 a_15170_3829# a_15128_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12861 a_27149_25071# a_26983_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12862 a_17497_5737# _0622_.B2 a_17415_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12865 a_26877_13103# _1066_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12866 a_27149_23983# a_26983_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12867 a_22580_22729# a_22181_22357# a_22454_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12869 a_4248_29673# _0845_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12870 a_2773_25615# _1078_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12871 a_27847_8029# a_27149_7663# a_27590_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12872 a_6813_19087# _0869_.B1 a_6559_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12873 vssd1 _0464_.X a_3523_13655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12874 a_5547_25615# _0839_.B _0839_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12875 a_12723_3561# _0532_.A2 a_12805_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12877 a_10359_4765# a_9577_4399# a_10275_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12878 _0471_.X a_9503_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12879 a_14453_9839# a_14287_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12880 a_18179_23261# a_17397_22895# a_18095_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12881 a_10703_19407# _0761_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X12883 vssd1 a_18611_14735# _0662_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12884 a_26229_20719# a_26063_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12885 a_24021_1685# a_23855_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12887 a_23833_6575# _1064_.Q a_23487_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X12888 vssd1 _0579_.C a_17625_16161# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X12889 a_22741_11471# _0505_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12891 vssd1 _0758_.B1 a_6336_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X12892 a_7090_5853# a_6651_5487# a_7005_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12893 a_19329_26709# a_19163_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12894 a_21502_15529# _0662_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X12895 a_19689_9269# _0512_.A a_19942_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X12896 a_20977_10901# _0643_.B1 a_21134_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12897 vssd1 a_8175_11989# _0655_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12898 vccd1 fanout10.A a_10791_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12899 vccd1 a_16553_15425# _0580_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X12904 vccd1 a_10643_4943# a_10811_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12906 vssd1 a_25842_10357# a_25800_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12907 vssd1 a_23415_3579# a_23373_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12908 vssd1 a_2686_28879# _0845_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12910 a_19208_16143# _0582_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X12911 a_6354_2589# a_5915_2223# a_6269_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12912 a_13544_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12914 vccd1 a_1766_29423# clkbuf_1_1__f_net57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12915 vssd1 a_19773_18689# _0584_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X12916 a_20709_3311# a_20543_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12917 vccd1 _1030_.CLK a_18151_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12918 vssd1 _0572_.A2 a_23936_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X12919 a_16097_14013# _1050_.Q a_16025_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12920 a_22373_16617# _1067_.Q a_22291_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12921 a_9997_12061# a_9595_12015# a_9911_12061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X12922 vccd1 _0972_.CLK a_16955_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12924 vccd1 a_2686_27791# _0798_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12926 _0999_.CLK a_22659_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X12930 _0623_.D a_17415_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X12931 a_25842_15797# a_25674_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12932 a_25658_17567# a_25490_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12933 a_5989_3677# a_5455_3311# a_5894_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12934 a_6663_8751# _0746_.A2 a_6556_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X12935 a_26137_10927# a_25971_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12936 vssd1 _0577_.C a_15821_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12937 a_16553_15425# _0579_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X12941 _0523_.X a_17691_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X12942 vssd1 _1030_.CLK a_20543_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12943 a_17838_23007# a_17670_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12944 a_25674_10383# a_25235_10389# a_25589_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12945 vssd1 a_25915_17821# a_26083_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12946 a_11067_14191# _0747_.B1 a_11245_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X12947 vssd1 _0489_.C1 a_19531_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12948 vssd1 a_1674_32143# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12949 vccd1 a_1674_31599# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X12950 a_25455_2589# a_24757_2223# a_25198_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12951 temp1.capload\[13\].cap.B a_1766_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12952 a_24512_3145# a_24113_2773# a_24386_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12953 a_8193_4399# a_7203_4399# a_8067_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12954 a_10727_4943# a_9945_4949# a_10643_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12955 vssd1 a_12575_8207# a_12743_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12956 a_13544_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12957 a_26689_13103# a_26523_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12958 vccd1 a_10535_21237# a_10451_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12959 a_7745_15529# _0760_.B1 a_7829_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12960 a_15002_23439# a_14563_23445# a_14917_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12961 vccd1 _0577_.C a_11929_9633# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X12962 vccd1 _0460_.C a_1867_15831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X12963 a_15005_2223# a_14839_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12964 vccd1 a_2623_5755# a_2539_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12966 a_15002_3855# a_14563_3861# a_14917_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12967 a_6863_2589# a_6081_2223# a_6779_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12968 vccd1 _0487_.X a_15105_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X12971 _0441_.B a_5015_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12972 vssd1 a_27590_3423# a_27548_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12973 temp1.capload\[13\].cap.B a_1766_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12974 _0952_.Q a_14307_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12975 vccd1 a_13514_22325# a_13441_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12976 vccd1 a_20027_6031# a_20195_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12977 a_19429_8207# _0515_.B2 a_19347_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12978 vccd1 _0647_.X a_22449_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X12979 vccd1 a_7623_10901# _0776_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X12980 vccd1 fanout10.A a_9871_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12981 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A a_15016_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12982 vccd1 _0999_.CLK a_26983_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12983 vccd1 a_10533_18776# a_10202_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X12984 vccd1 a_10167_1403# a_10083_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12985 vssd1 _0995_.CLK a_23027_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12986 _0761_.B a_5642_19637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X12987 vccd1 a_9190_3829# a_9117_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12988 _0831_.B clkbuf_1_0__f_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12989 vccd1 a_21867_24349# a_22035_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12990 a_9758_9295# a_9485_9301# a_9673_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12991 _0440_.A a_2623_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12993 _0633_.X a_20543_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12994 vccd1 _0860_.B a_15575_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12995 vccd1 a_2823_3677# a_2991_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12996 vccd1 a_2198_9269# a_2132_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X12998 _0825_.S _0444_.B a_11711_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12999 a_18409_21269# a_18243_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13000 _0669_.X a_21279_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13001 _1019_.D a_20195_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13002 a_1674_26159# clkbuf_1_1__f_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13003 _0861_.A2 a_16904_24643# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13004 vssd1 clkbuf_1_0__f_io_in[0].X a_1959_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13005 _0695_.A1 _0656_.Y a_5621_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X13006 a_13303_4765# a_12521_4399# a_13219_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13007 _0645_.B1 a_15793_6603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X13008 vssd1 _0515_.B1 a_12333_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X13009 vccd1 _0763_.A2 a_8305_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X13010 a_4167_17999# _0722_.B a_4589_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13012 clkbuf_1_0__f_net57.X a_1674_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X13013 a_20204_18793# _0584_.B1 a_20102_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X13014 a_12659_8207# a_11877_8213# a_12575_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13015 vssd1 _0686_.A a_6653_10933# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X13016 vssd1 _0658_.B1 a_17864_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X13017 vccd1 a_19402_13621# a_19329_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13018 vssd1 fanout27.A a_15575_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13019 vssd1 a_10535_11445# a_10493_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13020 a_22281_12265# _0563_.B1 a_22365_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13021 vccd1 _0511_.D a_15115_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X13022 a_14621_8897# _0601_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13023 vssd1 a_26175_10107# a_26133_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13024 _0928_.D a_28015_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13025 vssd1 a_9184_25223# _0817_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X13026 a_22829_20719# _0963_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13034 a_5443_29967# _0827_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X13035 vssd1 a_17895_3829# a_17853_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13036 vccd1 a_27847_12381# a_28015_12283# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13038 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A _0819_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13039 a_12809_7663# _0924_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X13040 vccd1 _0717_.A2 a_7393_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13041 a_13311_2767# a_12613_2773# a_13054_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13042 vssd1 a_2686_10383# clkbuf_1_0__f_io_in[0].X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13043 a_18497_10927# a_17507_10927# a_18371_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13044 a_22737_19087# _1016_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13045 _0838_.A0 _0472_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13046 a_21361_6575# _0669_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X13048 a_15749_12559# _0667_.B1 a_15833_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13049 vccd1 a_24059_26677# a_23975_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13050 vssd1 _0999_.CLK a_22475_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13051 _0587_.C1 a_12723_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X13052 a_10876_21813# a_10689_21853# a_10789_22071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X13053 vssd1 a_25623_15547# a_25581_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13054 vssd1 _0444_.A a_3983_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13055 vssd1 _0722_.A a_4170_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X13056 vccd1 a_4774_1653# a_4701_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13057 _0515_.X a_19347_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X13059 vccd1 a_5549_17719# _0797_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13060 a_27847_16733# a_27149_16367# a_27590_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13061 a_15235_8029# a_14453_7663# a_15151_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13063 a_4863_23413# _0813_.A2 a_5081_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X13064 vccd1 a_10198_7351# _0567_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X13066 a_22917_3677# a_22383_3311# a_22822_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13067 _0924_.D a_12743_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13068 a_21767_9117# a_20985_8751# a_21683_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13069 a_25198_4511# a_25030_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13071 _0440_.C a_5547_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X13072 a_7216_5487# a_6817_5487# a_7090_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13073 vccd1 _0824_.Y a_13183_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13074 a_14710_20149# a_14542_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13075 _0577_.C a_10202_18517# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X13076 a_14559_15823# _0797_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13077 _0924_.D a_12743_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13078 _1027_.Q a_13847_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13079 vccd1 _0831_.D a_10055_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X13081 a_3327_16367# _0873_.A _0877_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X13083 a_11983_22351# _0861_.B1 a_11765_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X13085 a_6480_2223# a_6081_2223# a_6354_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13086 a_12886_15823# a_12447_15829# a_12801_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13087 a_22549_14191# a_22383_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13088 a_14542_20175# a_14269_20181# a_14457_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13089 vccd1 _0807_.C a_6559_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13090 a_7192_27497# _0836_.Y a_6937_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13092 _0798_.A1 a_2686_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13096 vssd1 a_2686_15823# _0444_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X13097 _0770_.B2 _0461_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13098 a_7801_11079# _0438_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X13101 _0506_.A2 a_20761_9633# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X13102 vccd1 _1047_.D a_22606_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X13103 _1061_.Q a_19367_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13104 a_14559_15823# _0798_.A2 a_14341_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X13106 vccd1 a_28015_3579# a_27931_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13108 vssd1 a_20839_7931# a_20797_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13109 a_19329_6037# a_19163_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13111 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z a_10048_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13112 a_25401_15829# a_25235_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13114 vssd1 a_10735_2589# a_10903_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13115 vssd1 _0917_.CLK a_12907_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13116 _1061_.Q a_19367_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13118 vssd1 _0735_.A2 a_7928_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X13119 vccd1 a_21039_5853# a_21207_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13120 a_12333_15279# a_11343_15279# a_12207_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13121 vssd1 _1033_.CLK a_25235_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13122 a_7734_6031# a_7461_6037# a_7649_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13126 a_20801_1679# _0946_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X13127 a_24949_18319# _0993_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X13129 a_4590_28447# a_4422_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13131 vssd1 _0561_.C1 a_19531_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13132 vccd1 _0893_.CLK a_26983_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13133 vccd1 a_14729_16911# _0582_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X13134 a_19689_9001# _0517_.B a_19617_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13135 vccd1 a_5692_13077# _0714_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X13136 a_23661_14735# _0662_.X a_23579_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13137 vssd1 _0972_.CLK a_17415_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13138 a_22833_7913# _0506_.A2 a_22917_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13139 a_6376_7913# _0680_.Y a_6815_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X13140 vssd1 a_4847_28701# a_5015_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13141 a_15916_29967# a_15667_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X13142 vccd1 a_26267_21237# a_26183_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13143 a_11371_11293# a_10589_10927# a_11287_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13144 vssd1 a_26911_23163# a_26869_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13145 vccd1 _0445_.A a_7843_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X13146 _0622_.A1 a_18539_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13147 vccd1 _0644_.A2 a_14829_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13148 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A a_15023_28887# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X13149 a_12777_24501# _0444_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X13150 a_12245_7119# _0899_.Q a_12161_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13151 a_18053_10089# a_17865_9845# a_17971_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X13152 a_2915_25437# a_2051_25071# a_2658_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13153 vssd1 _0461_.A a_6467_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13154 vccd1 _0845_.A2 a_4984_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13155 _0850_.Y _0850_.A a_12815_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
D6 vssd1 _0880_.Y sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X13156 _0845_.B1 _0844_.B a_4811_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13158 vssd1 _0776_.A2 a_4468_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X13159 a_16929_17973# _0662_.A1 a_17182_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X13161 a_16439_4765# a_15741_4399# a_16182_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13162 a_15759_9001# _0587_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13163 a_24673_11177# _0562_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X13164 vssd1 a_14805_10357# _0614_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X13165 a_15922_21085# a_15483_20719# a_15837_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13166 _0474_.X a_10147_15529# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X13168 io_out[0] a_5047_21781# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13169 vccd1 a_15595_3829# a_15511_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13170 a_13817_4221# _0842_.A0 a_13735_3968# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13171 a_23013_8751# _0488_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13173 a_2585_25437# a_2051_25071# a_2490_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13174 a_13717_6031# _1027_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X13176 a_11693_6825# _0674_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X13177 a_21683_19997# a_20819_19631# a_21426_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13178 _1062_.CLK a_19439_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13179 a_20801_1679# _1041_.Q a_20717_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13180 a_4701_1679# a_4167_1685# a_4606_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13181 a_22622_16885# a_22454_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13182 _0553_.C1 a_23487_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X13183 a_17158_12265# _0557_.X a_17078_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13184 a_14967_20175# a_14269_20181# a_14710_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13185 a_18187_6031# a_17323_6037# a_17930_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13186 _0624_.C a_22751_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X13187 vccd1 a_26267_3829# a_26183_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13188 a_25765_23817# a_24775_23445# a_25639_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13189 vssd1 _0444_.A a_1959_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13190 _0723_.X a_6416_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13191 a_19602_3855# a_19329_3861# a_19517_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13192 vccd1 a_12318_6005# a_12245_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13193 _0840_.A1 a_2991_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13194 vssd1 _0836_.A _0529_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13195 vssd1 _0866_.B a_6437_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13196 a_21353_19997# a_20819_19631# a_21258_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13197 a_4517_26525# a_3983_26159# a_4422_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13198 _0749_.B1 a_11067_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X13199 a_24719_20175# a_24021_20181# a_24462_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13200 a_7607_3855# a_6743_3861# a_7350_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13201 a_7037_29177# _0825_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X13202 a_23757_15055# _0963_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X13203 vccd1 _0999_.CLK a_22475_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13204 _0566_.B1 a_15115_5059# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X13205 a_26045_22895# a_25879_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13206 vccd1 _0491_.X a_12069_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13207 a_19283_25615# a_18501_25621# a_19199_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13208 a_11333_5737# _0907_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X13209 vccd1 _0652_.A a_15115_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13210 a_14805_10357# _0612_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X13211 vccd1 _0837_.A1 a_7192_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13212 vccd1 a_27038_4511# a_26965_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13213 a_8661_7119# _0653_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13214 vssd1 a_2566_27359# a_2524_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13215 a_5329_21807# _0809_.B2 a_5245_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X13216 a_7461_6037# a_7295_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13217 _0843_.B a_4035_25045# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13218 vccd1 _0583_.A a_23303_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13219 a_15611_3677# a_14747_3311# a_15354_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13220 vssd1 a_7258_5599# a_7216_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13221 vccd1 _0847_.A3 a_11711_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X13222 _0694_.A2 _0689_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13223 vssd1 _0758_.A1 _0758_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13224 vccd1 _0506_.A2 a_19981_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13226 a_16863_14848# _0919_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13227 vssd1 a_15538_27765# a_15496_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13229 a_17121_1685# a_16955_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13232 a_5547_17027# _0807_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X13234 vssd1 a_7350_3829# a_7308_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13237 a_16882_15529# _0580_.C1 a_16802_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X13238 vccd1 a_22879_1679# a_23047_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13240 a_25030_16733# a_24591_16367# a_24945_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13241 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13242 a_16127_7663# _0644_.A2 a_16305_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
C0 a_25589_1135# vssd1 0.23fF $ **FLOATING
C1 a_26099_1501# vssd1 0.61fF $ **FLOATING
C2 a_26267_1403# vssd1 0.82fF $ **FLOATING
C3 a_25674_1501# vssd1 0.63fF $ **FLOATING
C4 a_25842_1247# vssd1 0.58fF $ **FLOATING
C5 a_25401_1135# vssd1 1.43fF $ **FLOATING
C6 a_25235_1135# vssd1 1.81fF $ **FLOATING
C7 a_22737_1135# vssd1 0.23fF $ **FLOATING
C8 a_23247_1501# vssd1 0.61fF $ **FLOATING
C9 a_23415_1403# vssd1 0.82fF $ **FLOATING
C10 a_22822_1501# vssd1 0.63fF $ **FLOATING
C11 a_22990_1247# vssd1 0.58fF $ **FLOATING
C12 a_22549_1135# vssd1 1.43fF $ **FLOATING
C13 a_22383_1135# vssd1 1.81fF $ **FLOATING
C14 a_20993_1385# vssd1 0.21fF $ **FLOATING
C15 a_19981_1385# vssd1 0.21fF $ **FLOATING
C16 a_12428_1135# vssd1 0.34fF $ **FLOATING
C17 a_11895_1135# vssd1 0.28fF $ **FLOATING
C18 a_17861_1135# vssd1 0.23fF $ **FLOATING
C19 a_20911_1385# vssd1 0.80fF $ **FLOATING
C20 a_19899_1385# vssd1 0.80fF $ **FLOATING
C21 a_18371_1501# vssd1 0.61fF $ **FLOATING
C22 a_18539_1403# vssd1 0.82fF $ **FLOATING
C23 a_17946_1501# vssd1 0.63fF $ **FLOATING
C24 a_18114_1247# vssd1 0.58fF $ **FLOATING
C25 a_17673_1135# vssd1 1.43fF $ **FLOATING
C26 a_17507_1135# vssd1 1.81fF $ **FLOATING
C27 a_15841_1385# vssd1 0.21fF $ **FLOATING
C28 a_14772_1385# vssd1 0.24fF $ **FLOATING
C29 a_12342_1385# vssd1 0.32fF $ **FLOATING
C30 a_9489_1135# vssd1 0.23fF $ **FLOATING
C31 a_15759_1385# vssd1 0.80fF $ **FLOATING
C32 a_11895_1385# vssd1 1.14fF $ **FLOATING
C33 a_9999_1501# vssd1 0.61fF $ **FLOATING
C34 a_10167_1403# vssd1 0.82fF $ **FLOATING
C35 a_9574_1501# vssd1 0.63fF $ **FLOATING
C36 a_9742_1247# vssd1 0.58fF $ **FLOATING
C37 a_9301_1135# vssd1 1.43fF $ **FLOATING
C38 a_9135_1135# vssd1 1.81fF $ **FLOATING
C39 a_4337_1135# vssd1 0.23fF $ **FLOATING
C40 a_4847_1501# vssd1 0.61fF $ **FLOATING
C41 a_5015_1403# vssd1 0.82fF $ **FLOATING
C42 a_4422_1501# vssd1 0.63fF $ **FLOATING
C43 a_4590_1247# vssd1 0.58fF $ **FLOATING
C44 a_4149_1135# vssd1 1.43fF $ **FLOATING
C45 a_3983_1135# vssd1 1.81fF $ **FLOATING
C46 a_2313_1135# vssd1 0.23fF $ **FLOATING
C47 a_2823_1501# vssd1 0.61fF $ **FLOATING
C48 a_2991_1403# vssd1 0.97fF $ **FLOATING
C49 a_2398_1501# vssd1 0.63fF $ **FLOATING
C50 a_2566_1247# vssd1 0.58fF $ **FLOATING
C51 a_2125_1135# vssd1 1.43fF $ **FLOATING
C52 a_1959_1135# vssd1 1.81fF $ **FLOATING
C53 a_25777_1679# vssd1 0.21fF $ **FLOATING
C54 a_24209_1679# vssd1 0.23fF $ **FLOATING
C55 a_20801_1679# vssd1 0.21fF $ **FLOATING
C56 a_20717_1679# vssd1 0.17fF $ **FLOATING
C57 a_22369_1679# vssd1 0.23fF $ **FLOATING
C58 a_19149_1679# vssd1 0.23fF $ **FLOATING
C59 a_17309_1679# vssd1 0.23fF $ **FLOATING
C60 a_15285_1679# vssd1 0.23fF $ **FLOATING
C61 a_12893_1679# vssd1 0.23fF $ **FLOATING
C62 _0641_.D1 vssd1 1.87fF $ **FLOATING
C63 a_10133_1679# vssd1 0.23fF $ **FLOATING
C64 a_8293_1679# vssd1 0.23fF $ **FLOATING
C65 a_4521_1679# vssd1 0.23fF $ **FLOATING
C66 a_3326_2057# vssd1 0.22fF $ **FLOATING
C67 a_25695_1679# vssd1 0.80fF $ **FLOATING
C68 a_24719_1679# vssd1 0.61fF $ **FLOATING
C69 a_24887_1653# vssd1 0.82fF $ **FLOATING
C70 a_24294_1679# vssd1 0.63fF $ **FLOATING
C71 a_24462_1653# vssd1 0.58fF $ **FLOATING
C72 a_24021_1685# vssd1 1.43fF $ **FLOATING
C73 a_23855_1685# vssd1 1.81fF $ **FLOATING
C74 a_22879_1679# vssd1 0.61fF $ **FLOATING
C75 a_23047_1653# vssd1 0.82fF $ **FLOATING
C76 a_22454_1679# vssd1 0.63fF $ **FLOATING
C77 a_22622_1653# vssd1 0.58fF $ **FLOATING
C78 a_22181_1685# vssd1 1.43fF $ **FLOATING
C79 a_22015_1685# vssd1 1.81fF $ **FLOATING
C80 a_20635_1679# vssd1 0.97fF $ **FLOATING
C81 _0660_.X vssd1 2.99fF $ **FLOATING
C82 a_19659_1679# vssd1 0.61fF $ **FLOATING
C83 a_19827_1653# vssd1 0.82fF $ **FLOATING
C84 a_19234_1679# vssd1 0.63fF $ **FLOATING
C85 a_19402_1653# vssd1 0.58fF $ **FLOATING
C86 a_18961_1685# vssd1 1.43fF $ **FLOATING
C87 a_18795_1685# vssd1 1.81fF $ **FLOATING
C88 a_17819_1679# vssd1 0.61fF $ **FLOATING
C89 a_17987_1653# vssd1 0.82fF $ **FLOATING
C90 a_17394_1679# vssd1 0.63fF $ **FLOATING
C91 a_17562_1653# vssd1 0.58fF $ **FLOATING
C92 a_17121_1685# vssd1 1.43fF $ **FLOATING
C93 a_16955_1685# vssd1 1.81fF $ **FLOATING
C94 a_15795_1679# vssd1 0.61fF $ **FLOATING
C95 a_15963_1653# vssd1 0.82fF $ **FLOATING
C96 a_15370_1679# vssd1 0.63fF $ **FLOATING
C97 a_15538_1653# vssd1 0.58fF $ **FLOATING
C98 a_15097_1685# vssd1 1.43fF $ **FLOATING
C99 a_14931_1685# vssd1 1.81fF $ **FLOATING
C100 a_13403_1679# vssd1 0.61fF $ **FLOATING
C101 a_13571_1653# vssd1 0.82fF $ **FLOATING
C102 a_12978_1679# vssd1 0.63fF $ **FLOATING
C103 a_13146_1653# vssd1 0.58fF $ **FLOATING
C104 a_12705_1685# vssd1 1.43fF $ **FLOATING
C105 a_12539_1685# vssd1 1.81fF $ **FLOATING
C106 a_11711_1792# vssd1 0.62fF $ **FLOATING
C107 a_10643_1679# vssd1 0.61fF $ **FLOATING
C108 a_10811_1653# vssd1 0.82fF $ **FLOATING
C109 a_10218_1679# vssd1 0.63fF $ **FLOATING
C110 a_10386_1653# vssd1 0.58fF $ **FLOATING
C111 a_9945_1685# vssd1 1.43fF $ **FLOATING
C112 a_9779_1685# vssd1 1.81fF $ **FLOATING
C113 a_8803_1679# vssd1 0.61fF $ **FLOATING
C114 a_8971_1653# vssd1 0.82fF $ **FLOATING
C115 a_8378_1679# vssd1 0.63fF $ **FLOATING
C116 a_8546_1653# vssd1 0.58fF $ **FLOATING
C117 a_8105_1685# vssd1 1.43fF $ **FLOATING
C118 a_7939_1685# vssd1 1.81fF $ **FLOATING
C119 a_5031_1679# vssd1 0.61fF $ **FLOATING
C120 a_5199_1653# vssd1 0.82fF $ **FLOATING
C121 a_4606_1679# vssd1 0.63fF $ **FLOATING
C122 a_4774_1653# vssd1 0.58fF $ **FLOATING
C123 a_4333_1685# vssd1 1.43fF $ **FLOATING
C124 a_4167_1685# vssd1 1.81fF $ **FLOATING
C125 a_2885_2057# vssd1 0.59fF $ **FLOATING
C126 a_2956_1956# vssd1 0.63fF $ **FLOATING
C127 a_2762_1801# vssd1 1.39fF $ **FLOATING
C128 a_2752_1897# vssd1 1.77fF $ **FLOATING
C129 a_2464_1653# vssd1 0.60fF $ **FLOATING
C130 a_2114_1653# vssd1 1.41fF $ **FLOATING
C131 _0976_.Q vssd1 5.65fF $ **FLOATING
C132 a_27337_2223# vssd1 0.23fF $ **FLOATING
C133 a_27847_2589# vssd1 0.61fF $ **FLOATING
C134 a_28015_2491# vssd1 0.82fF $ **FLOATING
C135 a_27422_2589# vssd1 0.63fF $ **FLOATING
C136 a_27590_2335# vssd1 0.58fF $ **FLOATING
C137 a_27149_2223# vssd1 1.43fF $ **FLOATING
C138 a_26983_2223# vssd1 1.81fF $ **FLOATING
C139 a_24945_2223# vssd1 0.23fF $ **FLOATING
C140 a_25455_2589# vssd1 0.61fF $ **FLOATING
C141 a_25623_2491# vssd1 0.82fF $ **FLOATING
C142 a_25030_2589# vssd1 0.63fF $ **FLOATING
C143 a_25198_2335# vssd1 0.58fF $ **FLOATING
C144 a_24757_2223# vssd1 1.43fF $ **FLOATING
C145 a_24591_2223# vssd1 1.81fF $ **FLOATING
C146 a_21633_2223# vssd1 0.23fF $ **FLOATING
C147 a_22143_2589# vssd1 0.61fF $ **FLOATING
C148 a_22311_2491# vssd1 0.82fF $ **FLOATING
C149 a_21718_2589# vssd1 0.63fF $ **FLOATING
C150 a_21886_2335# vssd1 0.58fF $ **FLOATING
C151 a_21445_2223# vssd1 1.43fF $ **FLOATING
C152 a_21279_2223# vssd1 1.81fF $ **FLOATING
C153 _0594_.C vssd1 2.16fF $ **FLOATING
C154 _0594_.D vssd1 2.01fF $ **FLOATING
C155 a_17489_2473# vssd1 0.21fF $ **FLOATING
C156 a_17405_2473# vssd1 0.17fF $ **FLOATING
C157 a_15193_2223# vssd1 0.23fF $ **FLOATING
C158 a_18427_2473# vssd1 0.70fF $ **FLOATING
C159 a_17323_2223# vssd1 0.97fF $ **FLOATING
C160 _0551_.C1 vssd1 3.20fF $ **FLOATING
C161 a_15703_2589# vssd1 0.61fF $ **FLOATING
C162 a_15871_2491# vssd1 0.82fF $ **FLOATING
C163 a_15278_2589# vssd1 0.63fF $ **FLOATING
C164 a_15446_2335# vssd1 0.58fF $ **FLOATING
C165 a_15005_2223# vssd1 1.43fF $ **FLOATING
C166 a_14839_2223# vssd1 1.81fF $ **FLOATING
C167 a_13165_2473# vssd1 0.21fF $ **FLOATING
C168 a_13081_2473# vssd1 0.17fF $ **FLOATING
C169 a_12069_2473# vssd1 0.21fF $ **FLOATING
C170 a_10225_2223# vssd1 0.23fF $ **FLOATING
C171 a_12999_2223# vssd1 0.97fF $ **FLOATING
C172 _0555_.C1 vssd1 0.78fF $ **FLOATING
C173 a_11987_2473# vssd1 0.80fF $ **FLOATING
C174 _0945_.D vssd1 3.79fF $ **FLOATING
C175 a_10735_2589# vssd1 0.61fF $ **FLOATING
C176 a_10903_2491# vssd1 0.82fF $ **FLOATING
C177 a_10310_2589# vssd1 0.63fF $ **FLOATING
C178 a_10478_2335# vssd1 0.58fF $ **FLOATING
C179 a_10037_2223# vssd1 1.43fF $ **FLOATING
C180 a_9871_2223# vssd1 1.81fF $ **FLOATING
C181 a_6269_2223# vssd1 0.23fF $ **FLOATING
C182 a_6779_2589# vssd1 0.61fF $ **FLOATING
C183 a_6947_2491# vssd1 0.82fF $ **FLOATING
C184 a_6354_2589# vssd1 0.63fF $ **FLOATING
C185 a_6522_2335# vssd1 0.58fF $ **FLOATING
C186 a_6081_2223# vssd1 1.43fF $ **FLOATING
C187 a_5915_2223# vssd1 1.81fF $ **FLOATING
C188 a_4337_2223# vssd1 0.23fF $ **FLOATING
C189 a_4847_2589# vssd1 0.61fF $ **FLOATING
C190 a_5015_2491# vssd1 0.97fF $ **FLOATING
C191 a_4422_2589# vssd1 0.63fF $ **FLOATING
C192 a_4590_2335# vssd1 0.58fF $ **FLOATING
C193 a_4149_2223# vssd1 1.43fF $ **FLOATING
C194 a_3983_2223# vssd1 1.81fF $ **FLOATING
C195 a_2313_2223# vssd1 0.23fF $ **FLOATING
C196 a_2823_2589# vssd1 0.61fF $ **FLOATING
C197 a_2991_2491# vssd1 0.97fF $ **FLOATING
C198 a_2398_2589# vssd1 0.63fF $ **FLOATING
C199 a_2566_2335# vssd1 0.58fF $ **FLOATING
C200 a_2125_2223# vssd1 1.43fF $ **FLOATING
C201 a_1959_2223# vssd1 1.81fF $ **FLOATING
C202 _1035_.Q vssd1 2.16fF $ **FLOATING
C203 a_24301_2767# vssd1 0.23fF $ **FLOATING
C204 a_22461_2767# vssd1 0.23fF $ **FLOATING
C205 a_19885_2767# vssd1 0.23fF $ **FLOATING
C206 a_14737_2767# vssd1 0.21fF $ **FLOATING
C207 a_17217_2767# vssd1 0.23fF $ **FLOATING
C208 _0591_.X vssd1 2.31fF $ **FLOATING
C209 a_12801_2767# vssd1 0.23fF $ **FLOATING
C210 a_10133_2767# vssd1 0.23fF $ **FLOATING
C211 _0905_.Q vssd1 5.14fF $ **FLOATING
C212 a_4705_2767# vssd1 0.23fF $ **FLOATING
C213 a_2589_2767# vssd1 0.22fF $ **FLOATING
C214 a_24811_2767# vssd1 0.61fF $ **FLOATING
C215 a_24979_2741# vssd1 0.82fF $ **FLOATING
C216 a_24386_2767# vssd1 0.63fF $ **FLOATING
C217 a_24554_2741# vssd1 0.58fF $ **FLOATING
C218 a_24113_2773# vssd1 1.43fF $ **FLOATING
C219 a_23947_2773# vssd1 1.81fF $ **FLOATING
C220 a_22971_2767# vssd1 0.61fF $ **FLOATING
C221 a_23139_2741# vssd1 0.82fF $ **FLOATING
C222 a_22546_2767# vssd1 0.63fF $ **FLOATING
C223 a_22714_2741# vssd1 0.58fF $ **FLOATING
C224 a_22273_2773# vssd1 1.43fF $ **FLOATING
C225 a_22107_2773# vssd1 1.81fF $ **FLOATING
C226 a_20395_2767# vssd1 0.61fF $ **FLOATING
C227 a_20563_2741# vssd1 0.82fF $ **FLOATING
C228 a_19970_2767# vssd1 0.63fF $ **FLOATING
C229 a_20138_2741# vssd1 0.58fF $ **FLOATING
C230 a_19697_2773# vssd1 1.43fF $ **FLOATING
C231 a_19531_2773# vssd1 1.81fF $ **FLOATING
C232 a_17727_2767# vssd1 0.61fF $ **FLOATING
C233 a_17895_2741# vssd1 0.82fF $ **FLOATING
C234 a_17302_2767# vssd1 0.63fF $ **FLOATING
C235 a_17470_2741# vssd1 0.58fF $ **FLOATING
C236 a_17029_2773# vssd1 1.43fF $ **FLOATING
C237 a_16863_2773# vssd1 1.81fF $ **FLOATING
C238 a_15667_2767# vssd1 0.70fF $ **FLOATING
C239 a_14655_2767# vssd1 0.80fF $ **FLOATING
C240 a_13311_2767# vssd1 0.61fF $ **FLOATING
C241 a_13479_2741# vssd1 0.82fF $ **FLOATING
C242 a_12886_2767# vssd1 0.63fF $ **FLOATING
C243 a_13054_2741# vssd1 0.58fF $ **FLOATING
C244 a_12613_2773# vssd1 1.43fF $ **FLOATING
C245 a_12447_2773# vssd1 1.81fF $ **FLOATING
C246 a_10643_2767# vssd1 0.61fF $ **FLOATING
C247 a_10811_2741# vssd1 0.82fF $ **FLOATING
C248 a_10218_2767# vssd1 0.63fF $ **FLOATING
C249 a_10386_2741# vssd1 0.58fF $ **FLOATING
C250 a_9945_2773# vssd1 1.43fF $ **FLOATING
C251 a_9779_2773# vssd1 1.81fF $ **FLOATING
C252 a_5215_2767# vssd1 0.61fF $ **FLOATING
C253 a_5383_2741# vssd1 0.82fF $ **FLOATING
C254 a_4790_2767# vssd1 0.63fF $ **FLOATING
C255 a_4958_2741# vssd1 0.58fF $ **FLOATING
C256 a_4517_2773# vssd1 1.43fF $ **FLOATING
C257 a_4351_2773# vssd1 1.81fF $ **FLOATING
C258 a_3099_2767# vssd1 0.60fF $ **FLOATING
C259 a_3270_2741# vssd1 1.41fF $ **FLOATING
C260 a_2683_2767# vssd1 0.63fF $ **FLOATING
C261 a_2842_2741# vssd1 0.59fF $ **FLOATING
C262 a_2401_2773# vssd1 1.39fF $ **FLOATING
C263 a_2235_2773# vssd1 1.77fF $ **FLOATING
C264 a_27337_3311# vssd1 0.23fF $ **FLOATING
C265 a_27847_3677# vssd1 0.61fF $ **FLOATING
C266 a_28015_3579# vssd1 0.82fF $ **FLOATING
C267 a_27422_3677# vssd1 0.63fF $ **FLOATING
C268 a_27590_3423# vssd1 0.58fF $ **FLOATING
C269 a_27149_3311# vssd1 1.43fF $ **FLOATING
C270 a_26983_3311# vssd1 1.81fF $ **FLOATING
C271 _1034_.Q vssd1 4.30fF $ **FLOATING
C272 a_25497_3311# vssd1 0.23fF $ **FLOATING
C273 a_26007_3677# vssd1 0.61fF $ **FLOATING
C274 a_26175_3579# vssd1 0.82fF $ **FLOATING
C275 a_25582_3677# vssd1 0.63fF $ **FLOATING
C276 a_25750_3423# vssd1 0.58fF $ **FLOATING
C277 a_25309_3311# vssd1 1.43fF $ **FLOATING
C278 a_25143_3311# vssd1 1.81fF $ **FLOATING
C279 a_22737_3311# vssd1 0.23fF $ **FLOATING
C280 a_23247_3677# vssd1 0.61fF $ **FLOATING
C281 a_23415_3579# vssd1 0.82fF $ **FLOATING
C282 a_22822_3677# vssd1 0.63fF $ **FLOATING
C283 a_22990_3423# vssd1 0.58fF $ **FLOATING
C284 a_22549_3311# vssd1 1.43fF $ **FLOATING
C285 a_22383_3311# vssd1 1.81fF $ **FLOATING
C286 a_20897_3311# vssd1 0.23fF $ **FLOATING
C287 a_21407_3677# vssd1 0.61fF $ **FLOATING
C288 a_21575_3579# vssd1 0.82fF $ **FLOATING
C289 a_20982_3677# vssd1 0.63fF $ **FLOATING
C290 a_21150_3423# vssd1 0.58fF $ **FLOATING
C291 a_20709_3311# vssd1 1.43fF $ **FLOATING
C292 a_20543_3311# vssd1 1.81fF $ **FLOATING
C293 _1042_.Q vssd1 3.50fF $ **FLOATING
C294 a_17769_3311# vssd1 0.23fF $ **FLOATING
C295 a_18279_3677# vssd1 0.61fF $ **FLOATING
C296 a_18447_3579# vssd1 0.82fF $ **FLOATING
C297 a_17854_3677# vssd1 0.63fF $ **FLOATING
C298 a_18022_3423# vssd1 0.58fF $ **FLOATING
C299 a_17581_3311# vssd1 1.43fF $ **FLOATING
C300 _1041_.Q vssd1 3.66fF $ **FLOATING
C301 a_17415_3311# vssd1 1.81fF $ **FLOATING
C302 _0946_.Q vssd1 3.57fF $ **FLOATING
C303 a_15101_3311# vssd1 0.23fF $ **FLOATING
C304 a_15611_3677# vssd1 0.61fF $ **FLOATING
C305 a_15779_3579# vssd1 0.82fF $ **FLOATING
C306 a_15186_3677# vssd1 0.63fF $ **FLOATING
C307 a_15354_3423# vssd1 0.58fF $ **FLOATING
C308 a_14913_3311# vssd1 1.43fF $ **FLOATING
C309 _0946_.D vssd1 4.33fF $ **FLOATING
C310 a_14747_3311# vssd1 1.81fF $ **FLOATING
C311 a_12805_3561# vssd1 0.21fF $ **FLOATING
C312 a_11237_3311# vssd1 0.23fF $ **FLOATING
C313 a_12723_3561# vssd1 0.80fF $ **FLOATING
C314 _0586_.B2 vssd1 5.12fF $ **FLOATING
C315 a_11747_3677# vssd1 0.61fF $ **FLOATING
C316 a_11915_3579# vssd1 0.82fF $ **FLOATING
C317 a_11322_3677# vssd1 0.63fF $ **FLOATING
C318 a_11490_3423# vssd1 0.58fF $ **FLOATING
C319 a_11049_3311# vssd1 1.43fF $ **FLOATING
C320 a_10883_3311# vssd1 1.81fF $ **FLOATING
C321 a_5809_3311# vssd1 0.23fF $ **FLOATING
C322 a_6319_3677# vssd1 0.61fF $ **FLOATING
C323 a_6487_3579# vssd1 0.82fF $ **FLOATING
C324 a_5894_3677# vssd1 0.63fF $ **FLOATING
C325 a_6062_3423# vssd1 0.58fF $ **FLOATING
C326 a_5621_3311# vssd1 1.43fF $ **FLOATING
C327 a_5455_3311# vssd1 1.81fF $ **FLOATING
C328 a_2313_3311# vssd1 0.23fF $ **FLOATING
C329 a_3983_3311# vssd1 0.70fF $ **FLOATING
C330 io_in[1] vssd1 2.32fF
C331 a_2823_3677# vssd1 0.61fF $ **FLOATING
C332 a_2991_3579# vssd1 0.97fF $ **FLOATING
C333 a_2398_3677# vssd1 0.63fF $ **FLOATING
C334 a_2566_3423# vssd1 0.58fF $ **FLOATING
C335 a_2125_3311# vssd1 1.43fF $ **FLOATING
C336 a_1959_3311# vssd1 1.81fF $ **FLOATING
C337 a_25589_3855# vssd1 0.23fF $ **FLOATING
C338 a_19517_3855# vssd1 0.23fF $ **FLOATING
C339 _0970_.Q vssd1 2.94fF $ **FLOATING
C340 a_17217_3855# vssd1 0.23fF $ **FLOATING
C341 a_14917_3855# vssd1 0.23fF $ **FLOATING
C342 _0639_.X vssd1 1.92fF $ **FLOATING
C343 a_12249_3855# vssd1 0.23fF $ **FLOATING
C344 a_8937_3855# vssd1 0.23fF $ **FLOATING
C345 a_7097_3855# vssd1 0.23fF $ **FLOATING
C346 a_4153_3855# vssd1 0.23fF $ **FLOATING
C347 a_2037_3855# vssd1 0.23fF $ **FLOATING
C348 a_26099_3855# vssd1 0.61fF $ **FLOATING
C349 a_26267_3829# vssd1 0.82fF $ **FLOATING
C350 a_25674_3855# vssd1 0.63fF $ **FLOATING
C351 a_25842_3829# vssd1 0.58fF $ **FLOATING
C352 a_25401_3861# vssd1 1.43fF $ **FLOATING
C353 _1072_.D vssd1 2.78fF $ **FLOATING
C354 a_25235_3861# vssd1 1.81fF $ **FLOATING
C355 a_22015_3855# vssd1 0.70fF $ **FLOATING
C356 a_20027_3855# vssd1 0.61fF $ **FLOATING
C357 a_20195_3829# vssd1 0.82fF $ **FLOATING
C358 a_19602_3855# vssd1 0.63fF $ **FLOATING
C359 a_19770_3829# vssd1 0.58fF $ **FLOATING
C360 a_19329_3861# vssd1 1.43fF $ **FLOATING
C361 _0969_.D vssd1 5.65fF $ **FLOATING
C362 a_19163_3861# vssd1 1.81fF $ **FLOATING
C363 a_17727_3855# vssd1 0.61fF $ **FLOATING
C364 a_17895_3829# vssd1 0.82fF $ **FLOATING
C365 a_17302_3855# vssd1 0.63fF $ **FLOATING
C366 a_17470_3829# vssd1 0.58fF $ **FLOATING
C367 a_17029_3861# vssd1 1.43fF $ **FLOATING
C368 a_16863_3861# vssd1 1.81fF $ **FLOATING
C369 a_15427_3855# vssd1 0.61fF $ **FLOATING
C370 a_15595_3829# vssd1 0.82fF $ **FLOATING
C371 a_15002_3855# vssd1 0.63fF $ **FLOATING
C372 a_15170_3829# vssd1 0.58fF $ **FLOATING
C373 a_14729_3861# vssd1 1.43fF $ **FLOATING
C374 a_14563_3861# vssd1 1.81fF $ **FLOATING
C375 a_13735_3968# vssd1 0.62fF $ **FLOATING
C376 _0639_.B vssd1 3.74fF $ **FLOATING
C377 a_12759_3855# vssd1 0.61fF $ **FLOATING
C378 a_12927_3829# vssd1 0.82fF $ **FLOATING
C379 a_12334_3855# vssd1 0.63fF $ **FLOATING
C380 a_12502_3829# vssd1 0.58fF $ **FLOATING
C381 a_12061_3861# vssd1 1.43fF $ **FLOATING
C382 a_11895_3861# vssd1 1.81fF $ **FLOATING
C383 a_10423_3855# vssd1 0.70fF $ **FLOATING
C384 a_9447_3855# vssd1 0.61fF $ **FLOATING
C385 a_9615_3829# vssd1 0.82fF $ **FLOATING
C386 a_9022_3855# vssd1 0.63fF $ **FLOATING
C387 a_9190_3829# vssd1 0.58fF $ **FLOATING
C388 a_8749_3861# vssd1 1.43fF $ **FLOATING
C389 a_8583_3861# vssd1 1.81fF $ **FLOATING
C390 a_7607_3855# vssd1 0.61fF $ **FLOATING
C391 a_7775_3829# vssd1 0.82fF $ **FLOATING
C392 a_7182_3855# vssd1 0.63fF $ **FLOATING
C393 a_7350_3829# vssd1 0.58fF $ **FLOATING
C394 a_6909_3861# vssd1 1.43fF $ **FLOATING
C395 a_6743_3861# vssd1 1.81fF $ **FLOATING
C396 a_4663_3855# vssd1 0.61fF $ **FLOATING
C397 a_4831_3829# vssd1 0.82fF $ **FLOATING
C398 a_4238_3855# vssd1 0.63fF $ **FLOATING
C399 a_4406_3829# vssd1 0.58fF $ **FLOATING
C400 a_3965_3861# vssd1 1.43fF $ **FLOATING
C401 a_3799_3861# vssd1 1.81fF $ **FLOATING
C402 a_2547_3855# vssd1 0.61fF $ **FLOATING
C403 a_2715_3829# vssd1 0.82fF $ **FLOATING
C404 a_2122_3855# vssd1 0.63fF $ **FLOATING
C405 a_2290_3829# vssd1 0.58fF $ **FLOATING
C406 a_1849_3861# vssd1 1.43fF $ **FLOATING
C407 a_1683_3861# vssd1 1.81fF $ **FLOATING
C408 a_26785_4399# vssd1 0.23fF $ **FLOATING
C409 a_27295_4765# vssd1 0.61fF $ **FLOATING
C410 a_27463_4667# vssd1 0.82fF $ **FLOATING
C411 a_26870_4765# vssd1 0.63fF $ **FLOATING
C412 a_27038_4511# vssd1 0.58fF $ **FLOATING
C413 a_26597_4399# vssd1 1.43fF $ **FLOATING
C414 a_26431_4399# vssd1 1.81fF $ **FLOATING
C415 a_24945_4399# vssd1 0.23fF $ **FLOATING
C416 a_25455_4765# vssd1 0.61fF $ **FLOATING
C417 a_25623_4667# vssd1 0.82fF $ **FLOATING
C418 a_25030_4765# vssd1 0.63fF $ **FLOATING
C419 a_25198_4511# vssd1 0.58fF $ **FLOATING
C420 a_24757_4399# vssd1 1.43fF $ **FLOATING
C421 a_24591_4399# vssd1 1.81fF $ **FLOATING
C422 a_23013_4399# vssd1 0.23fF $ **FLOATING
C423 a_23523_4765# vssd1 0.61fF $ **FLOATING
C424 a_23691_4667# vssd1 0.82fF $ **FLOATING
C425 a_23098_4765# vssd1 0.63fF $ **FLOATING
C426 a_23266_4511# vssd1 0.58fF $ **FLOATING
C427 a_22825_4399# vssd1 1.43fF $ **FLOATING
C428 a_22659_4399# vssd1 1.81fF $ **FLOATING
C429 _0975_.CLK vssd1 9.39fF $ **FLOATING
C430 a_20897_4399# vssd1 0.23fF $ **FLOATING
C431 a_21407_4765# vssd1 0.61fF $ **FLOATING
C432 a_21575_4667# vssd1 0.82fF $ **FLOATING
C433 a_20982_4765# vssd1 0.63fF $ **FLOATING
C434 a_21150_4511# vssd1 0.58fF $ **FLOATING
C435 a_20709_4399# vssd1 1.43fF $ **FLOATING
C436 a_20543_4399# vssd1 1.81fF $ **FLOATING
C437 a_19605_4649# vssd1 0.21fF $ **FLOATING
C438 a_19521_4649# vssd1 0.17fF $ **FLOATING
C439 _0638_.X vssd1 3.54fF $ **FLOATING
C440 _0956_.Q vssd1 4.56fF $ **FLOATING
C441 a_15929_4399# vssd1 0.23fF $ **FLOATING
C442 a_19439_4399# vssd1 0.97fF $ **FLOATING
C443 _0497_.B2 vssd1 3.84fF $ **FLOATING
C444 a_18059_4399# vssd1 0.62fF $ **FLOATING
C445 a_16439_4765# vssd1 0.61fF $ **FLOATING
C446 a_16607_4667# vssd1 0.82fF $ **FLOATING
C447 a_16014_4765# vssd1 0.63fF $ **FLOATING
C448 a_16182_4511# vssd1 0.58fF $ **FLOATING
C449 a_15741_4399# vssd1 1.43fF $ **FLOATING
C450 _0497_.A1 vssd1 3.03fF $ **FLOATING
C451 a_15575_4399# vssd1 1.81fF $ **FLOATING
C452 _0972_.CLK vssd1 11.23fF $ **FLOATING
C453 a_12709_4399# vssd1 0.23fF $ **FLOATING
C454 a_14655_4399# vssd1 0.62fF $ **FLOATING
C455 a_13219_4765# vssd1 0.61fF $ **FLOATING
C456 a_13387_4667# vssd1 0.82fF $ **FLOATING
C457 a_12794_4765# vssd1 0.63fF $ **FLOATING
C458 a_12962_4511# vssd1 0.58fF $ **FLOATING
C459 a_12521_4399# vssd1 1.43fF $ **FLOATING
C460 _0951_.D vssd1 2.56fF $ **FLOATING
C461 a_12355_4399# vssd1 1.81fF $ **FLOATING
C462 a_9765_4399# vssd1 0.23fF $ **FLOATING
C463 a_10275_4765# vssd1 0.61fF $ **FLOATING
C464 a_10443_4667# vssd1 0.82fF $ **FLOATING
C465 a_9850_4765# vssd1 0.63fF $ **FLOATING
C466 a_10018_4511# vssd1 0.58fF $ **FLOATING
C467 a_9577_4399# vssd1 1.43fF $ **FLOATING
C468 _0959_.D vssd1 4.19fF $ **FLOATING
C469 a_9411_4399# vssd1 1.81fF $ **FLOATING
C470 _0908_.Q vssd1 5.94fF $ **FLOATING
C471 a_7557_4399# vssd1 0.23fF $ **FLOATING
C472 a_8067_4765# vssd1 0.61fF $ **FLOATING
C473 a_8235_4667# vssd1 0.82fF $ **FLOATING
C474 a_7642_4765# vssd1 0.63fF $ **FLOATING
C475 a_7810_4511# vssd1 0.58fF $ **FLOATING
C476 a_7369_4399# vssd1 1.43fF $ **FLOATING
C477 a_7203_4399# vssd1 1.81fF $ **FLOATING
C478 a_4889_4399# vssd1 0.23fF $ **FLOATING
C479 a_5399_4765# vssd1 0.61fF $ **FLOATING
C480 a_5567_4667# vssd1 0.82fF $ **FLOATING
C481 a_4974_4765# vssd1 0.63fF $ **FLOATING
C482 a_5142_4511# vssd1 0.58fF $ **FLOATING
C483 a_4701_4399# vssd1 1.43fF $ **FLOATING
C484 a_4535_4399# vssd1 1.81fF $ **FLOATING
C485 a_2129_4399# vssd1 0.23fF $ **FLOATING
C486 a_2639_4765# vssd1 0.61fF $ **FLOATING
C487 a_2807_4667# vssd1 0.82fF $ **FLOATING
C488 a_2214_4765# vssd1 0.63fF $ **FLOATING
C489 a_2382_4511# vssd1 0.58fF $ **FLOATING
C490 a_1941_4399# vssd1 1.43fF $ **FLOATING
C491 a_1775_4399# vssd1 1.81fF $ **FLOATING
C492 a_27981_4943# vssd1 0.23fF $ **FLOATING
C493 a_25589_4943# vssd1 0.23fF $ **FLOATING
C494 _1040_.Q vssd1 3.28fF $ **FLOATING
C495 a_18505_4943# vssd1 0.23fF $ **FLOATING
C496 a_27804_4943# vssd1 0.50fF $ **FLOATING
C497 a_27698_4943# vssd1 0.58fF $ **FLOATING
C498 a_27521_4943# vssd1 0.50fF $ **FLOATING
C499 fanout23.X vssd1 7.41fF $ **FLOATING
C500 a_27202_4943# vssd1 0.54fF $ **FLOATING
C501 a_26099_4943# vssd1 0.61fF $ **FLOATING
C502 a_26267_4917# vssd1 0.82fF $ **FLOATING
C503 a_25674_4943# vssd1 0.63fF $ **FLOATING
C504 a_25842_4917# vssd1 0.58fF $ **FLOATING
C505 a_25401_4949# vssd1 1.43fF $ **FLOATING
C506 a_25235_4949# vssd1 1.81fF $ **FLOATING
C507 a_19991_5056# vssd1 0.62fF $ **FLOATING
C508 _0632_.B vssd1 4.68fF $ **FLOATING
C509 a_19015_4943# vssd1 0.61fF $ **FLOATING
C510 a_19183_4917# vssd1 0.82fF $ **FLOATING
C511 a_18590_4943# vssd1 0.63fF $ **FLOATING
C512 a_18758_4917# vssd1 0.58fF $ **FLOATING
C513 a_18317_4949# vssd1 1.43fF $ **FLOATING
C514 a_18151_4949# vssd1 1.81fF $ **FLOATING
C515 a_16895_5281# vssd1 0.56fF $ **FLOATING
C516 a_16035_4943# vssd1 0.70fF $ **FLOATING
C517 a_15115_5059# vssd1 0.70fF $ **FLOATING
C518 _0556_.B vssd1 2.90fF $ **FLOATING
C519 _0556_.D vssd1 2.33fF $ **FLOATING
C520 a_12069_4943# vssd1 0.21fF $ **FLOATING
C521 a_13629_4943# vssd1 0.23fF $ **FLOATING
C522 a_10133_4943# vssd1 0.23fF $ **FLOATING
C523 a_8293_4943# vssd1 0.23fF $ **FLOATING
C524 a_4981_4943# vssd1 0.23fF $ **FLOATING
C525 _0910_.Q vssd1 6.07fF $ **FLOATING
C526 a_3049_4943# vssd1 0.23fF $ **FLOATING
C527 _0908_.CLK vssd1 12.16fF $ **FLOATING
C528 a_14139_4943# vssd1 0.61fF $ **FLOATING
C529 a_14307_4917# vssd1 0.82fF $ **FLOATING
C530 a_13714_4943# vssd1 0.63fF $ **FLOATING
C531 a_13882_4917# vssd1 0.58fF $ **FLOATING
C532 a_13441_4949# vssd1 1.43fF $ **FLOATING
C533 a_13275_4949# vssd1 1.81fF $ **FLOATING
C534 a_11987_4943# vssd1 0.80fF $ **FLOATING
C535 _0673_.A1 vssd1 3.41fF $ **FLOATING
C536 a_10643_4943# vssd1 0.61fF $ **FLOATING
C537 a_10811_4917# vssd1 0.82fF $ **FLOATING
C538 a_10218_4943# vssd1 0.63fF $ **FLOATING
C539 a_10386_4917# vssd1 0.58fF $ **FLOATING
C540 a_9945_4949# vssd1 1.43fF $ **FLOATING
C541 _0952_.Q vssd1 3.92fF $ **FLOATING
C542 a_9779_4949# vssd1 1.81fF $ **FLOATING
C543 _0959_.CLK vssd1 10.06fF $ **FLOATING
C544 a_8803_4943# vssd1 0.61fF $ **FLOATING
C545 a_8971_4917# vssd1 0.82fF $ **FLOATING
C546 a_8378_4943# vssd1 0.63fF $ **FLOATING
C547 a_8546_4917# vssd1 0.58fF $ **FLOATING
C548 a_8105_4949# vssd1 1.43fF $ **FLOATING
C549 a_7939_4949# vssd1 1.81fF $ **FLOATING
C550 a_5491_4943# vssd1 0.61fF $ **FLOATING
C551 a_5659_4917# vssd1 0.82fF $ **FLOATING
C552 a_5066_4943# vssd1 0.63fF $ **FLOATING
C553 a_5234_4917# vssd1 0.58fF $ **FLOATING
C554 a_4793_4949# vssd1 1.43fF $ **FLOATING
C555 a_4627_4949# vssd1 1.81fF $ **FLOATING
C556 a_3559_4943# vssd1 0.61fF $ **FLOATING
C557 a_3727_4917# vssd1 0.82fF $ **FLOATING
C558 a_3134_4943# vssd1 0.63fF $ **FLOATING
C559 a_3302_4917# vssd1 0.58fF $ **FLOATING
C560 a_2861_4949# vssd1 1.43fF $ **FLOATING
C561 _0673_.B2 vssd1 5.32fF $ **FLOATING
C562 a_2695_4949# vssd1 1.81fF $ **FLOATING
C563 a_1959_4951# vssd1 0.65fF $ **FLOATING
C564 a_27337_5487# vssd1 0.23fF $ **FLOATING
C565 a_27847_5853# vssd1 0.61fF $ **FLOATING
C566 a_28015_5755# vssd1 0.82fF $ **FLOATING
C567 a_27422_5853# vssd1 0.63fF $ **FLOATING
C568 a_27590_5599# vssd1 0.58fF $ **FLOATING
C569 a_27149_5487# vssd1 1.43fF $ **FLOATING
C570 a_26983_5487# vssd1 1.81fF $ **FLOATING
C571 a_24945_5487# vssd1 0.23fF $ **FLOATING
C572 a_25455_5853# vssd1 0.61fF $ **FLOATING
C573 a_25623_5755# vssd1 0.82fF $ **FLOATING
C574 a_25030_5853# vssd1 0.63fF $ **FLOATING
C575 a_25198_5599# vssd1 0.58fF $ **FLOATING
C576 a_24757_5487# vssd1 1.43fF $ **FLOATING
C577 a_24591_5487# vssd1 1.81fF $ **FLOATING
C578 a_22097_5737# vssd1 0.21fF $ **FLOATING
C579 a_20529_5487# vssd1 0.23fF $ **FLOATING
C580 a_22015_5737# vssd1 0.80fF $ **FLOATING
C581 _1008_.Q vssd1 4.27fF $ **FLOATING
C582 a_21039_5853# vssd1 0.61fF $ **FLOATING
C583 a_21207_5755# vssd1 0.82fF $ **FLOATING
C584 a_20614_5853# vssd1 0.63fF $ **FLOATING
C585 a_20782_5599# vssd1 0.58fF $ **FLOATING
C586 a_20341_5487# vssd1 1.43fF $ **FLOATING
C587 a_20175_5487# vssd1 1.81fF $ **FLOATING
C588 _0631_.B vssd1 5.19fF $ **FLOATING
C589 a_17497_5737# vssd1 0.21fF $ **FLOATING
C590 a_15005_5737# vssd1 0.21fF $ **FLOATING
C591 a_14921_5737# vssd1 0.17fF $ **FLOATING
C592 a_11333_5737# vssd1 0.21fF $ **FLOATING
C593 a_9489_5487# vssd1 0.23fF $ **FLOATING
C594 a_18519_5487# vssd1 0.62fF $ **FLOATING
C595 a_17415_5737# vssd1 0.80fF $ **FLOATING
C596 _0622_.A1 vssd1 3.69fF $ **FLOATING
C597 _0622_.B2 vssd1 7.68fF $ **FLOATING
C598 a_16495_5487# vssd1 0.70fF $ **FLOATING
C599 a_14839_5487# vssd1 0.97fF $ **FLOATING
C600 _0543_.A1 vssd1 4.33fF $ **FLOATING
C601 _0543_.B2 vssd1 3.89fF $ **FLOATING
C602 a_13309_5515# vssd1 0.71fF $ **FLOATING
C603 a_12479_5515# vssd1 0.56fF $ **FLOATING
C604 a_11251_5737# vssd1 0.80fF $ **FLOATING
C605 a_9999_5853# vssd1 0.61fF $ **FLOATING
C606 a_10167_5755# vssd1 0.82fF $ **FLOATING
C607 a_9574_5853# vssd1 0.63fF $ **FLOATING
C608 a_9742_5599# vssd1 0.58fF $ **FLOATING
C609 a_9301_5487# vssd1 1.43fF $ **FLOATING
C610 a_9135_5487# vssd1 1.81fF $ **FLOATING
C611 a_7005_5487# vssd1 0.23fF $ **FLOATING
C612 a_7515_5853# vssd1 0.61fF $ **FLOATING
C613 a_7683_5755# vssd1 0.82fF $ **FLOATING
C614 a_7090_5853# vssd1 0.63fF $ **FLOATING
C615 a_7258_5599# vssd1 0.58fF $ **FLOATING
C616 a_6817_5487# vssd1 1.43fF $ **FLOATING
C617 a_6651_5487# vssd1 1.81fF $ **FLOATING
C618 a_1945_5487# vssd1 0.23fF $ **FLOATING
C619 a_4852_5737# vssd1 0.50fF $ **FLOATING
C620 a_4015_5515# vssd1 0.56fF $ **FLOATING
C621 a_2455_5853# vssd1 0.61fF $ **FLOATING
C622 a_2623_5755# vssd1 0.82fF $ **FLOATING
C623 a_2030_5853# vssd1 0.63fF $ **FLOATING
C624 a_2198_5599# vssd1 0.58fF $ **FLOATING
C625 a_1757_5487# vssd1 1.43fF $ **FLOATING
C626 a_1591_5487# vssd1 1.81fF $ **FLOATING
C627 a_25497_6031# vssd1 0.23fF $ **FLOATING
C628 a_23657_6031# vssd1 0.23fF $ **FLOATING
C629 a_19517_6031# vssd1 0.23fF $ **FLOATING
C630 a_15949_6031# vssd1 0.19fF $ **FLOATING
C631 a_14829_6031# vssd1 0.21fF $ **FLOATING
C632 a_13717_6031# vssd1 0.21fF $ **FLOATING
C633 a_13633_6031# vssd1 0.17fF $ **FLOATING
C634 a_17677_6031# vssd1 0.23fF $ **FLOATING
C635 _0954_.Q vssd1 2.90fF $ **FLOATING
C636 a_12065_6031# vssd1 0.23fF $ **FLOATING
C637 _0902_.Q vssd1 3.95fF $ **FLOATING
C638 a_10041_6031# vssd1 0.23fF $ **FLOATING
C639 _0907_.Q vssd1 3.79fF $ **FLOATING
C640 a_7649_6031# vssd1 0.23fF $ **FLOATING
C641 a_5817_6351# vssd1 0.17fF $ **FLOATING
C642 a_1945_6031# vssd1 0.23fF $ **FLOATING
C643 a_26007_6031# vssd1 0.61fF $ **FLOATING
C644 a_26175_6005# vssd1 0.82fF $ **FLOATING
C645 a_25582_6031# vssd1 0.63fF $ **FLOATING
C646 a_25750_6005# vssd1 0.58fF $ **FLOATING
C647 a_25309_6037# vssd1 1.43fF $ **FLOATING
C648 a_25143_6037# vssd1 1.81fF $ **FLOATING
C649 a_24167_6031# vssd1 0.61fF $ **FLOATING
C650 a_24335_6005# vssd1 0.82fF $ **FLOATING
C651 a_23742_6031# vssd1 0.63fF $ **FLOATING
C652 a_23910_6005# vssd1 0.58fF $ **FLOATING
C653 a_23469_6037# vssd1 1.43fF $ **FLOATING
C654 a_23303_6037# vssd1 1.81fF $ **FLOATING
C655 a_22015_6144# vssd1 0.62fF $ **FLOATING
C656 _0575_.B vssd1 4.61fF $ **FLOATING
C657 a_20027_6031# vssd1 0.61fF $ **FLOATING
C658 a_20195_6005# vssd1 0.82fF $ **FLOATING
C659 a_19602_6031# vssd1 0.63fF $ **FLOATING
C660 a_19770_6005# vssd1 0.58fF $ **FLOATING
C661 a_19329_6037# vssd1 1.43fF $ **FLOATING
C662 a_19163_6037# vssd1 1.81fF $ **FLOATING
C663 a_18187_6031# vssd1 0.61fF $ **FLOATING
C664 a_18355_6005# vssd1 0.82fF $ **FLOATING
C665 a_17762_6031# vssd1 0.63fF $ **FLOATING
C666 a_17930_6005# vssd1 0.58fF $ **FLOATING
C667 a_17489_6037# vssd1 1.43fF $ **FLOATING
C668 a_17323_6037# vssd1 1.81fF $ **FLOATING
C669 _0670_.A1 vssd1 3.15fF $ **FLOATING
C670 _0670_.A2 vssd1 6.05fF $ **FLOATING
C671 a_15812_6005# vssd1 0.85fF $ **FLOATING
C672 a_14747_6031# vssd1 0.80fF $ **FLOATING
C673 _0671_.B2 vssd1 4.84fF $ **FLOATING
C674 a_13551_6031# vssd1 0.97fF $ **FLOATING
C675 _0538_.B2 vssd1 4.53fF $ **FLOATING
C676 _0538_.C1 vssd1 1.53fF $ **FLOATING
C677 a_12575_6031# vssd1 0.61fF $ **FLOATING
C678 a_12743_6005# vssd1 0.82fF $ **FLOATING
C679 a_12150_6031# vssd1 0.63fF $ **FLOATING
C680 a_12318_6005# vssd1 0.58fF $ **FLOATING
C681 a_11877_6037# vssd1 1.43fF $ **FLOATING
C682 _0954_.D vssd1 4.86fF $ **FLOATING
C683 a_11711_6037# vssd1 1.81fF $ **FLOATING
C684 a_10551_6031# vssd1 0.61fF $ **FLOATING
C685 a_10719_6005# vssd1 0.82fF $ **FLOATING
C686 a_10126_6031# vssd1 0.63fF $ **FLOATING
C687 a_10294_6005# vssd1 0.58fF $ **FLOATING
C688 a_9853_6037# vssd1 1.43fF $ **FLOATING
C689 a_9687_6037# vssd1 1.81fF $ **FLOATING
C690 a_8159_6031# vssd1 0.61fF $ **FLOATING
C691 a_8327_6005# vssd1 0.82fF $ **FLOATING
C692 a_7734_6031# vssd1 0.63fF $ **FLOATING
C693 a_7902_6005# vssd1 0.58fF $ **FLOATING
C694 a_7461_6037# vssd1 1.43fF $ **FLOATING
C695 a_7295_6037# vssd1 1.81fF $ **FLOATING
C696 a_5599_6263# vssd1 0.55fF $ **FLOATING
C697 a_4259_6031# vssd1 0.70fF $ **FLOATING
C698 a_3523_6039# vssd1 0.65fF $ **FLOATING
C699 a_2455_6031# vssd1 0.61fF $ **FLOATING
C700 a_2623_6005# vssd1 0.82fF $ **FLOATING
C701 a_2030_6031# vssd1 0.63fF $ **FLOATING
C702 a_2198_6005# vssd1 0.58fF $ **FLOATING
C703 a_1757_6037# vssd1 1.43fF $ **FLOATING
C704 a_1591_6037# vssd1 1.81fF $ **FLOATING
C705 a_27061_6575# vssd1 0.23fF $ **FLOATING
C706 a_27571_6941# vssd1 0.61fF $ **FLOATING
C707 a_27739_6843# vssd1 0.82fF $ **FLOATING
C708 a_27146_6941# vssd1 0.63fF $ **FLOATING
C709 a_27314_6687# vssd1 0.58fF $ **FLOATING
C710 a_26873_6575# vssd1 1.43fF $ **FLOATING
C711 a_26707_6575# vssd1 1.81fF $ **FLOATING
C712 a_25221_6575# vssd1 0.23fF $ **FLOATING
C713 a_25731_6941# vssd1 0.61fF $ **FLOATING
C714 a_25899_6843# vssd1 0.82fF $ **FLOATING
C715 a_25306_6941# vssd1 0.63fF $ **FLOATING
C716 a_25474_6687# vssd1 0.58fF $ **FLOATING
C717 a_25033_6575# vssd1 1.43fF $ **FLOATING
C718 a_24867_6575# vssd1 1.81fF $ **FLOATING
C719 a_23569_6825# vssd1 0.21fF $ **FLOATING
C720 _0669_.X vssd1 3.12fF $ **FLOATING
C721 a_21361_6825# vssd1 0.21fF $ **FLOATING
C722 a_20349_6825# vssd1 0.21fF $ **FLOATING
C723 a_16902_6825# vssd1 0.33fF $ **FLOATING
C724 a_14661_6825# vssd1 0.19fF $ **FLOATING
C725 _0604_.B vssd1 4.21fF $ **FLOATING
C726 a_11693_6825# vssd1 0.21fF $ **FLOATING
C727 a_11609_6825# vssd1 0.17fF $ **FLOATING
C728 a_23487_6825# vssd1 0.80fF $ **FLOATING
C729 _0552_.B2 vssd1 5.53fF $ **FLOATING
C730 a_22325_6603# vssd1 0.71fF $ **FLOATING
C731 a_21279_6825# vssd1 0.80fF $ **FLOATING
C732 _0669_.B2 vssd1 3.51fF $ **FLOATING
C733 a_20267_6825# vssd1 0.80fF $ **FLOATING
C734 _0548_.A1 vssd1 5.08fF $ **FLOATING
C735 _0548_.B2 vssd1 4.02fF $ **FLOATING
C736 a_19471_6603# vssd1 0.56fF $ **FLOATING
C737 _0645_.B2 vssd1 4.34fF $ **FLOATING
C738 _0645_.B1 vssd1 10.39fF $ **FLOATING
C739 a_16745_6549# vssd1 0.72fF $ **FLOATING
C740 a_15793_6603# vssd1 0.71fF $ **FLOATING
C741 a_14524_6549# vssd1 0.85fF $ **FLOATING
C742 a_13367_6575# vssd1 0.62fF $ **FLOATING
C743 a_11527_6575# vssd1 0.97fF $ **FLOATING
C744 _0532_.A2 vssd1 4.83fF $ **FLOATING
C745 _0674_.A1 vssd1 4.60fF $ **FLOATING
C746 _0674_.C1 vssd1 1.68fF $ **FLOATING
C747 a_9919_6740# vssd1 0.52fF $ **FLOATING
C748 a_9135_6575# vssd1 0.65fF $ **FLOATING
C749 a_6821_6575# vssd1 0.23fF $ **FLOATING
C750 a_7331_6941# vssd1 0.61fF $ **FLOATING
C751 a_7499_6843# vssd1 0.82fF $ **FLOATING
C752 a_6906_6941# vssd1 0.63fF $ **FLOATING
C753 a_7074_6687# vssd1 0.58fF $ **FLOATING
C754 a_6633_6575# vssd1 1.43fF $ **FLOATING
C755 a_6467_6575# vssd1 1.81fF $ **FLOATING
C756 a_1945_6575# vssd1 0.23fF $ **FLOATING
C757 a_2455_6941# vssd1 0.61fF $ **FLOATING
C758 a_2623_6843# vssd1 0.82fF $ **FLOATING
C759 a_2030_6941# vssd1 0.63fF $ **FLOATING
C760 a_2198_6687# vssd1 0.58fF $ **FLOATING
C761 a_1757_6575# vssd1 1.43fF $ **FLOATING
C762 a_1591_6575# vssd1 1.81fF $ **FLOATING
C763 a_25589_7119# vssd1 0.23fF $ **FLOATING
C764 a_20257_7119# vssd1 0.21fF $ **FLOATING
C765 a_22921_7119# vssd1 0.23fF $ **FLOATING
C766 a_17029_7119# vssd1 0.21fF $ **FLOATING
C767 a_16945_7119# vssd1 0.17fF $ **FLOATING
C768 a_26099_7119# vssd1 0.61fF $ **FLOATING
C769 a_26267_7093# vssd1 0.82fF $ **FLOATING
C770 a_25674_7119# vssd1 0.63fF $ **FLOATING
C771 a_25842_7093# vssd1 0.58fF $ **FLOATING
C772 a_25401_7125# vssd1 1.43fF $ **FLOATING
C773 a_25235_7125# vssd1 1.81fF $ **FLOATING
C774 a_23431_7119# vssd1 0.61fF $ **FLOATING
C775 a_23599_7093# vssd1 0.82fF $ **FLOATING
C776 a_23006_7119# vssd1 0.63fF $ **FLOATING
C777 a_23174_7093# vssd1 0.58fF $ **FLOATING
C778 a_22733_7125# vssd1 1.43fF $ **FLOATING
C779 _1045_.D vssd1 4.53fF $ **FLOATING
C780 a_22567_7125# vssd1 1.81fF $ **FLOATING
C781 a_20175_7119# vssd1 0.80fF $ **FLOATING
C782 _0649_.B2 vssd1 3.16fF $ **FLOATING
C783 a_18645_7457# vssd1 0.71fF $ **FLOATING
C784 a_16863_7119# vssd1 0.97fF $ **FLOATING
C785 _0672_.C1 vssd1 1.67fF $ **FLOATING
C786 a_15671_7235# vssd1 0.70fF $ **FLOATING
C787 a_15565_7235# vssd1 0.43fF $ **FLOATING
C788 _0642_.D_N vssd1 3.80fF $ **FLOATING
C789 a_14011_7235# vssd1 0.70fF $ **FLOATING
C790 _0544_.B vssd1 0.99fF $ **FLOATING
C791 _0544_.C vssd1 1.18fF $ **FLOATING
C792 _0544_.D vssd1 1.93fF $ **FLOATING
C793 a_12245_7119# vssd1 0.21fF $ **FLOATING
C794 a_12161_7119# vssd1 0.17fF $ **FLOATING
C795 _0642_.C vssd1 1.95fF $ **FLOATING
C796 a_10335_7439# vssd1 0.27fF $ **FLOATING
C797 a_5727_7119# vssd1 0.25fF $ **FLOATING
C798 a_8661_7119# vssd1 0.23fF $ **FLOATING
C799 input2.X vssd1 1.89fF $ **FLOATING
C800 a_13183_7232# vssd1 0.62fF $ **FLOATING
C801 _0611_.B vssd1 6.77fF $ **FLOATING
C802 a_12079_7119# vssd1 0.97fF $ **FLOATING
C803 _0637_.A1 vssd1 4.15fF $ **FLOATING
C804 _0566_.A1 vssd1 4.89fF $ **FLOATING
C805 _0566_.B1 vssd1 3.78fF $ **FLOATING
C806 a_10198_7351# vssd1 0.60fF $ **FLOATING
C807 a_9171_7119# vssd1 0.61fF $ **FLOATING
C808 a_9339_7093# vssd1 0.82fF $ **FLOATING
C809 a_8746_7119# vssd1 0.63fF $ **FLOATING
C810 a_8914_7093# vssd1 0.58fF $ **FLOATING
C811 a_8473_7125# vssd1 1.43fF $ **FLOATING
C812 a_8307_7125# vssd1 1.81fF $ **FLOATING
C813 _0888_.CLK vssd1 10.04fF $ **FLOATING
C814 a_5509_7093# vssd1 0.55fF $ **FLOATING
C815 a_2787_7119# vssd1 0.70fF $ **FLOATING
C816 io_in[2] vssd1 1.88fF
C817 a_1639_7338# vssd1 0.52fF $ **FLOATING
C818 a_27337_7663# vssd1 0.23fF $ **FLOATING
C819 a_27847_8029# vssd1 0.61fF $ **FLOATING
C820 a_28015_7931# vssd1 0.82fF $ **FLOATING
C821 a_27422_8029# vssd1 0.63fF $ **FLOATING
C822 a_27590_7775# vssd1 0.58fF $ **FLOATING
C823 a_27149_7663# vssd1 1.43fF $ **FLOATING
C824 a_26983_7663# vssd1 1.81fF $ **FLOATING
C825 a_25405_7663# vssd1 0.23fF $ **FLOATING
C826 a_25915_8029# vssd1 0.61fF $ **FLOATING
C827 a_26083_7931# vssd1 0.82fF $ **FLOATING
C828 a_25490_8029# vssd1 0.63fF $ **FLOATING
C829 a_25658_7775# vssd1 0.58fF $ **FLOATING
C830 a_25217_7663# vssd1 1.43fF $ **FLOATING
C831 a_25051_7663# vssd1 1.81fF $ **FLOATING
C832 a_22917_7913# vssd1 0.21fF $ **FLOATING
C833 a_22833_7913# vssd1 0.17fF $ **FLOATING
C834 a_21813_7913# vssd1 0.21fF $ **FLOATING
C835 a_21729_7913# vssd1 0.17fF $ **FLOATING
C836 a_20161_7663# vssd1 0.23fF $ **FLOATING
C837 a_22751_7663# vssd1 0.97fF $ **FLOATING
C838 _0618_.B2 vssd1 4.11fF $ **FLOATING
C839 _0618_.C1 vssd1 1.48fF $ **FLOATING
C840 a_21647_7663# vssd1 0.97fF $ **FLOATING
C841 _1003_.Q vssd1 3.89fF $ **FLOATING
C842 _0516_.B1 vssd1 9.23fF $ **FLOATING
C843 a_20671_8029# vssd1 0.61fF $ **FLOATING
C844 a_20839_7931# vssd1 0.82fF $ **FLOATING
C845 a_20246_8029# vssd1 0.63fF $ **FLOATING
C846 a_20414_7775# vssd1 0.58fF $ **FLOATING
C847 a_19973_7663# vssd1 1.43fF $ **FLOATING
C848 a_19807_7663# vssd1 1.81fF $ **FLOATING
C849 _1030_.CLK vssd1 11.98fF $ **FLOATING
C850 a_18456_7913# vssd1 0.26fF $ **FLOATING
C851 _0634_.X vssd1 1.94fF $ **FLOATING
C852 _0549_.X vssd1 2.22fF $ **FLOATING
C853 a_16293_7913# vssd1 0.21fF $ **FLOATING
C854 a_16209_7913# vssd1 0.17fF $ **FLOATING
C855 a_14641_7663# vssd1 0.23fF $ **FLOATING
C856 _0634_.B1 vssd1 1.72fF $ **FLOATING
C857 _0634_.C1 vssd1 2.71fF $ **FLOATING
C858 a_18025_7809# vssd1 0.67fF $ **FLOATING
C859 a_16127_7663# vssd1 0.97fF $ **FLOATING
C860 _0549_.B2 vssd1 5.66fF $ **FLOATING
C861 _0549_.C1 vssd1 3.02fF $ **FLOATING
C862 a_15151_8029# vssd1 0.61fF $ **FLOATING
C863 a_15319_7931# vssd1 0.82fF $ **FLOATING
C864 a_14726_8029# vssd1 0.63fF $ **FLOATING
C865 a_14894_7775# vssd1 0.58fF $ **FLOATING
C866 a_14453_7663# vssd1 1.43fF $ **FLOATING
C867 a_14287_7663# vssd1 1.81fF $ **FLOATING
C868 a_12797_7913# vssd1 0.21fF $ **FLOATING
C869 a_12713_7913# vssd1 0.17fF $ **FLOATING
C870 _0901_.Q vssd1 3.98fF $ **FLOATING
C871 a_9581_7663# vssd1 0.23fF $ **FLOATING
C872 a_12631_7663# vssd1 0.97fF $ **FLOATING
C873 _0646_.A1 vssd1 6.27fF $ **FLOATING
C874 _0646_.C1 vssd1 2.71fF $ **FLOATING
C875 a_10091_8029# vssd1 0.61fF $ **FLOATING
C876 a_10259_7931# vssd1 0.82fF $ **FLOATING
C877 a_9666_8029# vssd1 0.63fF $ **FLOATING
C878 a_9834_7775# vssd1 0.58fF $ **FLOATING
C879 a_9393_7663# vssd1 1.43fF $ **FLOATING
C880 a_9227_7663# vssd1 1.81fF $ **FLOATING
C881 _1028_.CLK vssd1 12.54fF $ **FLOATING
C882 a_6815_7913# vssd1 0.41fF $ **FLOATING
C883 a_6376_7913# vssd1 0.32fF $ **FLOATING
C884 a_4259_7669# vssd1 0.48fF $ **FLOATING
C885 input3.X vssd1 3.41fF $ **FLOATING
C886 a_4451_7913# vssd1 0.48fF $ **FLOATING
C887 io_in[3] vssd1 1.26fF
C888 a_1639_7828# vssd1 0.52fF $ **FLOATING
C889 a_25129_8207# vssd1 0.23fF $ **FLOATING
C890 _1031_.Q vssd1 5.35fF $ **FLOATING
C891 a_23105_8207# vssd1 0.23fF $ **FLOATING
C892 a_19429_8207# vssd1 0.21fF $ **FLOATING
C893 a_18065_8207# vssd1 0.19fF $ **FLOATING
C894 _0515_.X vssd1 1.53fF $ **FLOATING
C895 a_25639_8207# vssd1 0.61fF $ **FLOATING
C896 a_25807_8181# vssd1 0.82fF $ **FLOATING
C897 a_25214_8207# vssd1 0.63fF $ **FLOATING
C898 a_25382_8181# vssd1 0.58fF $ **FLOATING
C899 a_24941_8213# vssd1 1.43fF $ **FLOATING
C900 a_24775_8213# vssd1 1.81fF $ **FLOATING
C901 a_23615_8207# vssd1 0.61fF $ **FLOATING
C902 a_23783_8181# vssd1 0.82fF $ **FLOATING
C903 a_23190_8207# vssd1 0.63fF $ **FLOATING
C904 a_23358_8181# vssd1 0.58fF $ **FLOATING
C905 a_22917_8213# vssd1 1.43fF $ **FLOATING
C906 a_22751_8213# vssd1 1.81fF $ **FLOATING
C907 _1033_.CLK vssd1 9.60fF $ **FLOATING
C908 a_22015_8215# vssd1 0.65fF $ **FLOATING
C909 fanout24.A vssd1 12.10fF $ **FLOATING
C910 a_20393_8545# vssd1 0.71fF $ **FLOATING
C911 a_19347_8207# vssd1 0.80fF $ **FLOATING
C912 _0515_.B1 vssd1 11.16fF $ **FLOATING
C913 _0515_.B2 vssd1 4.60fF $ **FLOATING
C914 _0587_.C1 vssd1 5.11fF $ **FLOATING
C915 a_17928_8181# vssd1 0.85fF $ **FLOATING
C916 a_15391_8323# vssd1 0.70fF $ **FLOATING
C917 _0675_.B vssd1 1.59fF $ **FLOATING
C918 _0675_.C vssd1 1.87fF $ **FLOATING
C919 _0675_.D vssd1 2.80fF $ **FLOATING
C920 a_6749_8207# vssd1 0.19fF $ **FLOATING
C921 a_12065_8207# vssd1 0.23fF $ **FLOATING
C922 a_7663_8527# vssd1 0.18fF $ **FLOATING
C923 a_5510_8527# vssd1 0.20fF $ **FLOATING
C924 a_13551_8215# vssd1 0.65fF $ **FLOATING
C925 a_12575_8207# vssd1 0.61fF $ **FLOATING
C926 a_12743_8181# vssd1 0.82fF $ **FLOATING
C927 a_12150_8207# vssd1 0.63fF $ **FLOATING
C928 a_12318_8181# vssd1 0.58fF $ **FLOATING
C929 a_11877_8213# vssd1 1.43fF $ **FLOATING
C930 _0916_.D vssd1 5.00fF $ **FLOATING
C931 a_11711_8213# vssd1 1.81fF $ **FLOATING
C932 _0677_.A1 vssd1 4.17fF $ **FLOATING
C933 a_6612_8181# vssd1 0.85fF $ **FLOATING
C934 _0694_.A2 vssd1 3.52fF $ **FLOATING
C935 _0694_.A1 vssd1 2.29fF $ **FLOATING
C936 a_5325_8181# vssd1 0.89fF $ **FLOATING
C937 a_27245_8751# vssd1 0.23fF $ **FLOATING
C938 a_27755_9117# vssd1 0.61fF $ **FLOATING
C939 a_27923_9019# vssd1 0.82fF $ **FLOATING
C940 a_27330_9117# vssd1 0.63fF $ **FLOATING
C941 a_27498_8863# vssd1 0.58fF $ **FLOATING
C942 a_27057_8751# vssd1 1.43fF $ **FLOATING
C943 a_26891_8751# vssd1 1.81fF $ **FLOATING
C944 a_25405_8751# vssd1 0.23fF $ **FLOATING
C945 a_25915_9117# vssd1 0.61fF $ **FLOATING
C946 a_26083_9019# vssd1 0.82fF $ **FLOATING
C947 a_25490_9117# vssd1 0.63fF $ **FLOATING
C948 a_25658_8863# vssd1 0.58fF $ **FLOATING
C949 a_25217_8751# vssd1 1.43fF $ **FLOATING
C950 a_25051_8751# vssd1 1.81fF $ **FLOATING
C951 a_23013_8751# vssd1 0.23fF $ **FLOATING
C952 a_23523_9117# vssd1 0.61fF $ **FLOATING
C953 a_23691_9019# vssd1 0.82fF $ **FLOATING
C954 a_23098_9117# vssd1 0.63fF $ **FLOATING
C955 a_23266_8863# vssd1 0.58fF $ **FLOATING
C956 a_22825_8751# vssd1 1.43fF $ **FLOATING
C957 a_22659_8751# vssd1 1.81fF $ **FLOATING
C958 _0941_.Q vssd1 3.37fF $ **FLOATING
C959 a_21173_8751# vssd1 0.23fF $ **FLOATING
C960 a_21683_9117# vssd1 0.61fF $ **FLOATING
C961 a_21851_9019# vssd1 0.82fF $ **FLOATING
C962 a_21258_9117# vssd1 0.63fF $ **FLOATING
C963 a_21426_8863# vssd1 0.58fF $ **FLOATING
C964 a_20985_8751# vssd1 1.43fF $ **FLOATING
C965 a_20819_8751# vssd1 1.81fF $ **FLOATING
C966 _0517_.D vssd1 2.34fF $ **FLOATING
C967 _0517_.B vssd1 2.78fF $ **FLOATING
C968 _0553_.X vssd1 3.78fF $ **FLOATING
C969 a_18409_9001# vssd1 0.21fF $ **FLOATING
C970 a_18325_9001# vssd1 0.17fF $ **FLOATING
C971 a_16853_9001# vssd1 0.21fF $ **FLOATING
C972 _0595_.D vssd1 4.57fF $ **FLOATING
C973 _0587_.X vssd1 1.83fF $ **FLOATING
C974 a_15052_9001# vssd1 0.26fF $ **FLOATING
C975 a_19439_9001# vssd1 0.70fF $ **FLOATING
C976 a_18243_8751# vssd1 0.97fF $ **FLOATING
C977 _0553_.C1 vssd1 4.08fF $ **FLOATING
C978 a_16771_9001# vssd1 0.80fF $ **FLOATING
C979 _0615_.A1 vssd1 3.67fF $ **FLOATING
C980 a_15759_9001# vssd1 0.70fF $ **FLOATING
C981 _0601_.B1 vssd1 2.64fF $ **FLOATING
C982 a_14621_8897# vssd1 0.67fF $ **FLOATING
C983 a_13459_8751# vssd1 0.65fF $ **FLOATING
C984 _0535_.X vssd1 8.14fF $ **FLOATING
C985 a_12355_8751# vssd1 0.89fF $ **FLOATING
C986 a_11435_8751# vssd1 1.20fF $ **FLOATING
C987 a_9411_8751# vssd1 0.65fF $ **FLOATING
C988 a_6549_9001# vssd1 0.23fF $ **FLOATING
C989 a_4439_9001# vssd1 0.25fF $ **FLOATING
C990 a_1945_8751# vssd1 0.23fF $ **FLOATING
C991 a_6423_8903# vssd1 0.95fF $ **FLOATING
C992 a_5128_9001# vssd1 0.50fF $ **FLOATING
C993 _0695_.A2 vssd1 2.95fF $ **FLOATING
C994 _0695_.A1 vssd1 3.68fF $ **FLOATING
C995 a_4221_8725# vssd1 0.55fF $ **FLOATING
C996 a_2455_9117# vssd1 0.61fF $ **FLOATING
C997 a_2623_9019# vssd1 0.82fF $ **FLOATING
C998 a_2030_9117# vssd1 0.63fF $ **FLOATING
C999 a_2198_8863# vssd1 0.58fF $ **FLOATING
C1000 a_1757_8751# vssd1 1.43fF $ **FLOATING
C1001 a_1591_8751# vssd1 1.81fF $ **FLOATING
C1002 a_25309_9295# vssd1 0.21fF $ **FLOATING
C1003 a_25225_9295# vssd1 0.17fF $ **FLOATING
C1004 a_23657_9295# vssd1 0.23fF $ **FLOATING
C1005 a_19846_9295# vssd1 0.33fF $ **FLOATING
C1006 a_15563_9295# vssd1 0.35fF $ **FLOATING
C1007 a_15369_9295# vssd1 0.25fF $ **FLOATING
C1008 a_15115_9295# vssd1 0.38fF $ **FLOATING
C1009 _0590_.X vssd1 3.76fF $ **FLOATING
C1010 _1027_.Q vssd1 2.75fF $ **FLOATING
C1011 a_13169_9295# vssd1 0.23fF $ **FLOATING
C1012 _0491_.X vssd1 11.00fF $ **FLOATING
C1013 a_9673_9295# vssd1 0.23fF $ **FLOATING
C1014 a_8393_9615# vssd1 0.17fF $ **FLOATING
C1015 _0689_.X vssd1 4.21fF $ **FLOATING
C1016 _0681_.X vssd1 4.46fF $ **FLOATING
C1017 a_5445_9295# vssd1 0.18fF $ **FLOATING
C1018 a_4530_9295# vssd1 0.19fF $ **FLOATING
C1019 a_1945_9295# vssd1 0.22fF $ **FLOATING
C1020 a_25143_9295# vssd1 0.97fF $ **FLOATING
C1021 _0665_.B2 vssd1 4.76fF $ **FLOATING
C1022 a_24167_9295# vssd1 0.61fF $ **FLOATING
C1023 a_24335_9269# vssd1 0.82fF $ **FLOATING
C1024 a_23742_9295# vssd1 0.63fF $ **FLOATING
C1025 a_23910_9269# vssd1 0.58fF $ **FLOATING
C1026 a_23469_9301# vssd1 1.43fF $ **FLOATING
C1027 a_23303_9301# vssd1 1.81fF $ **FLOATING
C1028 _0623_.D vssd1 4.19fF $ **FLOATING
C1029 a_20761_9633# vssd1 0.71fF $ **FLOATING
C1030 _0590_.B2 vssd1 3.06fF $ **FLOATING
C1031 a_19689_9269# vssd1 0.72fF $ **FLOATING
C1032 _0652_.C vssd1 2.45fF $ **FLOATING
C1033 _0652_.A vssd1 2.03fF $ **FLOATING
C1034 a_13679_9295# vssd1 0.61fF $ **FLOATING
C1035 a_13847_9269# vssd1 0.82fF $ **FLOATING
C1036 a_13254_9295# vssd1 0.63fF $ **FLOATING
C1037 a_13422_9269# vssd1 0.58fF $ **FLOATING
C1038 a_12981_9301# vssd1 1.43fF $ **FLOATING
C1039 a_12815_9301# vssd1 1.81fF $ **FLOATING
C1040 a_11929_9633# vssd1 0.71fF $ **FLOATING
C1041 a_10183_9295# vssd1 0.61fF $ **FLOATING
C1042 a_10351_9269# vssd1 0.82fF $ **FLOATING
C1043 a_9758_9295# vssd1 0.63fF $ **FLOATING
C1044 a_9926_9269# vssd1 0.58fF $ **FLOATING
C1045 a_9485_9301# vssd1 1.43fF $ **FLOATING
C1046 a_9319_9301# vssd1 1.81fF $ **FLOATING
C1047 a_8175_9527# vssd1 0.55fF $ **FLOATING
C1048 a_7203_9408# vssd1 0.62fF $ **FLOATING
C1049 _0710_.A2 vssd1 2.58fF $ **FLOATING
C1050 _0710_.A1 vssd1 1.77fF $ **FLOATING
C1051 _0710_.B1 vssd1 3.08fF $ **FLOATING
C1052 _0710_.B2 vssd1 2.30fF $ **FLOATING
C1053 a_4447_9295# vssd1 0.63fF $ **FLOATING
C1054 a_4259_9295# vssd1 0.55fF $ **FLOATING
C1055 _0702_.B1_N vssd1 3.16fF $ **FLOATING
C1056 a_2455_9295# vssd1 0.60fF $ **FLOATING
C1057 a_2626_9269# vssd1 1.41fF $ **FLOATING
C1058 a_2039_9295# vssd1 0.63fF $ **FLOATING
C1059 a_2198_9269# vssd1 0.59fF $ **FLOATING
C1060 a_1757_9301# vssd1 1.39fF $ **FLOATING
C1061 _1084_.D vssd1 5.39fF $ **FLOATING
C1062 a_1591_9301# vssd1 1.77fF $ **FLOATING
C1063 a_27337_9839# vssd1 0.23fF $ **FLOATING
C1064 a_27847_10205# vssd1 0.61fF $ **FLOATING
C1065 a_28015_10107# vssd1 0.82fF $ **FLOATING
C1066 a_27422_10205# vssd1 0.63fF $ **FLOATING
C1067 a_27590_9951# vssd1 0.58fF $ **FLOATING
C1068 a_27149_9839# vssd1 1.43fF $ **FLOATING
C1069 a_26983_9839# vssd1 1.81fF $ **FLOATING
C1070 a_25497_9839# vssd1 0.23fF $ **FLOATING
C1071 a_26007_10205# vssd1 0.61fF $ **FLOATING
C1072 a_26175_10107# vssd1 0.82fF $ **FLOATING
C1073 a_25582_10205# vssd1 0.63fF $ **FLOATING
C1074 a_25750_9951# vssd1 0.58fF $ **FLOATING
C1075 a_25309_9839# vssd1 1.43fF $ **FLOATING
C1076 a_25143_9839# vssd1 1.81fF $ **FLOATING
C1077 a_23201_10089# vssd1 0.21fF $ **FLOATING
C1078 _0666_.D vssd1 2.61fF $ **FLOATING
C1079 _0666_.B vssd1 4.24fF $ **FLOATING
C1080 _0633_.X vssd1 2.64fF $ **FLOATING
C1081 _0589_.X vssd1 2.94fF $ **FLOATING
C1082 a_19605_10089# vssd1 0.21fF $ **FLOATING
C1083 a_19521_10089# vssd1 0.17fF $ **FLOATING
C1084 _0624_.C vssd1 3.80fF $ **FLOATING
C1085 a_17865_9845# vssd1 0.43fF $ **FLOATING
C1086 _0624_.D_N vssd1 3.29fF $ **FLOATING
C1087 a_14641_9839# vssd1 0.23fF $ **FLOATING
C1088 a_23119_10089# vssd1 0.80fF $ **FLOATING
C1089 _1069_.Q vssd1 5.27fF $ **FLOATING
C1090 _0488_.B2 vssd1 2.32fF $ **FLOATING
C1091 a_21831_10089# vssd1 0.70fF $ **FLOATING
C1092 a_20543_9839# vssd1 0.62fF $ **FLOATING
C1093 a_19439_9839# vssd1 0.97fF $ **FLOATING
C1094 a_17971_10089# vssd1 0.70fF $ **FLOATING
C1095 _0666_.X vssd1 3.37fF $ **FLOATING
C1096 _0676_.B vssd1 1.30fF $ **FLOATING
C1097 a_15151_10205# vssd1 0.61fF $ **FLOATING
C1098 a_15319_10107# vssd1 0.82fF $ **FLOATING
C1099 a_14726_10205# vssd1 0.63fF $ **FLOATING
C1100 a_14894_9951# vssd1 0.58fF $ **FLOATING
C1101 a_14453_9839# vssd1 1.43fF $ **FLOATING
C1102 _0961_.D vssd1 6.02fF $ **FLOATING
C1103 a_14287_9839# vssd1 1.81fF $ **FLOATING
C1104 a_10084_9839# vssd1 0.22fF $ **FLOATING
C1105 a_9993_9839# vssd1 0.12fF $ **FLOATING
C1106 a_9135_9839# vssd1 0.18fF $ **FLOATING
C1107 a_11789_9839# vssd1 0.23fF $ **FLOATING
C1108 a_12299_10205# vssd1 0.61fF $ **FLOATING
C1109 a_12467_10107# vssd1 0.82fF $ **FLOATING
C1110 a_11874_10205# vssd1 0.63fF $ **FLOATING
C1111 a_12042_9951# vssd1 0.58fF $ **FLOATING
C1112 a_11601_9839# vssd1 1.43fF $ **FLOATING
C1113 a_11435_9839# vssd1 1.81fF $ **FLOATING
C1114 a_4253_9839# vssd1 0.17fF $ **FLOATING
C1115 _0680_.Y vssd1 4.43fF $ **FLOATING
C1116 a_7457_10089# vssd1 0.33fF $ **FLOATING
C1117 a_7203_10089# vssd1 0.38fF $ **FLOATING
C1118 _0657_.X vssd1 2.34fF $ **FLOATING
C1119 a_9895_10089# vssd1 0.87fF $ **FLOATING
C1120 _0545_.A1 vssd1 5.32fF $ **FLOATING
C1121 _0545_.B2 vssd1 3.95fF $ **FLOATING
C1122 _0545_.B1 vssd1 5.64fF $ **FLOATING
C1123 _0653_.A1 vssd1 3.06fF $ **FLOATING
C1124 a_6416_10089# vssd1 0.50fF $ **FLOATING
C1125 a_4035_9813# vssd1 0.55fF $ **FLOATING
C1126 _0696_.A1 vssd1 3.18fF $ **FLOATING
C1127 a_1591_9839# vssd1 0.65fF $ **FLOATING
C1128 io_in[4] vssd1 1.27fF
C1129 a_27249_10383# vssd1 0.21fF $ **FLOATING
C1130 a_25589_10383# vssd1 0.23fF $ **FLOATING
C1131 a_23385_10383# vssd1 0.21fF $ **FLOATING
C1132 a_20717_10383# vssd1 0.21fF $ **FLOATING
C1133 _0621_.X vssd1 1.65fF $ **FLOATING
C1134 _0651_.X vssd1 4.15fF $ **FLOATING
C1135 a_27167_10383# vssd1 0.80fF $ **FLOATING
C1136 _0647_.B2 vssd1 2.62fF $ **FLOATING
C1137 a_26099_10383# vssd1 0.61fF $ **FLOATING
C1138 a_26267_10357# vssd1 0.82fF $ **FLOATING
C1139 a_25674_10383# vssd1 0.63fF $ **FLOATING
C1140 a_25842_10357# vssd1 0.58fF $ **FLOATING
C1141 a_25401_10389# vssd1 1.43fF $ **FLOATING
C1142 _1006_.D vssd1 6.42fF $ **FLOATING
C1143 a_25235_10389# vssd1 1.81fF $ **FLOATING
C1144 a_24315_10496# vssd1 0.62fF $ **FLOATING
C1145 _0573_.B vssd1 4.71fF $ **FLOATING
C1146 a_23303_10383# vssd1 0.80fF $ **FLOATING
C1147 _0621_.A1 vssd1 4.11fF $ **FLOATING
C1148 _0621_.B2 vssd1 3.86fF $ **FLOATING
C1149 a_22199_10499# vssd1 0.70fF $ **FLOATING
C1150 _0647_.X vssd1 3.07fF $ **FLOATING
C1151 _0651_.C vssd1 2.61fF $ **FLOATING
C1152 _0531_.X vssd1 4.82fF $ **FLOATING
C1153 a_17217_10383# vssd1 0.23fF $ **FLOATING
C1154 a_15236_10383# vssd1 0.26fF $ **FLOATING
C1155 a_8116_10383# vssd1 0.17fF $ **FLOATING
C1156 a_6559_10383# vssd1 0.44fF $ **FLOATING
C1157 a_13261_10383# vssd1 0.23fF $ **FLOATING
C1158 a_10325_10703# vssd1 0.17fF $ **FLOATING
C1159 a_9313_10703# vssd1 0.17fF $ **FLOATING
C1160 a_8033_10703# vssd1 0.42fF $ **FLOATING
C1161 _0656_.Y vssd1 4.41fF $ **FLOATING
C1162 a_5731_10703# vssd1 0.18fF $ **FLOATING
C1163 clkbuf_1_0__f_io_in[0].X vssd1 15.85fF $ **FLOATING
C1164 a_20635_10383# vssd1 0.80fF $ **FLOATING
C1165 _0531_.A1 vssd1 6.83fF $ **FLOATING
C1166 a_19439_10496# vssd1 0.62fF $ **FLOATING
C1167 _0607_.B vssd1 5.56fF $ **FLOATING
C1168 a_17727_10383# vssd1 0.61fF $ **FLOATING
C1169 a_17895_10357# vssd1 0.82fF $ **FLOATING
C1170 a_17302_10383# vssd1 0.63fF $ **FLOATING
C1171 a_17470_10357# vssd1 0.58fF $ **FLOATING
C1172 a_17029_10389# vssd1 1.43fF $ **FLOATING
C1173 _0983_.D vssd1 5.11fF $ **FLOATING
C1174 a_16863_10389# vssd1 1.81fF $ **FLOATING
C1175 a_15975_10721# vssd1 0.56fF $ **FLOATING
C1176 _0613_.A1 vssd1 4.89fF $ **FLOATING
C1177 _0613_.C1 vssd1 2.67fF $ **FLOATING
C1178 a_14805_10357# vssd1 0.67fF $ **FLOATING
C1179 a_13771_10383# vssd1 0.61fF $ **FLOATING
C1180 a_13939_10357# vssd1 0.82fF $ **FLOATING
C1181 a_13346_10383# vssd1 0.63fF $ **FLOATING
C1182 a_13514_10357# vssd1 0.58fF $ **FLOATING
C1183 a_13073_10389# vssd1 1.43fF $ **FLOATING
C1184 a_12907_10389# vssd1 1.81fF $ **FLOATING
C1185 _0625_.A1 vssd1 3.69fF $ **FLOATING
C1186 a_10107_10615# vssd1 0.55fF $ **FLOATING
C1187 _0596_.A1 vssd1 4.76fF $ **FLOATING
C1188 a_9095_10615# vssd1 0.55fF $ **FLOATING
C1189 _0679_.A2 vssd1 2.61fF $ **FLOATING
C1190 _0679_.A1 vssd1 5.23fF $ **FLOATING
C1191 a_4811_10383# vssd1 0.99fF $ **FLOATING
C1192 a_2686_10383# vssd1 4.03fF $ **FLOATING
C1193 _1064_.Q vssd1 4.52fF $ **FLOATING
C1194 a_26325_10927# vssd1 0.23fF $ **FLOATING
C1195 a_26835_11293# vssd1 0.61fF $ **FLOATING
C1196 a_27003_11195# vssd1 0.82fF $ **FLOATING
C1197 a_26410_11293# vssd1 0.63fF $ **FLOATING
C1198 a_26578_11039# vssd1 0.58fF $ **FLOATING
C1199 a_26137_10927# vssd1 1.43fF $ **FLOATING
C1200 a_25971_10927# vssd1 1.81fF $ **FLOATING
C1201 a_24673_11177# vssd1 0.21fF $ **FLOATING
C1202 _0506_.X vssd1 3.09fF $ **FLOATING
C1203 a_22825_11177# vssd1 0.21fF $ **FLOATING
C1204 a_22741_11177# vssd1 0.17fF $ **FLOATING
C1205 a_21134_11177# vssd1 0.33fF $ **FLOATING
C1206 _0496_.X vssd1 4.02fF $ **FLOATING
C1207 _1029_.Q vssd1 4.22fF $ **FLOATING
C1208 a_17861_10927# vssd1 0.23fF $ **FLOATING
C1209 a_24591_11177# vssd1 0.80fF $ **FLOATING
C1210 _0562_.A1 vssd1 3.74fF $ **FLOATING
C1211 a_23763_10927# vssd1 0.70fF $ **FLOATING
C1212 a_22659_10927# vssd1 0.97fF $ **FLOATING
C1213 _0506_.A2 vssd1 9.51fF $ **FLOATING
C1214 _0506_.A1 vssd1 4.04fF $ **FLOATING
C1215 a_20977_10901# vssd1 0.72fF $ **FLOATING
C1216 a_20025_10955# vssd1 0.71fF $ **FLOATING
C1217 a_18371_11293# vssd1 0.61fF $ **FLOATING
C1218 a_18539_11195# vssd1 0.82fF $ **FLOATING
C1219 a_17946_11293# vssd1 0.63fF $ **FLOATING
C1220 a_18114_11039# vssd1 0.58fF $ **FLOATING
C1221 a_17673_10927# vssd1 1.43fF $ **FLOATING
C1222 a_17507_10927# vssd1 1.81fF $ **FLOATING
C1223 a_16685_11177# vssd1 0.19fF $ **FLOATING
C1224 _0616_.X vssd1 1.81fF $ **FLOATING
C1225 _0614_.X vssd1 2.12fF $ **FLOATING
C1226 _0614_.A vssd1 2.07fF $ **FLOATING
C1227 _0614_.D vssd1 1.11fF $ **FLOATING
C1228 a_14655_11177# vssd1 0.39fF $ **FLOATING
C1229 _0899_.Q vssd1 4.04fF $ **FLOATING
C1230 a_9781_10927# vssd1 0.18fF $ **FLOATING
C1231 a_10777_10927# vssd1 0.23fF $ **FLOATING
C1232 _0616_.B1 vssd1 1.55fF $ **FLOATING
C1233 a_16548_10901# vssd1 0.85fF $ **FLOATING
C1234 a_15483_11177# vssd1 0.70fF $ **FLOATING
C1235 a_11287_11293# vssd1 0.61fF $ **FLOATING
C1236 a_11455_11195# vssd1 0.82fF $ **FLOATING
C1237 a_10862_11293# vssd1 0.63fF $ **FLOATING
C1238 a_11030_11039# vssd1 0.58fF $ **FLOATING
C1239 a_10589_10927# vssd1 1.43fF $ **FLOATING
C1240 a_10423_10927# vssd1 1.81fF $ **FLOATING
C1241 a_4537_10927# vssd1 0.18fF $ **FLOATING
C1242 _0686_.X vssd1 3.47fF $ **FLOATING
C1243 _0686_.A vssd1 2.55fF $ **FLOATING
C1244 a_6001_11177# vssd1 0.24fF $ **FLOATING
C1245 a_9495_11249# vssd1 0.54fF $ **FLOATING
C1246 _0597_.A2_N vssd1 1.03fF $ **FLOATING
C1247 _0597_.A1_N vssd1 4.33fF $ **FLOATING
C1248 a_9284_10901# vssd1 0.82fF $ **FLOATING
C1249 _0699_.A0 vssd1 5.66fF $ **FLOATING
C1250 a_7801_11079# vssd1 0.77fF $ **FLOATING
C1251 a_7623_10901# vssd1 0.83fF $ **FLOATING
C1252 a_6653_10933# vssd1 0.66fF $ **FLOATING
C1253 _0707_.A1 vssd1 0.97fF $ **FLOATING
C1254 _0698_.B1 vssd1 3.96fF $ **FLOATING
C1255 a_4251_11249# vssd1 0.54fF $ **FLOATING
C1256 _0698_.A2_N vssd1 1.82fF $ **FLOATING
C1257 _0698_.A1_N vssd1 1.14fF $ **FLOATING
C1258 a_4040_10901# vssd1 0.82fF $ **FLOATING
C1259 a_27249_11471# vssd1 0.21fF $ **FLOATING
C1260 a_25593_11471# vssd1 0.21fF $ **FLOATING
C1261 _0619_.X vssd1 3.70fF $ **FLOATING
C1262 _0650_.X vssd1 2.77fF $ **FLOATING
C1263 a_22741_11471# vssd1 0.21fF $ **FLOATING
C1264 a_24025_11471# vssd1 0.23fF $ **FLOATING
C1265 _0505_.X vssd1 1.02fF $ **FLOATING
C1266 a_19697_11471# vssd1 0.21fF $ **FLOATING
C1267 a_19613_11471# vssd1 0.17fF $ **FLOATING
C1268 _0489_.X vssd1 1.85fF $ **FLOATING
C1269 a_15105_11471# vssd1 0.21fF $ **FLOATING
C1270 a_14195_11471# vssd1 0.39fF $ **FLOATING
C1271 a_18045_11471# vssd1 0.23fF $ **FLOATING
C1272 _0588_.X vssd1 3.07fF $ **FLOATING
C1273 a_12065_11471# vssd1 0.23fF $ **FLOATING
C1274 a_9857_11471# vssd1 0.23fF $ **FLOATING
C1275 a_4993_11471# vssd1 0.20fF $ **FLOATING
C1276 a_27167_11471# vssd1 0.80fF $ **FLOATING
C1277 _0619_.B1 vssd1 9.35fF $ **FLOATING
C1278 _0619_.B2 vssd1 2.12fF $ **FLOATING
C1279 a_25511_11471# vssd1 0.80fF $ **FLOATING
C1280 _0650_.A1 vssd1 4.86fF $ **FLOATING
C1281 a_24535_11471# vssd1 0.61fF $ **FLOATING
C1282 a_24703_11445# vssd1 0.82fF $ **FLOATING
C1283 a_24110_11471# vssd1 0.63fF $ **FLOATING
C1284 a_24278_11445# vssd1 0.58fF $ **FLOATING
C1285 a_23837_11477# vssd1 1.43fF $ **FLOATING
C1286 a_23671_11477# vssd1 1.81fF $ **FLOATING
C1287 _1015_.CLK vssd1 10.38fF $ **FLOATING
C1288 a_22659_11471# vssd1 0.80fF $ **FLOATING
C1289 _0505_.A2 vssd1 11.33fF $ **FLOATING
C1290 _0505_.A1 vssd1 6.29fF $ **FLOATING
C1291 a_21127_11809# vssd1 0.56fF $ **FLOATING
C1292 a_19531_11471# vssd1 0.97fF $ **FLOATING
C1293 _0489_.C1 vssd1 3.01fF $ **FLOATING
C1294 a_18555_11471# vssd1 0.61fF $ **FLOATING
C1295 a_18723_11445# vssd1 0.82fF $ **FLOATING
C1296 a_18130_11471# vssd1 0.63fF $ **FLOATING
C1297 a_18298_11445# vssd1 0.58fF $ **FLOATING
C1298 a_17857_11477# vssd1 1.43fF $ **FLOATING
C1299 _0897_.D vssd1 5.60fF $ **FLOATING
C1300 a_17691_11477# vssd1 1.81fF $ **FLOATING
C1301 a_16863_11479# vssd1 0.65fF $ **FLOATING
C1302 a_15023_11471# vssd1 0.80fF $ **FLOATING
C1303 a_12575_11471# vssd1 0.61fF $ **FLOATING
C1304 a_12743_11445# vssd1 0.82fF $ **FLOATING
C1305 a_12150_11471# vssd1 0.63fF $ **FLOATING
C1306 a_12318_11445# vssd1 0.58fF $ **FLOATING
C1307 a_11877_11477# vssd1 1.43fF $ **FLOATING
C1308 a_11711_11477# vssd1 1.81fF $ **FLOATING
C1309 a_10367_11471# vssd1 0.61fF $ **FLOATING
C1310 a_10535_11445# vssd1 0.82fF $ **FLOATING
C1311 a_9942_11471# vssd1 0.63fF $ **FLOATING
C1312 a_10110_11445# vssd1 0.58fF $ **FLOATING
C1313 a_9669_11477# vssd1 1.43fF $ **FLOATING
C1314 _0985_.D vssd1 5.32fF $ **FLOATING
C1315 a_9503_11477# vssd1 1.81fF $ **FLOATING
C1316 a_8325_11769# vssd1 0.61fF $ **FLOATING
C1317 _0567_.A1 vssd1 3.40fF $ **FLOATING
C1318 a_7896_11703# vssd1 0.59fF $ **FLOATING
C1319 a_6600_11587# vssd1 0.50fF $ **FLOATING
C1320 _0708_.B1 vssd1 1.08fF $ **FLOATING
C1321 _0708_.A2 vssd1 1.52fF $ **FLOATING
C1322 _0708_.A3 vssd1 2.16fF $ **FLOATING
C1323 a_4864_11445# vssd1 0.65fF $ **FLOATING
C1324 a_3799_11471# vssd1 1.20fF $ **FLOATING
C1325 _1014_.Q vssd1 5.11fF $ **FLOATING
C1326 a_27337_12015# vssd1 0.23fF $ **FLOATING
C1327 a_27847_12381# vssd1 0.61fF $ **FLOATING
C1328 a_28015_12283# vssd1 0.82fF $ **FLOATING
C1329 a_27422_12381# vssd1 0.63fF $ **FLOATING
C1330 a_27590_12127# vssd1 0.58fF $ **FLOATING
C1331 a_27149_12015# vssd1 1.43fF $ **FLOATING
C1332 a_26983_12015# vssd1 1.81fF $ **FLOATING
C1333 a_25497_12015# vssd1 0.23fF $ **FLOATING
C1334 a_26007_12381# vssd1 0.61fF $ **FLOATING
C1335 a_26175_12283# vssd1 0.82fF $ **FLOATING
C1336 a_25582_12381# vssd1 0.63fF $ **FLOATING
C1337 a_25750_12127# vssd1 0.58fF $ **FLOATING
C1338 a_25309_12015# vssd1 1.43fF $ **FLOATING
C1339 a_25143_12015# vssd1 1.81fF $ **FLOATING
C1340 _0659_.X vssd1 1.76fF $ **FLOATING
C1341 a_22365_12265# vssd1 0.21fF $ **FLOATING
C1342 a_22281_12265# vssd1 0.17fF $ **FLOATING
C1343 _0612_.X vssd1 3.40fF $ **FLOATING
C1344 _0894_.Q vssd1 6.84fF $ **FLOATING
C1345 a_17260_12265# vssd1 0.26fF $ **FLOATING
C1346 _0565_.X vssd1 5.41fF $ **FLOATING
C1347 _0588_.A1 vssd1 3.77fF $ **FLOATING
C1348 a_14641_12015# vssd1 0.23fF $ **FLOATING
C1349 a_23303_12015# vssd1 0.62fF $ **FLOATING
C1350 a_22199_12015# vssd1 0.97fF $ **FLOATING
C1351 a_21127_12043# vssd1 0.56fF $ **FLOATING
C1352 a_20299_12043# vssd1 0.56fF $ **FLOATING
C1353 a_19439_12015# vssd1 0.62fF $ **FLOATING
C1354 a_18001_12043# vssd1 0.71fF $ **FLOATING
C1355 _0565_.A1 vssd1 3.91fF $ **FLOATING
C1356 _0565_.B1 vssd1 7.65fF $ **FLOATING
C1357 a_16829_12161# vssd1 0.67fF $ **FLOATING
C1358 a_15151_12381# vssd1 0.61fF $ **FLOATING
C1359 a_15319_12283# vssd1 0.82fF $ **FLOATING
C1360 a_14726_12381# vssd1 0.63fF $ **FLOATING
C1361 a_14894_12127# vssd1 0.58fF $ **FLOATING
C1362 a_14453_12015# vssd1 1.43fF $ **FLOATING
C1363 _0897_.Q vssd1 5.37fF $ **FLOATING
C1364 a_14287_12015# vssd1 1.81fF $ **FLOATING
C1365 _0475_.X vssd1 7.53fF $ **FLOATING
C1366 _0513_.X vssd1 7.69fF $ **FLOATING
C1367 a_8393_12015# vssd1 0.17fF $ **FLOATING
C1368 a_6563_12015# vssd1 0.21fF $ **FLOATING
C1369 _0655_.X vssd1 4.29fF $ **FLOATING
C1370 _0711_.A vssd1 2.96fF $ **FLOATING
C1371 a_4985_12061# vssd1 0.43fF $ **FLOATING
C1372 _0711_.B vssd1 3.08fF $ **FLOATING
C1373 a_4255_12265# vssd1 0.25fF $ **FLOATING
C1374 a_2405_12015# vssd1 0.23fF $ **FLOATING
C1375 a_11815_12265# vssd1 0.64fF $ **FLOATING
C1376 a_9911_12061# vssd1 0.71fF $ **FLOATING
C1377 a_9791_12015# vssd1 0.77fF $ **FLOATING
C1378 a_9595_12015# vssd1 0.74fF $ **FLOATING
C1379 a_8175_11989# vssd1 0.55fF $ **FLOATING
C1380 a_6427_11989# vssd1 0.79fF $ **FLOATING
C1381 a_5091_12021# vssd1 0.67fF $ **FLOATING
C1382 a_4037_11989# vssd1 0.55fF $ **FLOATING
C1383 a_2228_12015# vssd1 0.50fF $ **FLOATING
C1384 a_2122_12015# vssd1 0.58fF $ **FLOATING
C1385 a_1945_12015# vssd1 0.50fF $ **FLOATING
C1386 a_1626_12015# vssd1 0.54fF $ **FLOATING
C1387 io_in[5] vssd1 1.41fF
C1388 _1001_.Q vssd1 8.04fF $ **FLOATING
C1389 a_24068_12559# vssd1 0.26fF $ **FLOATING
C1390 a_22457_12559# vssd1 0.21fF $ **FLOATING
C1391 a_22373_12559# vssd1 0.17fF $ **FLOATING
C1392 a_25129_12559# vssd1 0.23fF $ **FLOATING
C1393 _0585_.X vssd1 3.85fF $ **FLOATING
C1394 a_25639_12559# vssd1 0.61fF $ **FLOATING
C1395 a_25807_12533# vssd1 0.82fF $ **FLOATING
C1396 a_25214_12559# vssd1 0.63fF $ **FLOATING
C1397 a_25382_12533# vssd1 0.58fF $ **FLOATING
C1398 a_24941_12565# vssd1 1.43fF $ **FLOATING
C1399 a_24775_12565# vssd1 1.81fF $ **FLOATING
C1400 _0576_.B1 vssd1 1.80fF $ **FLOATING
C1401 _0576_.D1 vssd1 4.43fF $ **FLOATING
C1402 a_23637_12533# vssd1 0.67fF $ **FLOATING
C1403 a_22291_12559# vssd1 0.97fF $ **FLOATING
C1404 _0563_.B1 vssd1 6.61fF $ **FLOATING
C1405 _0563_.C1 vssd1 2.53fF $ **FLOATING
C1406 a_19439_12675# vssd1 0.70fF $ **FLOATING
C1407 _0576_.X vssd1 2.42fF $ **FLOATING
C1408 _0533_.X vssd1 10.50fF $ **FLOATING
C1409 a_15833_12559# vssd1 0.21fF $ **FLOATING
C1410 a_15749_12559# vssd1 0.17fF $ **FLOATING
C1411 _0644_.X vssd1 2.60fF $ **FLOATING
C1412 _0502_.X vssd1 10.13fF $ **FLOATING
C1413 a_18703_12567# vssd1 0.65fF $ **FLOATING
C1414 a_17783_12672# vssd1 0.62fF $ **FLOATING
C1415 a_16897_12897# vssd1 0.71fF $ **FLOATING
C1416 a_15667_12559# vssd1 0.97fF $ **FLOATING
C1417 _0644_.A2 vssd1 5.48fF $ **FLOATING
C1418 a_13735_12925# vssd1 0.89fF $ **FLOATING
C1419 a_12763_12879# vssd1 0.71fF $ **FLOATING
C1420 a_12643_12559# vssd1 0.77fF $ **FLOATING
C1421 a_12447_12559# vssd1 0.74fF $ **FLOATING
C1422 _0479_.Y vssd1 7.91fF $ **FLOATING
C1423 _0678_.Y vssd1 2.51fF $ **FLOATING
C1424 a_7663_12879# vssd1 0.18fF $ **FLOATING
C1425 _0685_.X vssd1 3.04fF $ **FLOATING
C1426 a_5639_12879# vssd1 0.18fF $ **FLOATING
C1427 a_4989_12879# vssd1 0.17fF $ **FLOATING
C1428 a_9043_12567# vssd1 0.65fF $ **FLOATING
C1429 _0438_.A vssd1 7.57fF $ **FLOATING
C1430 _0684_.A2 vssd1 2.81fF $ **FLOATING
C1431 _0684_.A1 vssd1 6.55fF $ **FLOATING
C1432 a_6651_12672# vssd1 0.62fF $ **FLOATING
C1433 _0685_.B vssd1 8.51fF $ **FLOATING
C1434 _0756_.A2 vssd1 2.78fF $ **FLOATING
C1435 a_4771_12791# vssd1 0.55fF $ **FLOATING
C1436 a_26877_13103# vssd1 0.23fF $ **FLOATING
C1437 a_27387_13469# vssd1 0.61fF $ **FLOATING
C1438 a_27555_13371# vssd1 0.82fF $ **FLOATING
C1439 a_26962_13469# vssd1 0.63fF $ **FLOATING
C1440 a_27130_13215# vssd1 0.58fF $ **FLOATING
C1441 a_26689_13103# vssd1 1.43fF $ **FLOATING
C1442 _1066_.D vssd1 5.01fF $ **FLOATING
C1443 a_26523_13103# vssd1 1.81fF $ **FLOATING
C1444 a_25037_13103# vssd1 0.23fF $ **FLOATING
C1445 a_25547_13469# vssd1 0.61fF $ **FLOATING
C1446 a_25715_13371# vssd1 0.82fF $ **FLOATING
C1447 a_25122_13469# vssd1 0.63fF $ **FLOATING
C1448 a_25290_13215# vssd1 0.58fF $ **FLOATING
C1449 a_24849_13103# vssd1 1.43fF $ **FLOATING
C1450 _1011_.D vssd1 5.48fF $ **FLOATING
C1451 a_24683_13103# vssd1 1.81fF $ **FLOATING
C1452 a_23792_13353# vssd1 0.26fF $ **FLOATING
C1453 _0572_.X vssd1 2.53fF $ **FLOATING
C1454 a_21357_13103# vssd1 0.23fF $ **FLOATING
C1455 _0572_.A2 vssd1 13.33fF $ **FLOATING
C1456 _0572_.A1 vssd1 4.18fF $ **FLOATING
C1457 _0572_.D1 vssd1 1.12fF $ **FLOATING
C1458 a_23361_13249# vssd1 0.67fF $ **FLOATING
C1459 a_21867_13469# vssd1 0.61fF $ **FLOATING
C1460 a_22035_13371# vssd1 0.82fF $ **FLOATING
C1461 a_21442_13469# vssd1 0.63fF $ **FLOATING
C1462 a_21610_13215# vssd1 0.58fF $ **FLOATING
C1463 a_21169_13103# vssd1 1.43fF $ **FLOATING
C1464 _0890_.D vssd1 6.04fF $ **FLOATING
C1465 a_21003_13103# vssd1 1.81fF $ **FLOATING
C1466 a_17720_13353# vssd1 0.26fF $ **FLOATING
C1467 _0605_.X vssd1 2.23fF $ **FLOATING
C1468 _0483_.X vssd1 11.24fF $ **FLOATING
C1469 _0599_.X vssd1 2.44fF $ **FLOATING
C1470 _0524_.X vssd1 15.69fF $ **FLOATING
C1471 a_4468_13103# vssd1 0.20fF $ **FLOATING
C1472 a_10693_13353# vssd1 0.24fF $ **FLOATING
C1473 a_9497_13353# vssd1 0.24fF $ **FLOATING
C1474 _0654_.Y vssd1 1.69fF $ **FLOATING
C1475 a_6833_13353# vssd1 0.20fF $ **FLOATING
C1476 a_5821_13353# vssd1 0.20fF $ **FLOATING
C1477 a_19439_13103# vssd1 1.20fF $ **FLOATING
C1478 _0605_.C1 vssd1 1.09fF $ **FLOATING
C1479 _0605_.D1 vssd1 5.28fF $ **FLOATING
C1480 a_17289_13249# vssd1 0.67fF $ **FLOATING
C1481 a_16127_13103# vssd1 0.62fF $ **FLOATING
C1482 a_15115_13103# vssd1 0.73fF $ **FLOATING
C1483 a_14287_13103# vssd1 0.62fF $ **FLOATING
C1484 a_11913_13336# vssd1 0.70fF $ **FLOATING
C1485 a_11435_13103# vssd1 0.79fF $ **FLOATING
C1486 a_11582_13077# vssd1 0.80fF $ **FLOATING
C1487 _0746_.A2 vssd1 5.75fF $ **FLOATING
C1488 _0466_.A vssd1 11.99fF $ **FLOATING
C1489 _0745_.A1 vssd1 6.91fF $ **FLOATING
C1490 _0745_.A3 vssd1 4.78fF $ **FLOATING
C1491 a_6704_13077# vssd1 0.65fF $ **FLOATING
C1492 _0713_.A1 vssd1 2.08fF $ **FLOATING
C1493 _0713_.A3 vssd1 1.95fF $ **FLOATING
C1494 a_5692_13077# vssd1 0.65fF $ **FLOATING
C1495 _0745_.A2 vssd1 7.76fF $ **FLOATING
C1496 _0776_.A2 vssd1 5.86fF $ **FLOATING
C1497 a_4035_13077# vssd1 0.74fF $ **FLOATING
C1498 a_26053_13647# vssd1 0.21fF $ **FLOATING
C1499 _0664_.X vssd1 3.36fF $ **FLOATING
C1500 a_24485_13647# vssd1 0.23fF $ **FLOATING
C1501 _0570_.X vssd1 0.80fF $ **FLOATING
C1502 _1026_.Q vssd1 6.07fF $ **FLOATING
C1503 a_18088_13647# vssd1 0.26fF $ **FLOATING
C1504 a_19149_13647# vssd1 0.23fF $ **FLOATING
C1505 _0609_.X vssd1 2.52fF $ **FLOATING
C1506 _0600_.X vssd1 3.59fF $ **FLOATING
C1507 _0494_.X vssd1 6.93fF $ **FLOATING
C1508 _0610_.X vssd1 2.49fF $ **FLOATING
C1509 a_12065_13647# vssd1 0.23fF $ **FLOATING
C1510 a_8205_13647# vssd1 0.21fF $ **FLOATING
C1511 a_4901_13647# vssd1 0.20fF $ **FLOATING
C1512 a_9949_13647# vssd1 0.23fF $ **FLOATING
C1513 a_5731_13967# vssd1 0.18fF $ **FLOATING
C1514 a_25971_13647# vssd1 0.80fF $ **FLOATING
C1515 _0664_.A2 vssd1 7.72fF $ **FLOATING
C1516 a_24995_13647# vssd1 0.61fF $ **FLOATING
C1517 a_25163_13621# vssd1 0.82fF $ **FLOATING
C1518 a_24570_13647# vssd1 0.63fF $ **FLOATING
C1519 a_24738_13621# vssd1 0.58fF $ **FLOATING
C1520 a_24297_13653# vssd1 1.43fF $ **FLOATING
C1521 _1046_.D vssd1 5.73fF $ **FLOATING
C1522 a_24131_13653# vssd1 1.81fF $ **FLOATING
C1523 a_23303_13760# vssd1 0.62fF $ **FLOATING
C1524 a_22015_13760# vssd1 0.62fF $ **FLOATING
C1525 a_20635_13655# vssd1 0.65fF $ **FLOATING
C1526 a_19659_13647# vssd1 0.61fF $ **FLOATING
C1527 a_19827_13621# vssd1 0.82fF $ **FLOATING
C1528 a_19234_13647# vssd1 0.63fF $ **FLOATING
C1529 a_19402_13621# vssd1 0.58fF $ **FLOATING
C1530 a_18961_13653# vssd1 1.43fF $ **FLOATING
C1531 a_18795_13653# vssd1 1.81fF $ **FLOATING
C1532 _0609_.C1 vssd1 2.80fF $ **FLOATING
C1533 a_17657_13621# vssd1 0.67fF $ **FLOATING
C1534 a_15943_13760# vssd1 0.62fF $ **FLOATING
C1535 a_14637_13647# vssd1 0.67fF $ **FLOATING
C1536 a_14471_13647# vssd1 0.64fF $ **FLOATING
C1537 a_13551_13760# vssd1 0.62fF $ **FLOATING
C1538 a_12575_13647# vssd1 0.61fF $ **FLOATING
C1539 a_12743_13621# vssd1 0.82fF $ **FLOATING
C1540 a_12150_13647# vssd1 0.63fF $ **FLOATING
C1541 a_12318_13621# vssd1 0.58fF $ **FLOATING
C1542 a_11877_13653# vssd1 1.43fF $ **FLOATING
C1543 _0917_.D vssd1 5.59fF $ **FLOATING
C1544 a_11711_13653# vssd1 1.81fF $ **FLOATING
C1545 _0917_.CLK vssd1 12.78fF $ **FLOATING
C1546 a_10459_13647# vssd1 0.61fF $ **FLOATING
C1547 a_10627_13621# vssd1 0.82fF $ **FLOATING
C1548 a_10034_13647# vssd1 0.63fF $ **FLOATING
C1549 a_10202_13621# vssd1 0.58fF $ **FLOATING
C1550 a_9761_13653# vssd1 1.43fF $ **FLOATING
C1551 a_9595_13653# vssd1 1.81fF $ **FLOATING
C1552 _0922_.CLK vssd1 12.16fF $ **FLOATING
C1553 a_8123_13647# vssd1 1.01fF $ **FLOATING
C1554 _0626_.B1 vssd1 6.63fF $ **FLOATING
C1555 _0626_.B2 vssd1 3.01fF $ **FLOATING
C1556 a_7111_13655# vssd1 0.65fF $ **FLOATING
C1557 _0780_.A1 vssd1 1.52fF $ **FLOATING
C1558 _0791_.A1 vssd1 2.90fF $ **FLOATING
C1559 _0791_.A2 vssd1 2.68fF $ **FLOATING
C1560 _0791_.A3 vssd1 3.20fF $ **FLOATING
C1561 a_4772_13621# vssd1 0.65fF $ **FLOATING
C1562 a_3523_13655# vssd1 0.65fF $ **FLOATING
C1563 _1013_.Q vssd1 3.37fF $ **FLOATING
C1564 a_27337_14191# vssd1 0.23fF $ **FLOATING
C1565 a_27847_14557# vssd1 0.61fF $ **FLOATING
C1566 a_28015_14459# vssd1 0.82fF $ **FLOATING
C1567 a_27422_14557# vssd1 0.63fF $ **FLOATING
C1568 a_27590_14303# vssd1 0.58fF $ **FLOATING
C1569 a_27149_14191# vssd1 1.43fF $ **FLOATING
C1570 a_26983_14191# vssd1 1.81fF $ **FLOATING
C1571 _0620_.X vssd1 4.02fF $ **FLOATING
C1572 a_25225_14441# vssd1 0.21fF $ **FLOATING
C1573 _0940_.Q vssd1 5.21fF $ **FLOATING
C1574 a_22737_14191# vssd1 0.23fF $ **FLOATING
C1575 a_25143_14441# vssd1 0.80fF $ **FLOATING
C1576 a_23247_14557# vssd1 0.61fF $ **FLOATING
C1577 a_23415_14459# vssd1 0.82fF $ **FLOATING
C1578 a_22822_14557# vssd1 0.63fF $ **FLOATING
C1579 a_22990_14303# vssd1 0.58fF $ **FLOATING
C1580 a_22549_14191# vssd1 1.43fF $ **FLOATING
C1581 a_22383_14191# vssd1 1.81fF $ **FLOATING
C1582 a_21495_14219# vssd1 0.56fF $ **FLOATING
C1583 a_19439_14191# vssd1 0.70fF $ **FLOATING
C1584 a_18611_14191# vssd1 0.65fF $ **FLOATING
C1585 a_17904_14441# vssd1 0.26fF $ **FLOATING
C1586 _0630_.X vssd1 3.97fF $ **FLOATING
C1587 a_15929_14191# vssd1 0.23fF $ **FLOATING
C1588 _0630_.A2 vssd1 11.92fF $ **FLOATING
C1589 _0630_.A1 vssd1 4.97fF $ **FLOATING
C1590 a_17473_14337# vssd1 0.67fF $ **FLOATING
C1591 a_16439_14557# vssd1 0.61fF $ **FLOATING
C1592 a_16607_14459# vssd1 0.82fF $ **FLOATING
C1593 a_16014_14557# vssd1 0.63fF $ **FLOATING
C1594 a_16182_14303# vssd1 0.58fF $ **FLOATING
C1595 a_15741_14191# vssd1 1.43fF $ **FLOATING
C1596 a_15575_14191# vssd1 1.81fF $ **FLOATING
C1597 a_7164_14191# vssd1 0.20fF $ **FLOATING
C1598 a_12625_14441# vssd1 0.24fF $ **FLOATING
C1599 a_11233_14441# vssd1 0.21fF $ **FLOATING
C1600 a_11149_14441# vssd1 0.17fF $ **FLOATING
C1601 a_9301_14441# vssd1 0.21fF $ **FLOATING
C1602 a_9217_14441# vssd1 0.17fF $ **FLOATING
C1603 a_8037_14441# vssd1 0.19fF $ **FLOATING
C1604 _0779_.X vssd1 1.15fF $ **FLOATING
C1605 a_5737_14441# vssd1 0.19fF $ **FLOATING
C1606 a_14453_14557# vssd1 0.85fF $ **FLOATING
C1607 a_14287_14557# vssd1 0.60fF $ **FLOATING
C1608 a_11067_14191# vssd1 0.97fF $ **FLOATING
C1609 _0747_.B1 vssd1 3.13fF $ **FLOATING
C1610 _0747_.B2 vssd1 1.82fF $ **FLOATING
C1611 _0714_.B1 vssd1 1.64fF $ **FLOATING
C1612 _0714_.B2 vssd1 2.52fF $ **FLOATING
C1613 _0768_.C1 vssd1 2.29fF $ **FLOATING
C1614 _0768_.B1 vssd1 2.98fF $ **FLOATING
C1615 _0768_.A2 vssd1 2.29fF $ **FLOATING
C1616 a_7900_14165# vssd1 0.85fF $ **FLOATING
C1617 a_6938_14237# vssd1 0.44fF $ **FLOATING
C1618 a_6795_14343# vssd1 0.65fF $ **FLOATING
C1619 _0734_.C1 vssd1 1.80fF $ **FLOATING
C1620 _0768_.A1 vssd1 8.64fF $ **FLOATING
C1621 _0734_.A2 vssd1 6.23fF $ **FLOATING
C1622 a_5600_14165# vssd1 0.85fF $ **FLOATING
C1623 a_4165_14455# vssd1 0.60fF $ **FLOATING
C1624 a_4065_14237# vssd1 0.49fF $ **FLOATING
C1625 a_2879_14191# vssd1 0.73fF $ **FLOATING
C1626 a_3028_14165# vssd1 0.72fF $ **FLOATING
C1627 a_1591_14191# vssd1 0.65fF $ **FLOATING
C1628 io_in[6] vssd1 1.38fF
C1629 _0967_.Q vssd1 9.35fF $ **FLOATING
C1630 a_23745_14735# vssd1 0.21fF $ **FLOATING
C1631 a_23661_14735# vssd1 0.17fF $ **FLOATING
C1632 a_25589_14735# vssd1 0.23fF $ **FLOATING
C1633 _0663_.X vssd1 3.78fF $ **FLOATING
C1634 _0569_.X vssd1 1.69fF $ **FLOATING
C1635 _1025_.Q vssd1 4.36fF $ **FLOATING
C1636 a_20161_14735# vssd1 0.23fF $ **FLOATING
C1637 _0487_.X vssd1 14.16fF $ **FLOATING
C1638 _0606_.X vssd1 1.43fF $ **FLOATING
C1639 a_10313_14735# vssd1 0.21fF $ **FLOATING
C1640 a_10229_14735# vssd1 0.17fF $ **FLOATING
C1641 a_9497_14735# vssd1 0.24fF $ **FLOATING
C1642 a_8763_14735# vssd1 0.25fF $ **FLOATING
C1643 a_7843_14735# vssd1 0.25fF $ **FLOATING
C1644 a_6741_14735# vssd1 0.20fF $ **FLOATING
C1645 a_15101_14735# vssd1 0.23fF $ **FLOATING
C1646 _0546_.X vssd1 3.96fF $ **FLOATING
C1647 a_26099_14735# vssd1 0.61fF $ **FLOATING
C1648 a_26267_14709# vssd1 0.82fF $ **FLOATING
C1649 a_25674_14735# vssd1 0.63fF $ **FLOATING
C1650 a_25842_14709# vssd1 0.58fF $ **FLOATING
C1651 a_25401_14741# vssd1 1.43fF $ **FLOATING
C1652 a_25235_14741# vssd1 1.81fF $ **FLOATING
C1653 a_23579_14735# vssd1 0.97fF $ **FLOATING
C1654 a_22383_14848# vssd1 0.62fF $ **FLOATING
C1655 a_20671_14735# vssd1 0.61fF $ **FLOATING
C1656 a_20839_14709# vssd1 0.82fF $ **FLOATING
C1657 a_20246_14735# vssd1 0.63fF $ **FLOATING
C1658 a_20414_14709# vssd1 0.58fF $ **FLOATING
C1659 a_19973_14741# vssd1 1.43fF $ **FLOATING
C1660 a_19807_14741# vssd1 1.81fF $ **FLOATING
C1661 a_18611_14735# vssd1 1.20fF $ **FLOATING
C1662 a_17725_15073# vssd1 0.71fF $ **FLOATING
C1663 a_16863_14848# vssd1 0.62fF $ **FLOATING
C1664 a_15611_14735# vssd1 0.61fF $ **FLOATING
C1665 a_15779_14709# vssd1 0.82fF $ **FLOATING
C1666 a_15186_14735# vssd1 0.63fF $ **FLOATING
C1667 a_15354_14709# vssd1 0.58fF $ **FLOATING
C1668 a_14913_14741# vssd1 1.43fF $ **FLOATING
C1669 _0924_.D vssd1 4.92fF $ **FLOATING
C1670 a_14747_14741# vssd1 1.81fF $ **FLOATING
C1671 a_10147_14735# vssd1 0.97fF $ **FLOATING
C1672 _0770_.B1 vssd1 1.92fF $ **FLOATING
C1673 _0770_.B2 vssd1 0.90fF $ **FLOATING
C1674 _0546_.A2 vssd1 2.92fF $ **FLOATING
C1675 _0546_.B1 vssd1 3.41fF $ **FLOATING
C1676 a_8545_14709# vssd1 0.55fF $ **FLOATING
C1677 a_7625_14709# vssd1 0.55fF $ **FLOATING
C1678 _0793_.X vssd1 0.76fF $ **FLOATING
C1679 _0794_.A2 vssd1 1.93fF $ **FLOATING
C1680 _0794_.A3 vssd1 2.21fF $ **FLOATING
C1681 a_6612_14709# vssd1 0.65fF $ **FLOATING
C1682 a_5089_14851# vssd1 0.66fF $ **FLOATING
C1683 _0464_.X vssd1 1.53fF $ **FLOATING
C1684 a_2962_14735# vssd1 4.03fF $ **FLOATING
C1685 io_in[0] vssd1 7.45fF
C1686 a_2051_14848# vssd1 0.62fF $ **FLOATING
C1687 _0893_.Q vssd1 4.46fF $ **FLOATING
C1688 a_27337_15279# vssd1 0.23fF $ **FLOATING
C1689 a_27847_15645# vssd1 0.61fF $ **FLOATING
C1690 a_28015_15547# vssd1 0.82fF $ **FLOATING
C1691 a_27422_15645# vssd1 0.63fF $ **FLOATING
C1692 a_27590_15391# vssd1 0.58fF $ **FLOATING
C1693 a_27149_15279# vssd1 1.43fF $ **FLOATING
C1694 a_26983_15279# vssd1 1.81fF $ **FLOATING
C1695 a_24945_15279# vssd1 0.23fF $ **FLOATING
C1696 a_25455_15645# vssd1 0.61fF $ **FLOATING
C1697 a_25623_15547# vssd1 0.82fF $ **FLOATING
C1698 a_25030_15645# vssd1 0.63fF $ **FLOATING
C1699 a_25198_15391# vssd1 0.58fF $ **FLOATING
C1700 a_24757_15279# vssd1 1.43fF $ **FLOATING
C1701 _0891_.D vssd1 3.35fF $ **FLOATING
C1702 a_24591_15279# vssd1 1.81fF $ **FLOATING
C1703 _0893_.CLK vssd1 10.40fF $ **FLOATING
C1704 a_22606_15529# vssd1 0.33fF $ **FLOATING
C1705 a_21502_15529# vssd1 0.33fF $ **FLOATING
C1706 _0542_.X vssd1 7.53fF $ **FLOATING
C1707 a_19793_15279# vssd1 0.23fF $ **FLOATING
C1708 a_23487_15279# vssd1 0.70fF $ **FLOATING
C1709 fanout27.A vssd1 15.76fF $ **FLOATING
C1710 a_22449_15253# vssd1 0.72fF $ **FLOATING
C1711 a_21345_15253# vssd1 0.72fF $ **FLOATING
C1712 a_20303_15645# vssd1 0.61fF $ **FLOATING
C1713 a_20471_15547# vssd1 0.82fF $ **FLOATING
C1714 a_19878_15645# vssd1 0.63fF $ **FLOATING
C1715 a_20046_15391# vssd1 0.58fF $ **FLOATING
C1716 a_19605_15279# vssd1 1.43fF $ **FLOATING
C1717 _0962_.D vssd1 5.12fF $ **FLOATING
C1718 a_19439_15279# vssd1 1.81fF $ **FLOATING
C1719 _0523_.X vssd1 5.63fF $ **FLOATING
C1720 a_17857_15529# vssd1 0.21fF $ **FLOATING
C1721 a_17773_15529# vssd1 0.17fF $ **FLOATING
C1722 a_16984_15529# vssd1 0.26fF $ **FLOATING
C1723 _0580_.X vssd1 3.02fF $ **FLOATING
C1724 _0527_.X vssd1 9.33fF $ **FLOATING
C1725 a_11697_15279# vssd1 0.23fF $ **FLOATING
C1726 a_17691_15279# vssd1 0.97fF $ **FLOATING
C1727 _0523_.B1 vssd1 10.59fF $ **FLOATING
C1728 _0580_.A1 vssd1 5.45fF $ **FLOATING
C1729 _0580_.C1 vssd1 1.65fF $ **FLOATING
C1730 a_16553_15425# vssd1 0.67fF $ **FLOATING
C1731 a_15607_15307# vssd1 0.56fF $ **FLOATING
C1732 a_14603_15325# vssd1 0.71fF $ **FLOATING
C1733 a_14483_15279# vssd1 0.77fF $ **FLOATING
C1734 a_14287_15279# vssd1 0.74fF $ **FLOATING
C1735 a_12207_15645# vssd1 0.61fF $ **FLOATING
C1736 a_12375_15547# vssd1 0.82fF $ **FLOATING
C1737 a_11782_15645# vssd1 0.63fF $ **FLOATING
C1738 a_11950_15391# vssd1 0.58fF $ **FLOATING
C1739 a_11509_15279# vssd1 1.43fF $ **FLOATING
C1740 a_11343_15279# vssd1 1.81fF $ **FLOATING
C1741 _0474_.X vssd1 5.16fF $ **FLOATING
C1742 a_5455_15279# vssd1 0.18fF $ **FLOATING
C1743 a_10147_15529# vssd1 0.86fF $ **FLOATING
C1744 a_9411_15279# vssd1 0.65fF $ **FLOATING
C1745 a_7829_15529# vssd1 0.21fF $ **FLOATING
C1746 a_7745_15529# vssd1 0.17fF $ **FLOATING
C1747 a_6473_15529# vssd1 0.19fF $ **FLOATING
C1748 _0778_.Y vssd1 1.39fF $ **FLOATING
C1749 a_7663_15279# vssd1 0.97fF $ **FLOATING
C1750 _0760_.B1 vssd1 1.26fF $ **FLOATING
C1751 _0760_.B2 vssd1 3.12fF $ **FLOATING
C1752 _0758_.B1 vssd1 2.24fF $ **FLOATING
C1753 _0758_.A2 vssd1 1.88fF $ **FLOATING
C1754 a_6336_15253# vssd1 0.85fF $ **FLOATING
C1755 _0778_.B1 vssd1 2.61fF $ **FLOATING
C1756 _0778_.A2 vssd1 8.95fF $ **FLOATING
C1757 _0758_.A1 vssd1 6.95fF $ **FLOATING
C1758 a_3983_15279# vssd1 0.62fF $ **FLOATING
C1759 a_2693_15543# vssd1 0.60fF $ **FLOATING
C1760 a_2593_15325# vssd1 0.49fF $ **FLOATING
C1761 a_1775_15279# vssd1 0.65fF $ **FLOATING
C1762 _0715_.X vssd1 1.22fF $ **FLOATING
C1763 _0893_.D vssd1 4.74fF $ **FLOATING
C1764 a_25589_15823# vssd1 0.23fF $ **FLOATING
C1765 a_22369_15823# vssd1 0.23fF $ **FLOATING
C1766 _0627_.X vssd1 2.68fF $ **FLOATING
C1767 _0608_.X vssd1 2.80fF $ **FLOATING
C1768 a_19202_15823# vssd1 0.33fF $ **FLOATING
C1769 _0658_.X vssd1 3.49fF $ **FLOATING
C1770 _0628_.X vssd1 1.97fF $ **FLOATING
C1771 a_14559_15823# vssd1 0.25fF $ **FLOATING
C1772 _0921_.Q vssd1 6.71fF $ **FLOATING
C1773 a_10594_15823# vssd1 0.36fF $ **FLOATING
C1774 a_10397_15823# vssd1 0.25fF $ **FLOATING
C1775 a_10147_15823# vssd1 0.39fF $ **FLOATING
C1776 a_12801_15823# vssd1 0.23fF $ **FLOATING
C1777 _0529_.Y vssd1 9.40fF $ **FLOATING
C1778 a_9436_16143# vssd1 0.20fF $ **FLOATING
C1779 _0636_.X vssd1 5.35fF $ **FLOATING
C1780 a_6725_15823# vssd1 0.21fF $ **FLOATING
C1781 a_6641_15823# vssd1 0.17fF $ **FLOATING
C1782 a_5001_15823# vssd1 0.19fF $ **FLOATING
C1783 a_26099_15823# vssd1 0.61fF $ **FLOATING
C1784 a_26267_15797# vssd1 0.82fF $ **FLOATING
C1785 a_25674_15823# vssd1 0.63fF $ **FLOATING
C1786 a_25842_15797# vssd1 0.58fF $ **FLOATING
C1787 a_25401_15829# vssd1 1.43fF $ **FLOATING
C1788 _0892_.D vssd1 4.35fF $ **FLOATING
C1789 a_25235_15829# vssd1 1.81fF $ **FLOATING
C1790 a_23855_15831# vssd1 0.65fF $ **FLOATING
C1791 a_22879_15823# vssd1 0.61fF $ **FLOATING
C1792 a_23047_15797# vssd1 0.82fF $ **FLOATING
C1793 a_22454_15823# vssd1 0.63fF $ **FLOATING
C1794 a_22622_15797# vssd1 0.58fF $ **FLOATING
C1795 a_22181_15829# vssd1 1.43fF $ **FLOATING
C1796 _0925_.D vssd1 5.10fF $ **FLOATING
C1797 a_22015_15829# vssd1 1.81fF $ **FLOATING
C1798 a_20911_15936# vssd1 0.62fF $ **FLOATING
C1799 a_20083_15936# vssd1 0.62fF $ **FLOATING
C1800 _0658_.B1 vssd1 7.49fF $ **FLOATING
C1801 a_19045_15797# vssd1 0.72fF $ **FLOATING
C1802 a_17539_16161# vssd1 0.56fF $ **FLOATING
C1803 a_15667_15936# vssd1 0.62fF $ **FLOATING
C1804 a_14341_15797# vssd1 0.55fF $ **FLOATING
C1805 a_13311_15823# vssd1 0.61fF $ **FLOATING
C1806 a_13479_15797# vssd1 0.82fF $ **FLOATING
C1807 a_12886_15823# vssd1 0.63fF $ **FLOATING
C1808 a_13054_15797# vssd1 0.58fF $ **FLOATING
C1809 a_12613_15829# vssd1 1.43fF $ **FLOATING
C1810 a_12447_15829# vssd1 1.81fF $ **FLOATING
C1811 a_10814_15797# vssd1 0.65fF $ **FLOATING
C1812 _0508_.Y vssd1 6.39fF $ **FLOATING
C1813 a_9003_15797# vssd1 0.74fF $ **FLOATING
C1814 a_8155_16161# vssd1 0.56fF $ **FLOATING
C1815 a_6559_15823# vssd1 0.97fF $ **FLOATING
C1816 _0736_.B1 vssd1 1.80fF $ **FLOATING
C1817 a_4864_15797# vssd1 0.85fF $ **FLOATING
C1818 a_2686_15823# vssd1 4.03fF $ **FLOATING
C1819 clkbuf_1_1__f_io_in[0].A vssd1 6.74fF $ **FLOATING
C1820 a_1867_15831# vssd1 0.65fF $ **FLOATING
C1821 _0460_.C vssd1 6.70fF $ **FLOATING
C1822 _1012_.Q vssd1 4.49fF $ **FLOATING
C1823 a_27337_16367# vssd1 0.23fF $ **FLOATING
C1824 a_27847_16733# vssd1 0.61fF $ **FLOATING
C1825 a_28015_16635# vssd1 0.82fF $ **FLOATING
C1826 a_27422_16733# vssd1 0.63fF $ **FLOATING
C1827 a_27590_16479# vssd1 0.58fF $ **FLOATING
C1828 a_27149_16367# vssd1 1.43fF $ **FLOATING
C1829 _1012_.D vssd1 2.82fF $ **FLOATING
C1830 a_26983_16367# vssd1 1.81fF $ **FLOATING
C1831 _0939_.Q vssd1 4.29fF $ **FLOATING
C1832 a_24945_16367# vssd1 0.23fF $ **FLOATING
C1833 a_25455_16733# vssd1 0.61fF $ **FLOATING
C1834 a_25623_16635# vssd1 0.82fF $ **FLOATING
C1835 a_25030_16733# vssd1 0.63fF $ **FLOATING
C1836 a_25198_16479# vssd1 0.58fF $ **FLOATING
C1837 a_24757_16367# vssd1 1.43fF $ **FLOATING
C1838 a_24591_16367# vssd1 1.81fF $ **FLOATING
C1839 _0648_.X vssd1 4.14fF $ **FLOATING
C1840 a_23385_16617# vssd1 0.21fF $ **FLOATING
C1841 _0643_.X vssd1 5.30fF $ **FLOATING
C1842 a_22373_16617# vssd1 0.21fF $ **FLOATING
C1843 _0564_.X vssd1 4.42fF $ **FLOATING
C1844 _0564_.D vssd1 3.12fF $ **FLOATING
C1845 _0564_.C vssd1 0.95fF $ **FLOATING
C1846 a_19697_16617# vssd1 0.21fF $ **FLOATING
C1847 a_19613_16617# vssd1 0.17fF $ **FLOATING
C1848 _0521_.A vssd1 16.85fF $ **FLOATING
C1849 a_11269_16367# vssd1 0.44fF $ **FLOATING
C1850 a_15377_16367# vssd1 0.23fF $ **FLOATING
C1851 a_23303_16617# vssd1 0.80fF $ **FLOATING
C1852 _0648_.B1 vssd1 7.35fF $ **FLOATING
C1853 a_22291_16617# vssd1 0.80fF $ **FLOATING
C1854 _0643_.B1 vssd1 12.45fF $ **FLOATING
C1855 a_20819_16617# vssd1 0.70fF $ **FLOATING
C1856 a_19531_16367# vssd1 0.97fF $ **FLOATING
C1857 _0648_.A2 vssd1 11.58fF $ **FLOATING
C1858 _0561_.C1 vssd1 2.30fF $ **FLOATING
C1859 a_17909_16395# vssd1 0.71fF $ **FLOATING
C1860 a_16897_16395# vssd1 0.71fF $ **FLOATING
C1861 a_15887_16733# vssd1 0.61fF $ **FLOATING
C1862 a_16055_16635# vssd1 0.82fF $ **FLOATING
C1863 a_15462_16733# vssd1 0.63fF $ **FLOATING
C1864 a_15630_16479# vssd1 0.58fF $ **FLOATING
C1865 a_15189_16367# vssd1 1.43fF $ **FLOATING
C1866 _0990_.D vssd1 4.13fF $ **FLOATING
C1867 a_15023_16367# vssd1 1.81fF $ **FLOATING
C1868 a_9497_16367# vssd1 0.21fF $ **FLOATING
C1869 a_11437_16617# vssd1 0.39fF $ **FLOATING
C1870 _0882_.Y vssd1 11.15fF $ **FLOATING
C1871 _0880_.Y vssd1 8.81fF $ **FLOATING
C1872 _0882_.A2 vssd1 1.55fF $ **FLOATING
C1873 a_11068_16617# vssd1 0.63fF $ **FLOATING
C1874 _0880_.A1 vssd1 3.14fF $ **FLOATING
C1875 _0880_.A2 vssd1 2.50fF $ **FLOATING
C1876 a_9305_16672# vssd1 0.45fF $ **FLOATING
C1877 a_8393_16617# vssd1 0.24fF $ **FLOATING
C1878 _0735_.Y vssd1 1.51fF $ **FLOATING
C1879 _0735_.A2 vssd1 10.01fF $ **FLOATING
C1880 a_6467_16367# vssd1 0.65fF $ **FLOATING
C1881 _0461_.A vssd1 4.38fF $ **FLOATING
C1882 a_4621_16367# vssd1 0.21fF $ **FLOATING
C1883 _0877_.Y vssd1 5.89fF $ **FLOATING
C1884 a_5639_16367# vssd1 0.62fF $ **FLOATING
C1885 a_4429_16672# vssd1 0.45fF $ **FLOATING
C1886 a_3241_16617# vssd1 0.24fF $ **FLOATING
C1887 _0877_.A2 vssd1 1.20fF $ **FLOATING
C1888 a_1591_16367# vssd1 0.65fF $ **FLOATING
C1889 io_in[7] vssd1 1.43fF
C1890 _1000_.Q vssd1 4.95fF $ **FLOATING
C1891 a_25589_16911# vssd1 0.23fF $ **FLOATING
C1892 _1063_.Q vssd1 5.73fF $ **FLOATING
C1893 a_22369_16911# vssd1 0.23fF $ **FLOATING
C1894 a_20214_16911# vssd1 0.33fF $ **FLOATING
C1895 _0557_.X vssd1 3.94fF $ **FLOATING
C1896 _0602_.X vssd1 2.96fF $ **FLOATING
C1897 _0629_.X vssd1 2.04fF $ **FLOATING
C1898 a_12995_16911# vssd1 0.25fF $ **FLOATING
C1899 a_9305_16911# vssd1 0.23fF $ **FLOATING
C1900 a_7006_16911# vssd1 0.36fF $ **FLOATING
C1901 a_6809_16911# vssd1 0.25fF $ **FLOATING
C1902 a_6559_16911# vssd1 0.39fF $ **FLOATING
C1903 a_2599_16911# vssd1 0.25fF $ **FLOATING
C1904 _0518_.Y vssd1 8.66fF $ **FLOATING
C1905 a_26099_16911# vssd1 0.61fF $ **FLOATING
C1906 a_26267_16885# vssd1 0.82fF $ **FLOATING
C1907 a_25674_16911# vssd1 0.63fF $ **FLOATING
C1908 a_25842_16885# vssd1 0.58fF $ **FLOATING
C1909 a_25401_16917# vssd1 1.43fF $ **FLOATING
C1910 a_25235_16917# vssd1 1.81fF $ **FLOATING
C1911 a_22879_16911# vssd1 0.61fF $ **FLOATING
C1912 a_23047_16885# vssd1 0.82fF $ **FLOATING
C1913 a_22454_16911# vssd1 0.63fF $ **FLOATING
C1914 a_22622_16885# vssd1 0.58fF $ **FLOATING
C1915 a_22181_16917# vssd1 1.43fF $ **FLOATING
C1916 a_22015_16917# vssd1 1.81fF $ **FLOATING
C1917 a_21127_17249# vssd1 0.56fF $ **FLOATING
C1918 a_20057_16885# vssd1 0.72fF $ **FLOATING
C1919 a_18887_17024# vssd1 0.62fF $ **FLOATING
C1920 _0602_.A vssd1 18.80fF $ **FLOATING
C1921 a_18059_17024# vssd1 0.62fF $ **FLOATING
C1922 _0504_.A vssd1 18.35fF $ **FLOATING
C1923 a_14729_16911# vssd1 0.85fF $ **FLOATING
C1924 a_14563_16911# vssd1 0.60fF $ **FLOATING
C1925 a_12777_16885# vssd1 0.55fF $ **FLOATING
C1926 a_11936_17027# vssd1 0.50fF $ **FLOATING
C1927 a_10791_16919# vssd1 0.65fF $ **FLOATING
C1928 a_9815_16911# vssd1 0.61fF $ **FLOATING
C1929 a_9983_16885# vssd1 0.82fF $ **FLOATING
C1930 a_9390_16911# vssd1 0.63fF $ **FLOATING
C1931 a_9558_16885# vssd1 0.58fF $ **FLOATING
C1932 a_9117_16917# vssd1 1.43fF $ **FLOATING
C1933 _0986_.D vssd1 6.70fF $ **FLOATING
C1934 a_8951_16917# vssd1 1.81fF $ **FLOATING
C1935 a_8031_16911# vssd1 1.20fF $ **FLOATING
C1936 a_7226_16885# vssd1 0.65fF $ **FLOATING
C1937 a_5547_17027# vssd1 0.70fF $ **FLOATING
C1938 _0439_.A vssd1 8.93fF $ **FLOATING
C1939 a_3435_17231# vssd1 0.27fF $ **FLOATING
C1940 _0875_.X vssd1 4.16fF $ **FLOATING
C1941 a_4300_17027# vssd1 0.50fF $ **FLOATING
C1942 a_3298_17143# vssd1 0.60fF $ **FLOATING
C1943 _0874_.X vssd1 1.40fF $ **FLOATING
C1944 a_2381_16885# vssd1 0.55fF $ **FLOATING
C1945 a_27337_17455# vssd1 0.23fF $ **FLOATING
C1946 a_27847_17821# vssd1 0.61fF $ **FLOATING
C1947 a_28015_17723# vssd1 0.82fF $ **FLOATING
C1948 a_27422_17821# vssd1 0.63fF $ **FLOATING
C1949 a_27590_17567# vssd1 0.58fF $ **FLOATING
C1950 a_27149_17455# vssd1 1.43fF $ **FLOATING
C1951 a_26983_17455# vssd1 1.81fF $ **FLOATING
C1952 _0927_.D vssd1 3.68fF $ **FLOATING
C1953 a_25405_17455# vssd1 0.23fF $ **FLOATING
C1954 a_25915_17821# vssd1 0.61fF $ **FLOATING
C1955 a_26083_17723# vssd1 0.82fF $ **FLOATING
C1956 a_25490_17821# vssd1 0.63fF $ **FLOATING
C1957 a_25658_17567# vssd1 0.58fF $ **FLOATING
C1958 a_25217_17455# vssd1 1.43fF $ **FLOATING
C1959 _0926_.D vssd1 4.74fF $ **FLOATING
C1960 a_25051_17455# vssd1 1.81fF $ **FLOATING
C1961 _0574_.X vssd1 3.37fF $ **FLOATING
C1962 _0938_.Q vssd1 5.72fF $ **FLOATING
C1963 a_19793_17455# vssd1 0.23fF $ **FLOATING
C1964 a_22751_17455# vssd1 0.62fF $ **FLOATING
C1965 a_20303_17821# vssd1 0.61fF $ **FLOATING
C1966 a_20471_17723# vssd1 0.82fF $ **FLOATING
C1967 a_19878_17821# vssd1 0.63fF $ **FLOATING
C1968 a_20046_17567# vssd1 0.58fF $ **FLOATING
C1969 a_19605_17455# vssd1 1.43fF $ **FLOATING
C1970 a_19439_17455# vssd1 1.81fF $ **FLOATING
C1971 a_17401_17455# vssd1 0.23fF $ **FLOATING
C1972 a_17911_17821# vssd1 0.61fF $ **FLOATING
C1973 a_18079_17723# vssd1 0.82fF $ **FLOATING
C1974 a_17486_17821# vssd1 0.63fF $ **FLOATING
C1975 a_17654_17567# vssd1 0.58fF $ **FLOATING
C1976 a_17213_17455# vssd1 1.43fF $ **FLOATING
C1977 _1059_.D vssd1 5.52fF $ **FLOATING
C1978 a_17047_17455# vssd1 1.81fF $ **FLOATING
C1979 a_14559_17705# vssd1 0.25fF $ **FLOATING
C1980 a_12441_17705# vssd1 0.24fF $ **FLOATING
C1981 _0574_.C vssd1 9.83fF $ **FLOATING
C1982 a_11238_17705# vssd1 0.36fF $ **FLOATING
C1983 a_11041_17705# vssd1 0.25fF $ **FLOATING
C1984 a_10791_17705# vssd1 0.39fF $ **FLOATING
C1985 a_14341_17429# vssd1 0.55fF $ **FLOATING
C1986 a_13257_17821# vssd1 0.67fF $ **FLOATING
C1987 a_13091_17455# vssd1 0.64fF $ **FLOATING
C1988 a_11458_17429# vssd1 0.65fF $ **FLOATING
C1989 a_9963_17455# vssd1 0.65fF $ **FLOATING
C1990 a_9227_17455# vssd1 0.70fF $ **FLOATING
C1991 fanout37.A vssd1 18.39fF $ **FLOATING
C1992 a_8307_17455# vssd1 0.65fF $ **FLOATING
C1993 a_7393_17705# vssd1 0.19fF $ **FLOATING
C1994 a_6553_17705# vssd1 0.24fF $ **FLOATING
C1995 _0717_.B1 vssd1 3.03fF $ **FLOATING
C1996 a_7256_17429# vssd1 0.85fF $ **FLOATING
C1997 _0717_.A2 vssd1 9.71fF $ **FLOATING
C1998 a_5549_17719# vssd1 0.76fF $ **FLOATING
C1999 a_2869_17501# vssd1 0.43fF $ **FLOATING
C2000 a_3983_17455# vssd1 0.79fF $ **FLOATING
C2001 a_4132_17429# vssd1 1.17fF $ **FLOATING
C2002 a_2975_17461# vssd1 0.67fF $ **FLOATING
C2003 a_24949_17999# vssd1 0.21fF $ **FLOATING
C2004 _0558_.X vssd1 3.20fF $ **FLOATING
C2005 a_23381_17999# vssd1 0.23fF $ **FLOATING
C2006 a_18225_17999# vssd1 0.21fF $ **FLOATING
C2007 a_18141_17999# vssd1 0.17fF $ **FLOATING
C2008 a_17086_17999# vssd1 0.33fF $ **FLOATING
C2009 _0512_.A vssd1 17.02fF $ **FLOATING
C2010 _0668_.X vssd1 5.83fF $ **FLOATING
C2011 _0522_.X vssd1 1.99fF $ **FLOATING
C2012 _1057_.Q vssd1 5.50fF $ **FLOATING
C2013 a_10497_17999# vssd1 0.21fF $ **FLOATING
C2014 a_10413_17999# vssd1 0.17fF $ **FLOATING
C2015 a_7477_17999# vssd1 0.20fF $ **FLOATING
C2016 a_14825_17999# vssd1 0.23fF $ **FLOATING
C2017 a_4589_17999# vssd1 0.39fF $ **FLOATING
C2018 a_4167_17999# vssd1 0.86fF $ **FLOATING
C2019 _0873_.Y vssd1 1.20fF $ **FLOATING
C2020 a_24867_17999# vssd1 0.80fF $ **FLOATING
C2021 _0558_.A2 vssd1 7.39fF $ **FLOATING
C2022 a_23891_17999# vssd1 0.61fF $ **FLOATING
C2023 a_24059_17973# vssd1 0.82fF $ **FLOATING
C2024 a_23466_17999# vssd1 0.63fF $ **FLOATING
C2025 a_23634_17973# vssd1 0.58fF $ **FLOATING
C2026 a_23193_18005# vssd1 1.43fF $ **FLOATING
C2027 a_23027_18005# vssd1 1.81fF $ **FLOATING
C2028 _0964_.CLK vssd1 11.56fF $ **FLOATING
C2029 a_22015_18112# vssd1 0.62fF $ **FLOATING
C2030 _0582_.C vssd1 14.89fF $ **FLOATING
C2031 _0582_.A vssd1 18.39fF $ **FLOATING
C2032 a_19195_18337# vssd1 0.56fF $ **FLOATING
C2033 a_18059_17999# vssd1 0.97fF $ **FLOATING
C2034 _0512_.X vssd1 7.83fF $ **FLOATING
C2035 _0522_.B1 vssd1 11.68fF $ **FLOATING
C2036 a_16929_17973# vssd1 0.72fF $ **FLOATING
C2037 a_15335_17999# vssd1 0.61fF $ **FLOATING
C2038 a_15503_17973# vssd1 0.82fF $ **FLOATING
C2039 a_14910_17999# vssd1 0.63fF $ **FLOATING
C2040 a_15078_17973# vssd1 0.58fF $ **FLOATING
C2041 a_14637_18005# vssd1 1.43fF $ **FLOATING
C2042 a_14471_18005# vssd1 1.81fF $ **FLOATING
C2043 a_13367_17999# vssd1 0.70fF $ **FLOATING
C2044 a_10331_17999# vssd1 0.97fF $ **FLOATING
C2045 _0749_.A1 vssd1 1.41fF $ **FLOATING
C2046 _0749_.B1 vssd1 2.56fF $ **FLOATING
C2047 _0749_.B2 vssd1 2.53fF $ **FLOATING
C2048 a_8859_17999# vssd1 1.20fF $ **FLOATING
C2049 _0739_.B1 vssd1 3.09fF $ **FLOATING
C2050 _0739_.A2 vssd1 1.73fF $ **FLOATING
C2051 a_7348_17973# vssd1 0.65fF $ **FLOATING
C2052 _0472_.X vssd1 14.19fF $ **FLOATING
C2053 _0873_.A vssd1 8.54fF $ **FLOATING
C2054 _1068_.Q vssd1 5.64fF $ **FLOATING
C2055 a_26601_18543# vssd1 0.23fF $ **FLOATING
C2056 a_27111_18909# vssd1 0.61fF $ **FLOATING
C2057 a_27279_18811# vssd1 0.82fF $ **FLOATING
C2058 a_26686_18909# vssd1 0.63fF $ **FLOATING
C2059 a_26854_18655# vssd1 0.58fF $ **FLOATING
C2060 a_26413_18543# vssd1 1.43fF $ **FLOATING
C2061 a_26247_18543# vssd1 1.81fF $ **FLOATING
C2062 a_22974_18793# vssd1 0.33fF $ **FLOATING
C2063 _0662_.X vssd1 2.50fF $ **FLOATING
C2064 a_21265_18543# vssd1 0.23fF $ **FLOATING
C2065 _0662_.B1 vssd1 8.58fF $ **FLOATING
C2066 _0662_.A3 vssd1 16.89fF $ **FLOATING
C2067 a_22817_18517# vssd1 0.72fF $ **FLOATING
C2068 a_21775_18909# vssd1 0.61fF $ **FLOATING
C2069 a_21943_18811# vssd1 0.82fF $ **FLOATING
C2070 a_21350_18909# vssd1 0.63fF $ **FLOATING
C2071 a_21518_18655# vssd1 0.58fF $ **FLOATING
C2072 a_21077_18543# vssd1 1.43fF $ **FLOATING
C2073 _0991_.D vssd1 7.45fF $ **FLOATING
C2074 a_20911_18543# vssd1 1.81fF $ **FLOATING
C2075 a_20204_18793# vssd1 0.26fF $ **FLOATING
C2076 _0584_.X vssd1 3.40fF $ **FLOATING
C2077 a_18282_18793# vssd1 0.33fF $ **FLOATING
C2078 _0559_.X vssd1 2.82fF $ **FLOATING
C2079 _0577_.X vssd1 2.10fF $ **FLOATING
C2080 a_16258_18793# vssd1 0.33fF $ **FLOATING
C2081 _0667_.X vssd1 1.77fF $ **FLOATING
C2082 a_11697_18543# vssd1 0.23fF $ **FLOATING
C2083 _0584_.B1 vssd1 3.64fF $ **FLOATING
C2084 _0584_.C1 vssd1 1.84fF $ **FLOATING
C2085 a_19773_18689# vssd1 0.67fF $ **FLOATING
C2086 _0584_.A2 vssd1 4.81fF $ **FLOATING
C2087 a_18125_18517# vssd1 0.72fF $ **FLOATING
C2088 a_17139_18543# vssd1 0.62fF $ **FLOATING
C2089 _0667_.B1 vssd1 13.70fF $ **FLOATING
C2090 _0662_.A1 vssd1 19.48fF $ **FLOATING
C2091 a_16101_18517# vssd1 0.72fF $ **FLOATING
C2092 a_14603_18589# vssd1 0.71fF $ **FLOATING
C2093 a_14483_18543# vssd1 0.77fF $ **FLOATING
C2094 a_14287_18543# vssd1 0.74fF $ **FLOATING
C2095 a_12207_18909# vssd1 0.61fF $ **FLOATING
C2096 a_12375_18811# vssd1 0.82fF $ **FLOATING
C2097 a_11782_18909# vssd1 0.63fF $ **FLOATING
C2098 a_11950_18655# vssd1 0.58fF $ **FLOATING
C2099 a_11509_18543# vssd1 1.43fF $ **FLOATING
C2100 _0918_.D vssd1 5.54fF $ **FLOATING
C2101 a_11343_18543# vssd1 1.81fF $ **FLOATING
C2102 a_6929_18543# vssd1 0.19fF $ **FLOATING
C2103 _0577_.C vssd1 12.27fF $ **FLOATING
C2104 a_9407_18793# vssd1 0.25fF $ **FLOATING
C2105 a_8105_18793# vssd1 0.21fF $ **FLOATING
C2106 a_8021_18793# vssd1 0.17fF $ **FLOATING
C2107 a_6646_18865# vssd1 0.54fF $ **FLOATING
C2108 _0795_.A2_N vssd1 2.14fF $ **FLOATING
C2109 a_5819_18793# vssd1 0.25fF $ **FLOATING
C2110 _0511_.D vssd1 13.16fF $ **FLOATING
C2111 a_10533_18776# vssd1 0.70fF $ **FLOATING
C2112 a_10055_18543# vssd1 0.79fF $ **FLOATING
C2113 a_10202_18517# vssd1 0.80fF $ **FLOATING
C2114 a_9189_18517# vssd1 0.55fF $ **FLOATING
C2115 a_7939_18543# vssd1 0.97fF $ **FLOATING
C2116 _0719_.B2 vssd1 1.38fF $ **FLOATING
C2117 a_6516_18695# vssd1 0.64fF $ **FLOATING
C2118 _0795_.A1_N vssd1 2.70fF $ **FLOATING
C2119 _0783_.A1 vssd1 2.53fF $ **FLOATING
C2120 _0782_.X vssd1 2.04fF $ **FLOATING
C2121 a_5601_18517# vssd1 0.55fF $ **FLOATING
C2122 a_3983_18543# vssd1 0.62fF $ **FLOATING
C2123 _1067_.Q vssd1 4.41fF $ **FLOATING
C2124 a_25589_19087# vssd1 0.23fF $ **FLOATING
C2125 a_22737_19087# vssd1 0.23fF $ **FLOATING
C2126 _0583_.X vssd1 1.01fF $ **FLOATING
C2127 _0579_.X vssd1 2.57fF $ **FLOATING
C2128 _0937_.Q vssd1 4.88fF $ **FLOATING
C2129 a_12725_19087# vssd1 0.39fF $ **FLOATING
C2130 a_8305_19087# vssd1 0.20fF $ **FLOATING
C2131 a_6813_19087# vssd1 0.33fF $ **FLOATING
C2132 a_6559_19087# vssd1 0.38fF $ **FLOATING
C2133 a_14089_19087# vssd1 0.23fF $ **FLOATING
C2134 _0865_.Y vssd1 11.84fF $ **FLOATING
C2135 a_12557_19407# vssd1 0.44fF $ **FLOATING
C2136 a_10703_19407# vssd1 0.21fF $ **FLOATING
C2137 _0471_.X vssd1 14.32fF $ **FLOATING
C2138 a_5165_19087# vssd1 0.23fF $ **FLOATING
C2139 a_3333_19407# vssd1 0.21fF $ **FLOATING
C2140 _0872_.Y vssd1 6.94fF $ **FLOATING
C2141 a_26099_19087# vssd1 0.61fF $ **FLOATING
C2142 a_26267_19061# vssd1 0.82fF $ **FLOATING
C2143 a_25674_19087# vssd1 0.63fF $ **FLOATING
C2144 a_25842_19061# vssd1 0.58fF $ **FLOATING
C2145 a_25401_19093# vssd1 1.43fF $ **FLOATING
C2146 _1067_.D vssd1 5.80fF $ **FLOATING
C2147 a_25235_19093# vssd1 1.81fF $ **FLOATING
C2148 a_23247_19087# vssd1 0.61fF $ **FLOATING
C2149 a_23415_19061# vssd1 0.82fF $ **FLOATING
C2150 a_22822_19087# vssd1 0.63fF $ **FLOATING
C2151 a_22990_19061# vssd1 0.58fF $ **FLOATING
C2152 a_22549_19093# vssd1 1.43fF $ **FLOATING
C2153 _1016_.D vssd1 8.34fF $ **FLOATING
C2154 a_22383_19093# vssd1 1.81fF $ **FLOATING
C2155 a_20083_19200# vssd1 0.62fF $ **FLOATING
C2156 _0583_.C vssd1 6.21fF $ **FLOATING
C2157 a_17231_19200# vssd1 0.62fF $ **FLOATING
C2158 _0579_.C vssd1 5.46fF $ **FLOATING
C2159 _0583_.A vssd1 18.86fF $ **FLOATING
C2160 a_15575_19200# vssd1 0.62fF $ **FLOATING
C2161 a_14599_19087# vssd1 0.61fF $ **FLOATING
C2162 a_14767_19061# vssd1 0.82fF $ **FLOATING
C2163 a_14174_19087# vssd1 0.63fF $ **FLOATING
C2164 a_14342_19061# vssd1 0.58fF $ **FLOATING
C2165 a_13901_19093# vssd1 1.43fF $ **FLOATING
C2166 a_13735_19093# vssd1 1.81fF $ **FLOATING
C2167 a_12356_19203# vssd1 0.63fF $ **FLOATING
C2168 _0771_.C1 vssd1 2.58fF $ **FLOATING
C2169 a_10567_19061# vssd1 0.79fF $ **FLOATING
C2170 a_9503_19087# vssd1 1.20fF $ **FLOATING
C2171 _0763_.B1 vssd1 4.41fF $ **FLOATING
C2172 _0763_.A2 vssd1 2.09fF $ **FLOATING
C2173 a_8176_19061# vssd1 0.65fF $ **FLOATING
C2174 _0440_.C vssd1 1.99fF $ **FLOATING
C2175 a_4988_19087# vssd1 0.50fF $ **FLOATING
C2176 a_4882_19087# vssd1 0.58fF $ **FLOATING
C2177 a_4705_19087# vssd1 0.50fF $ **FLOATING
C2178 a_4386_19087# vssd1 0.54fF $ **FLOATING
C2179 _0872_.A1 vssd1 5.92fF $ **FLOATING
C2180 a_3141_19148# vssd1 0.45fF $ **FLOATING
C2181 a_25589_19631# vssd1 0.23fF $ **FLOATING
C2182 a_26099_19997# vssd1 0.61fF $ **FLOATING
C2183 a_26267_19899# vssd1 0.82fF $ **FLOATING
C2184 a_25674_19997# vssd1 0.63fF $ **FLOATING
C2185 a_25842_19743# vssd1 0.58fF $ **FLOATING
C2186 a_25401_19631# vssd1 1.43fF $ **FLOATING
C2187 _1047_.D vssd1 5.00fF $ **FLOATING
C2188 a_25235_19631# vssd1 1.81fF $ **FLOATING
C2189 a_22659_19631# vssd1 0.65fF $ **FLOATING
C2190 _1024_.Q vssd1 6.39fF $ **FLOATING
C2191 a_21173_19631# vssd1 0.23fF $ **FLOATING
C2192 a_21683_19997# vssd1 0.61fF $ **FLOATING
C2193 a_21851_19899# vssd1 0.82fF $ **FLOATING
C2194 a_21258_19997# vssd1 0.63fF $ **FLOATING
C2195 a_21426_19743# vssd1 0.58fF $ **FLOATING
C2196 a_20985_19631# vssd1 1.43fF $ **FLOATING
C2197 a_20819_19631# vssd1 1.81fF $ **FLOATING
C2198 a_17125_19631# vssd1 0.23fF $ **FLOATING
C2199 a_17635_19997# vssd1 0.61fF $ **FLOATING
C2200 a_17803_19899# vssd1 0.82fF $ **FLOATING
C2201 a_17210_19997# vssd1 0.63fF $ **FLOATING
C2202 a_17378_19743# vssd1 0.58fF $ **FLOATING
C2203 a_16937_19631# vssd1 1.43fF $ **FLOATING
C2204 a_16771_19631# vssd1 1.81fF $ **FLOATING
C2205 a_9769_19881# vssd1 0.21fF $ **FLOATING
C2206 _0807_.C vssd1 5.26fF $ **FLOATING
C2207 _0807_.A vssd1 12.35fF $ **FLOATING
C2208 _0807_.B vssd1 15.14fF $ **FLOATING
C2209 _0456_.A vssd1 8.54fF $ **FLOATING
C2210 _0456_.B vssd1 9.87fF $ **FLOATING
C2211 _0805_.A vssd1 1.33fF $ **FLOATING
C2212 _0872_.A2 vssd1 1.19fF $ **FLOATING
C2213 a_11067_19631# vssd1 0.89fF $ **FLOATING
C2214 a_9687_19881# vssd1 0.80fF $ **FLOATING
C2215 _0751_.B1 vssd1 1.66fF $ **FLOATING
C2216 _0751_.B2 vssd1 2.83fF $ **FLOATING
C2217 a_7939_19631# vssd1 1.20fF $ **FLOATING
C2218 a_6559_19631# vssd1 0.62fF $ **FLOATING
C2219 a_5642_19637# vssd1 0.82fF $ **FLOATING
C2220 a_4843_19659# vssd1 0.56fF $ **FLOATING
C2221 _0440_.A vssd1 10.01fF $ **FLOATING
C2222 a_24209_20175# vssd1 0.23fF $ **FLOATING
C2223 _1023_.Q vssd1 4.70fF $ **FLOATING
C2224 a_22369_20175# vssd1 0.23fF $ **FLOATING
C2225 _1062_.Q vssd1 8.18fF $ **FLOATING
C2226 a_20345_20175# vssd1 0.23fF $ **FLOATING
C2227 _1050_.Q vssd1 5.48fF $ **FLOATING
C2228 a_16029_20175# vssd1 0.24fF $ **FLOATING
C2229 a_18505_20175# vssd1 0.23fF $ **FLOATING
C2230 a_11893_20175# vssd1 0.20fF $ **FLOATING
C2231 a_10977_20175# vssd1 0.19fF $ **FLOATING
C2232 a_14457_20175# vssd1 0.23fF $ **FLOATING
C2233 a_7291_20175# vssd1 0.25fF $ **FLOATING
C2234 a_5635_20175# vssd1 0.25fF $ **FLOATING
C2235 a_9313_20495# vssd1 0.17fF $ **FLOATING
C2236 _0459_.X vssd1 2.05fF $ **FLOATING
C2237 _0737_.X vssd1 2.03fF $ **FLOATING
C2238 a_24719_20175# vssd1 0.61fF $ **FLOATING
C2239 a_24887_20149# vssd1 0.82fF $ **FLOATING
C2240 a_24294_20175# vssd1 0.63fF $ **FLOATING
C2241 a_24462_20149# vssd1 0.58fF $ **FLOATING
C2242 a_24021_20181# vssd1 1.43fF $ **FLOATING
C2243 _0965_.D vssd1 8.74fF $ **FLOATING
C2244 a_23855_20181# vssd1 1.81fF $ **FLOATING
C2245 a_22879_20175# vssd1 0.61fF $ **FLOATING
C2246 a_23047_20149# vssd1 0.82fF $ **FLOATING
C2247 a_22454_20175# vssd1 0.63fF $ **FLOATING
C2248 a_22622_20149# vssd1 0.58fF $ **FLOATING
C2249 a_22181_20181# vssd1 1.43fF $ **FLOATING
C2250 a_22015_20181# vssd1 1.81fF $ **FLOATING
C2251 a_20855_20175# vssd1 0.61fF $ **FLOATING
C2252 a_21023_20149# vssd1 0.82fF $ **FLOATING
C2253 a_20430_20175# vssd1 0.63fF $ **FLOATING
C2254 a_20598_20149# vssd1 0.58fF $ **FLOATING
C2255 a_20157_20181# vssd1 1.43fF $ **FLOATING
C2256 a_19991_20181# vssd1 1.81fF $ **FLOATING
C2257 _1062_.CLK vssd1 10.86fF $ **FLOATING
C2258 a_19015_20175# vssd1 0.61fF $ **FLOATING
C2259 a_19183_20149# vssd1 0.82fF $ **FLOATING
C2260 a_18590_20175# vssd1 0.63fF $ **FLOATING
C2261 a_18758_20149# vssd1 0.58fF $ **FLOATING
C2262 a_18317_20181# vssd1 1.43fF $ **FLOATING
C2263 a_18151_20181# vssd1 1.81fF $ **FLOATING
C2264 a_14967_20175# vssd1 0.61fF $ **FLOATING
C2265 a_15135_20149# vssd1 0.82fF $ **FLOATING
C2266 a_14542_20175# vssd1 0.63fF $ **FLOATING
C2267 a_14710_20149# vssd1 0.58fF $ **FLOATING
C2268 a_14269_20181# vssd1 1.43fF $ **FLOATING
C2269 _0919_.D vssd1 5.53fF $ **FLOATING
C2270 a_14103_20181# vssd1 1.81fF $ **FLOATING
C2271 a_11764_20149# vssd1 0.65fF $ **FLOATING
C2272 a_10714_20541# vssd1 0.59fF $ **FLOATING
C2273 _0773_.A2_N vssd1 3.14fF $ **FLOATING
C2274 _0773_.A1_N vssd1 1.12fF $ **FLOATING
C2275 a_10564_20407# vssd1 0.66fF $ **FLOATING
C2276 a_9095_20407# vssd1 0.55fF $ **FLOATING
C2277 a_8256_20291# vssd1 0.50fF $ **FLOATING
C2278 _0784_.A2 vssd1 2.14fF $ **FLOATING
C2279 _0784_.A1 vssd1 4.10fF $ **FLOATING
C2280 a_7073_20149# vssd1 0.55fF $ **FLOATING
C2281 _0812_.A2 vssd1 12.05fF $ **FLOATING
C2282 _0812_.B1 vssd1 2.89fF $ **FLOATING
C2283 a_5417_20149# vssd1 0.55fF $ **FLOATING
C2284 a_4170_20291# vssd1 0.82fF $ **FLOATING
C2285 _0722_.A vssd1 9.47fF $ **FLOATING
C2286 _0722_.B vssd1 9.68fF $ **FLOATING
C2287 _0722_.C vssd1 10.48fF $ **FLOATING
C2288 _0966_.Q vssd1 5.03fF $ **FLOATING
C2289 a_26417_20719# vssd1 0.23fF $ **FLOATING
C2290 a_26927_21085# vssd1 0.61fF $ **FLOATING
C2291 a_27095_20987# vssd1 0.82fF $ **FLOATING
C2292 a_26502_21085# vssd1 0.63fF $ **FLOATING
C2293 a_26670_20831# vssd1 0.58fF $ **FLOATING
C2294 a_26229_20719# vssd1 1.43fF $ **FLOATING
C2295 _0966_.D vssd1 4.07fF $ **FLOATING
C2296 a_26063_20719# vssd1 1.81fF $ **FLOATING
C2297 _0963_.Q vssd1 3.91fF $ **FLOATING
C2298 a_22829_20719# vssd1 0.23fF $ **FLOATING
C2299 a_23339_21085# vssd1 0.61fF $ **FLOATING
C2300 a_23507_20987# vssd1 0.82fF $ **FLOATING
C2301 a_22914_21085# vssd1 0.63fF $ **FLOATING
C2302 a_23082_20831# vssd1 0.58fF $ **FLOATING
C2303 a_22641_20719# vssd1 1.43fF $ **FLOATING
C2304 _0963_.D vssd1 5.11fF $ **FLOATING
C2305 a_22475_20719# vssd1 1.81fF $ **FLOATING
C2306 _1049_.Q vssd1 9.37fF $ **FLOATING
C2307 a_20989_20719# vssd1 0.23fF $ **FLOATING
C2308 a_21499_21085# vssd1 0.61fF $ **FLOATING
C2309 a_21667_20987# vssd1 0.82fF $ **FLOATING
C2310 a_21074_21085# vssd1 0.63fF $ **FLOATING
C2311 a_21242_20831# vssd1 0.58fF $ **FLOATING
C2312 a_20801_20719# vssd1 1.43fF $ **FLOATING
C2313 a_20635_20719# vssd1 1.81fF $ **FLOATING
C2314 _0920_.Q vssd1 6.67fF $ **FLOATING
C2315 a_15837_20719# vssd1 0.23fF $ **FLOATING
C2316 a_16347_21085# vssd1 0.61fF $ **FLOATING
C2317 a_16515_20987# vssd1 0.82fF $ **FLOATING
C2318 a_15922_21085# vssd1 0.63fF $ **FLOATING
C2319 a_16090_20831# vssd1 0.58fF $ **FLOATING
C2320 a_15649_20719# vssd1 1.43fF $ **FLOATING
C2321 _0920_.D vssd1 3.15fF $ **FLOATING
C2322 a_15483_20719# vssd1 1.81fF $ **FLOATING
C2323 _0801_.X vssd1 2.20fF $ **FLOATING
C2324 a_11697_20719# vssd1 0.23fF $ **FLOATING
C2325 a_14319_20747# vssd1 0.56fF $ **FLOATING
C2326 a_12207_21085# vssd1 0.61fF $ **FLOATING
C2327 a_12375_20987# vssd1 0.82fF $ **FLOATING
C2328 a_11782_21085# vssd1 0.63fF $ **FLOATING
C2329 a_11950_20831# vssd1 0.58fF $ **FLOATING
C2330 a_11509_20719# vssd1 1.43fF $ **FLOATING
C2331 _0987_.D vssd1 9.49fF $ **FLOATING
C2332 a_11343_20719# vssd1 1.81fF $ **FLOATING
C2333 _0761_.X vssd1 2.05fF $ **FLOATING
C2334 _0761_.B vssd1 5.80fF $ **FLOATING
C2335 a_7197_20969# vssd1 0.24fF $ **FLOATING
C2336 a_5173_20719# vssd1 0.21fF $ **FLOATING
C2337 _0870_.Y vssd1 8.90fF $ **FLOATING
C2338 a_9636_20969# vssd1 0.50fF $ **FLOATING
C2339 a_8123_20719# vssd1 1.20fF $ **FLOATING
C2340 _0808_.A vssd1 1.55fF $ **FLOATING
C2341 _0869_.B1 vssd1 10.97fF $ **FLOATING
C2342 a_6283_20719# vssd1 0.62fF $ **FLOATING
C2343 _0803_.X vssd1 2.79fF $ **FLOATING
C2344 _0869_.Y vssd1 1.43fF $ **FLOATING
C2345 a_4981_21024# vssd1 0.45fF $ **FLOATING
C2346 a_25589_21263# vssd1 0.23fF $ **FLOATING
C2347 _1048_.Q vssd1 5.50fF $ **FLOATING
C2348 a_23565_21263# vssd1 0.23fF $ **FLOATING
C2349 a_20437_21263# vssd1 0.23fF $ **FLOATING
C2350 a_15945_21263# vssd1 0.39fF $ **FLOATING
C2351 a_18597_21263# vssd1 0.23fF $ **FLOATING
C2352 _0863_.Y vssd1 15.55fF $ **FLOATING
C2353 a_15777_21583# vssd1 0.44fF $ **FLOATING
C2354 _0864_.Y vssd1 2.15fF $ **FLOATING
C2355 a_12525_21263# vssd1 0.23fF $ **FLOATING
C2356 _0988_.Q vssd1 7.18fF $ **FLOATING
C2357 a_9857_21263# vssd1 0.23fF $ **FLOATING
C2358 _0936_.Q vssd1 6.52fF $ **FLOATING
C2359 a_8017_21263# vssd1 0.23fF $ **FLOATING
C2360 a_26099_21263# vssd1 0.61fF $ **FLOATING
C2361 a_26267_21237# vssd1 0.82fF $ **FLOATING
C2362 a_25674_21263# vssd1 0.63fF $ **FLOATING
C2363 a_25842_21237# vssd1 0.58fF $ **FLOATING
C2364 a_25401_21269# vssd1 1.43fF $ **FLOATING
C2365 _0992_.D vssd1 6.99fF $ **FLOATING
C2366 a_25235_21269# vssd1 1.81fF $ **FLOATING
C2367 a_24075_21263# vssd1 0.61fF $ **FLOATING
C2368 a_24243_21237# vssd1 0.82fF $ **FLOATING
C2369 a_23650_21263# vssd1 0.63fF $ **FLOATING
C2370 a_23818_21237# vssd1 0.58fF $ **FLOATING
C2371 a_23377_21269# vssd1 1.43fF $ **FLOATING
C2372 _1048_.D vssd1 3.77fF $ **FLOATING
C2373 a_23211_21269# vssd1 1.81fF $ **FLOATING
C2374 a_20947_21263# vssd1 0.61fF $ **FLOATING
C2375 a_21115_21237# vssd1 0.82fF $ **FLOATING
C2376 a_20522_21263# vssd1 0.63fF $ **FLOATING
C2377 a_20690_21237# vssd1 0.58fF $ **FLOATING
C2378 a_20249_21269# vssd1 1.43fF $ **FLOATING
C2379 a_20083_21269# vssd1 1.81fF $ **FLOATING
C2380 _0931_.CLK vssd1 12.69fF $ **FLOATING
C2381 a_19107_21263# vssd1 0.61fF $ **FLOATING
C2382 a_19275_21237# vssd1 0.82fF $ **FLOATING
C2383 a_18682_21263# vssd1 0.63fF $ **FLOATING
C2384 a_18850_21237# vssd1 0.58fF $ **FLOATING
C2385 a_18409_21269# vssd1 1.43fF $ **FLOATING
C2386 _1060_.D vssd1 3.94fF $ **FLOATING
C2387 a_18243_21269# vssd1 1.81fF $ **FLOATING
C2388 _0863_.A2 vssd1 1.33fF $ **FLOATING
C2389 a_15576_21379# vssd1 0.63fF $ **FLOATING
C2390 _0863_.A1 vssd1 4.12fF $ **FLOATING
C2391 a_13035_21263# vssd1 0.61fF $ **FLOATING
C2392 a_13203_21237# vssd1 0.82fF $ **FLOATING
C2393 a_12610_21263# vssd1 0.63fF $ **FLOATING
C2394 a_12778_21237# vssd1 0.58fF $ **FLOATING
C2395 a_12337_21269# vssd1 1.43fF $ **FLOATING
C2396 a_12171_21269# vssd1 1.81fF $ **FLOATING
C2397 _0935_.CLK vssd1 13.65fF $ **FLOATING
C2398 a_10367_21263# vssd1 0.61fF $ **FLOATING
C2399 a_10535_21237# vssd1 0.82fF $ **FLOATING
C2400 a_9942_21263# vssd1 0.63fF $ **FLOATING
C2401 a_10110_21237# vssd1 0.58fF $ **FLOATING
C2402 a_9669_21269# vssd1 1.43fF $ **FLOATING
C2403 _0988_.D vssd1 5.61fF $ **FLOATING
C2404 a_9503_21269# vssd1 1.81fF $ **FLOATING
C2405 a_8527_21263# vssd1 0.61fF $ **FLOATING
C2406 a_8695_21237# vssd1 0.82fF $ **FLOATING
C2407 a_8102_21263# vssd1 0.63fF $ **FLOATING
C2408 a_8270_21237# vssd1 0.58fF $ **FLOATING
C2409 a_7829_21269# vssd1 1.43fF $ **FLOATING
C2410 _0935_.Q vssd1 6.05fF $ **FLOATING
C2411 a_7663_21269# vssd1 1.81fF $ **FLOATING
C2412 a_6876_21379# vssd1 0.50fF $ **FLOATING
C2413 a_3891_21263# vssd1 1.20fF $ **FLOATING
C2414 _0725_.A vssd1 1.84fF $ **FLOATING
C2415 a_3155_21271# vssd1 0.65fF $ **FLOATING
C2416 _0721_.A vssd1 2.22fF $ **FLOATING
C2417 _0999_.Q vssd1 5.74fF $ **FLOATING
C2418 a_27337_21807# vssd1 0.23fF $ **FLOATING
C2419 a_27847_22173# vssd1 0.61fF $ **FLOATING
C2420 a_28015_22075# vssd1 0.82fF $ **FLOATING
C2421 a_27422_22173# vssd1 0.63fF $ **FLOATING
C2422 a_27590_21919# vssd1 0.58fF $ **FLOATING
C2423 a_27149_21807# vssd1 1.43fF $ **FLOATING
C2424 a_26983_21807# vssd1 1.81fF $ **FLOATING
C2425 _0999_.CLK vssd1 11.42fF $ **FLOATING
C2426 _0930_.Q vssd1 6.05fF $ **FLOATING
C2427 a_24945_21807# vssd1 0.23fF $ **FLOATING
C2428 a_25455_22173# vssd1 0.61fF $ **FLOATING
C2429 a_25623_22075# vssd1 0.82fF $ **FLOATING
C2430 a_25030_22173# vssd1 0.63fF $ **FLOATING
C2431 a_25198_21919# vssd1 0.58fF $ **FLOATING
C2432 a_24757_21807# vssd1 1.43fF $ **FLOATING
C2433 a_24591_21807# vssd1 1.81fF $ **FLOATING
C2434 _1022_.Q vssd1 4.10fF $ **FLOATING
C2435 a_21909_21807# vssd1 0.23fF $ **FLOATING
C2436 a_22419_22173# vssd1 0.61fF $ **FLOATING
C2437 a_22587_22075# vssd1 0.82fF $ **FLOATING
C2438 a_21994_22173# vssd1 0.63fF $ **FLOATING
C2439 a_22162_21919# vssd1 0.58fF $ **FLOATING
C2440 a_21721_21807# vssd1 1.43fF $ **FLOATING
C2441 a_21555_21807# vssd1 1.81fF $ **FLOATING
C2442 _0934_.Q vssd1 5.92fF $ **FLOATING
C2443 a_16757_21807# vssd1 0.23fF $ **FLOATING
C2444 a_17267_22173# vssd1 0.61fF $ **FLOATING
C2445 a_17435_22075# vssd1 0.82fF $ **FLOATING
C2446 a_16842_22173# vssd1 0.63fF $ **FLOATING
C2447 a_17010_21919# vssd1 0.58fF $ **FLOATING
C2448 a_16569_21807# vssd1 1.43fF $ **FLOATING
C2449 a_16403_21807# vssd1 1.81fF $ **FLOATING
C2450 a_15667_21807# vssd1 0.65fF $ **FLOATING
C2451 a_12893_21807# vssd1 0.23fF $ **FLOATING
C2452 a_6287_21807# vssd1 0.21fF $ **FLOATING
C2453 a_1591_21807# vssd1 0.55fF $ **FLOATING
C2454 a_12716_21807# vssd1 0.50fF $ **FLOATING
C2455 a_12610_21807# vssd1 0.58fF $ **FLOATING
C2456 a_12433_21807# vssd1 0.50fF $ **FLOATING
C2457 _0849_.X vssd1 13.40fF $ **FLOATING
C2458 a_12114_21807# vssd1 0.54fF $ **FLOATING
C2459 a_10789_22071# vssd1 0.60fF $ **FLOATING
C2460 a_10689_21853# vssd1 0.49fF $ **FLOATING
C2461 a_5245_22057# vssd1 0.20fF $ **FLOATING
C2462 io_out[0] vssd1 4.15fF
C2463 a_2039_22057# vssd1 0.38fF $ **FLOATING
C2464 io_out[2] vssd1 1.50fF
C2465 a_1591_22057# vssd1 0.38fF $ **FLOATING
C2466 a_7244_22057# vssd1 0.50fF $ **FLOATING
C2467 _0797_.B1 vssd1 1.07fF $ **FLOATING
C2468 _0797_.A2 vssd1 1.82fF $ **FLOATING
C2469 _0797_.A1 vssd1 10.33fF $ **FLOATING
C2470 a_6151_21781# vssd1 0.79fF $ **FLOATING
C2471 _0727_.A1 vssd1 3.37fF $ **FLOATING
C2472 a_5047_21781# vssd1 0.80fF $ **FLOATING
C2473 _0753_.A2 vssd1 5.22fF $ **FLOATING
C2474 _0929_.Q vssd1 4.39fF $ **FLOATING
C2475 a_24209_22351# vssd1 0.23fF $ **FLOATING
C2476 a_22369_22351# vssd1 0.23fF $ **FLOATING
C2477 a_20345_22351# vssd1 0.23fF $ **FLOATING
C2478 a_11983_22351# vssd1 0.25fF $ **FLOATING
C2479 a_13261_22351# vssd1 0.23fF $ **FLOATING
C2480 _0858_.X vssd1 14.20fF $ **FLOATING
C2481 _1056_.Q vssd1 6.44fF $ **FLOATING
C2482 a_6831_22351# vssd1 0.25fF $ **FLOATING
C2483 a_10041_22351# vssd1 0.23fF $ **FLOATING
C2484 _0868_.X vssd1 10.72fF $ **FLOATING
C2485 a_24719_22351# vssd1 0.61fF $ **FLOATING
C2486 a_24887_22325# vssd1 0.82fF $ **FLOATING
C2487 a_24294_22351# vssd1 0.63fF $ **FLOATING
C2488 a_24462_22325# vssd1 0.58fF $ **FLOATING
C2489 a_24021_22357# vssd1 1.43fF $ **FLOATING
C2490 a_23855_22357# vssd1 1.81fF $ **FLOATING
C2491 a_22879_22351# vssd1 0.61fF $ **FLOATING
C2492 a_23047_22325# vssd1 0.82fF $ **FLOATING
C2493 a_22454_22351# vssd1 0.63fF $ **FLOATING
C2494 a_22622_22325# vssd1 0.58fF $ **FLOATING
C2495 a_22181_22357# vssd1 1.43fF $ **FLOATING
C2496 _1017_.D vssd1 5.11fF $ **FLOATING
C2497 a_22015_22357# vssd1 1.81fF $ **FLOATING
C2498 a_20855_22351# vssd1 0.61fF $ **FLOATING
C2499 a_21023_22325# vssd1 0.82fF $ **FLOATING
C2500 a_20430_22351# vssd1 0.63fF $ **FLOATING
C2501 a_20598_22325# vssd1 0.58fF $ **FLOATING
C2502 a_20157_22357# vssd1 1.43fF $ **FLOATING
C2503 _0932_.D vssd1 5.60fF $ **FLOATING
C2504 a_19991_22357# vssd1 1.81fF $ **FLOATING
C2505 a_13771_22351# vssd1 0.61fF $ **FLOATING
C2506 a_13939_22325# vssd1 0.82fF $ **FLOATING
C2507 a_13346_22351# vssd1 0.63fF $ **FLOATING
C2508 a_13514_22325# vssd1 0.58fF $ **FLOATING
C2509 a_13073_22357# vssd1 1.43fF $ **FLOATING
C2510 a_12907_22357# vssd1 1.81fF $ **FLOATING
C2511 _0858_.A2 vssd1 1.64fF $ **FLOATING
C2512 a_11765_22325# vssd1 0.55fF $ **FLOATING
C2513 a_10551_22351# vssd1 0.61fF $ **FLOATING
C2514 a_10719_22325# vssd1 0.82fF $ **FLOATING
C2515 a_10126_22351# vssd1 0.63fF $ **FLOATING
C2516 a_10294_22325# vssd1 0.58fF $ **FLOATING
C2517 a_9853_22357# vssd1 1.43fF $ **FLOATING
C2518 _1055_.Q vssd1 6.43fF $ **FLOATING
C2519 a_9687_22357# vssd1 1.81fF $ **FLOATING
C2520 _0866_.B vssd1 7.18fF $ **FLOATING
C2521 _0868_.A2 vssd1 1.09fF $ **FLOATING
C2522 _0866_.Y vssd1 0.91fF $ **FLOATING
C2523 a_6613_22325# vssd1 0.55fF $ **FLOATING
C2524 a_26233_22895# vssd1 0.23fF $ **FLOATING
C2525 a_26743_23261# vssd1 0.61fF $ **FLOATING
C2526 a_26911_23163# vssd1 0.82fF $ **FLOATING
C2527 a_26318_23261# vssd1 0.63fF $ **FLOATING
C2528 a_26486_23007# vssd1 0.58fF $ **FLOATING
C2529 a_26045_22895# vssd1 1.43fF $ **FLOATING
C2530 a_25879_22895# vssd1 1.81fF $ **FLOATING
C2531 a_21279_22895# vssd1 0.65fF $ **FLOATING
C2532 _0933_.Q vssd1 3.77fF $ **FLOATING
C2533 a_17585_22895# vssd1 0.23fF $ **FLOATING
C2534 a_18095_23261# vssd1 0.61fF $ **FLOATING
C2535 a_18263_23163# vssd1 0.82fF $ **FLOATING
C2536 a_17670_23261# vssd1 0.63fF $ **FLOATING
C2537 a_17838_23007# vssd1 0.58fF $ **FLOATING
C2538 a_17397_22895# vssd1 1.43fF $ **FLOATING
C2539 _0932_.Q vssd1 4.54fF $ **FLOATING
C2540 a_17231_22895# vssd1 1.81fF $ **FLOATING
C2541 _0856_.Y vssd1 1.33fF $ **FLOATING
C2542 _0848_.X vssd1 1.44fF $ **FLOATING
C2543 a_12355_22901# vssd1 0.48fF $ **FLOATING
C2544 a_5466_22895# vssd1 0.26fF $ **FLOATING
C2545 a_4959_22895# vssd1 0.19fF $ **FLOATING
C2546 a_4769_22895# vssd1 0.19fF $ **FLOATING
C2547 a_4769_23145# vssd1 0.67fF $ **FLOATING
C2548 io_out[1] vssd1 3.75fF
C2549 a_12547_23145# vssd1 0.48fF $ **FLOATING
C2550 a_11435_22895# vssd1 1.20fF $ **FLOATING
C2551 a_9811_22923# vssd1 0.56fF $ **FLOATING
C2552 _0742_.A2 vssd1 3.59fF $ **FLOATING
C2553 a_4403_22869# vssd1 1.57fF $ **FLOATING
C2554 _0996_.Q vssd1 5.13fF $ **FLOATING
C2555 a_25129_23439# vssd1 0.23fF $ **FLOATING
C2556 _1054_.Q vssd1 4.86fF $ **FLOATING
C2557 a_9687_23439# vssd1 0.44fF $ **FLOATING
C2558 a_14917_23439# vssd1 0.23fF $ **FLOATING
C2559 _0726_.X vssd1 1.86fF $ **FLOATING
C2560 a_4999_23759# vssd1 0.21fF $ **FLOATING
C2561 a_25639_23439# vssd1 0.61fF $ **FLOATING
C2562 a_25807_23413# vssd1 0.82fF $ **FLOATING
C2563 a_25214_23439# vssd1 0.63fF $ **FLOATING
C2564 a_25382_23413# vssd1 0.58fF $ **FLOATING
C2565 a_24941_23445# vssd1 1.43fF $ **FLOATING
C2566 a_24775_23445# vssd1 1.81fF $ **FLOATING
C2567 a_15427_23439# vssd1 0.61fF $ **FLOATING
C2568 a_15595_23413# vssd1 0.82fF $ **FLOATING
C2569 a_15002_23439# vssd1 0.63fF $ **FLOATING
C2570 a_15170_23413# vssd1 0.58fF $ **FLOATING
C2571 a_14729_23445# vssd1 1.43fF $ **FLOATING
C2572 a_14563_23445# vssd1 1.81fF $ **FLOATING
C2573 a_11803_23439# vssd1 1.20fF $ **FLOATING
C2574 _0443_.A vssd1 1.71fF $ **FLOATING
C2575 a_7520_23555# vssd1 0.50fF $ **FLOATING
C2576 _0441_.B vssd1 15.62fF $ **FLOATING
C2577 a_6559_23552# vssd1 0.62fF $ **FLOATING
C2578 _0813_.C1 vssd1 1.93fF $ **FLOATING
C2579 _0813_.A2 vssd1 11.70fF $ **FLOATING
C2580 a_4863_23413# vssd1 0.79fF $ **FLOATING
C2581 a_2686_23439# vssd1 4.03fF $ **FLOATING
C2582 temp1.capload\[10\].cap_40.HI vssd1 0.42fF $ **FLOATING
C2583 _0928_.Q vssd1 6.23fF $ **FLOATING
C2584 a_27337_23983# vssd1 0.23fF $ **FLOATING
C2585 a_27847_24349# vssd1 0.61fF $ **FLOATING
C2586 a_28015_24251# vssd1 0.82fF $ **FLOATING
C2587 a_27422_24349# vssd1 0.63fF $ **FLOATING
C2588 a_27590_24095# vssd1 0.58fF $ **FLOATING
C2589 a_27149_23983# vssd1 1.43fF $ **FLOATING
C2590 _0928_.D vssd1 6.29fF $ **FLOATING
C2591 a_26983_23983# vssd1 1.81fF $ **FLOATING
C2592 _1021_.Q vssd1 4.97fF $ **FLOATING
C2593 a_4356_23983# vssd1 0.54fF $ **FLOATING
C2594 a_21357_23983# vssd1 0.23fF $ **FLOATING
C2595 a_21867_24349# vssd1 0.61fF $ **FLOATING
C2596 a_22035_24251# vssd1 0.82fF $ **FLOATING
C2597 a_21442_24349# vssd1 0.63fF $ **FLOATING
C2598 a_21610_24095# vssd1 0.58fF $ **FLOATING
C2599 a_21169_23983# vssd1 1.43fF $ **FLOATING
C2600 a_21003_23983# vssd1 1.81fF $ **FLOATING
C2601 a_12622_24233# vssd1 0.22fF $ **FLOATING
C2602 a_11251_24233# vssd1 0.39fF $ **FLOATING
C2603 _0723_.X vssd1 2.16fF $ **FLOATING
C2604 io_out[4] vssd1 3.84fF
C2605 a_4439_24233# vssd1 0.34fF $ **FLOATING
C2606 a_1863_24233# vssd1 0.32fF $ **FLOATING
C2607 io_out[3] vssd1 1.22fF
C2608 a_12316_24135# vssd1 0.70fF $ **FLOATING
C2609 a_10055_23983# vssd1 1.20fF $ **FLOATING
C2610 a_6416_24233# vssd1 0.50fF $ **FLOATING
C2611 _0774_.A2 vssd1 5.07fF $ **FLOATING
C2612 _0765_.B1 vssd1 5.19fF $ **FLOATING
C2613 a_1585_24135# vssd1 0.77fF $ **FLOATING
C2614 a_14651_24527# vssd1 0.25fF $ **FLOATING
C2615 a_12995_24527# vssd1 0.25fF $ **FLOATING
C2616 a_11711_24527# vssd1 0.44fF $ **FLOATING
C2617 a_10055_24527# vssd1 0.44fF $ **FLOATING
C2618 _0852_.X vssd1 14.45fF $ **FLOATING
C2619 temp1.capload\[1\].cap.Y vssd1 0.28fF $ **FLOATING
C2620 temp1.capload\[11\].cap.Y vssd1 0.28fF $ **FLOATING
C2621 a_16904_24643# vssd1 0.50fF $ **FLOATING
C2622 _0860_.B vssd1 8.22fF $ **FLOATING
C2623 a_14433_24501# vssd1 0.55fF $ **FLOATING
C2624 a_12777_24501# vssd1 0.55fF $ **FLOATING
C2625 _0860_.A vssd1 25.51fF $ **FLOATING
C2626 _0838_.A0 vssd1 7.34fF $ **FLOATING
C2627 a_2833_24759# vssd1 0.77fF $ **FLOATING
C2628 a_2655_24501# vssd1 0.83fF $ **FLOATING
C2629 _0998_.Q vssd1 5.24fF $ **FLOATING
C2630 a_12815_25071# vssd1 0.28fF $ **FLOATING
C2631 a_27337_25071# vssd1 0.23fF $ **FLOATING
C2632 a_27847_25437# vssd1 0.61fF $ **FLOATING
C2633 a_28015_25339# vssd1 0.82fF $ **FLOATING
C2634 a_27422_25437# vssd1 0.63fF $ **FLOATING
C2635 a_27590_25183# vssd1 0.58fF $ **FLOATING
C2636 a_27149_25071# vssd1 1.43fF $ **FLOATING
C2637 _0998_.D vssd1 7.79fF $ **FLOATING
C2638 a_26983_25071# vssd1 1.81fF $ **FLOATING
C2639 _0854_.X vssd1 14.89fF $ **FLOATING
C2640 ANTENNA_7.DIODE vssd1 21.52fF $ **FLOATING
C2641 _0854_.B vssd1 16.12fF $ **FLOATING
C2642 _0850_.Y vssd1 12.52fF $ **FLOATING
C2643 a_11842_25321# vssd1 0.33fF $ **FLOATING
C2644 a_9613_25045# vssd1 0.61fF $ **FLOATING
C2645 a_25707_25321# vssd1 0.64fF $ **FLOATING
C2646 a_11685_25045# vssd1 0.72fF $ **FLOATING
C2647 a_9184_25223# vssd1 0.59fF $ **FLOATING
C2648 _0816_.S vssd1 4.79fF $ **FLOATING
C2649 a_7389_25335# vssd1 0.76fF $ **FLOATING
C2650 _0788_.C vssd1 2.44fF $ **FLOATING
C2651 a_5913_25335# vssd1 0.60fF $ **FLOATING
C2652 a_5813_25117# vssd1 0.49fF $ **FLOATING
C2653 _1077_.Q vssd1 6.88fF $ **FLOATING
C2654 a_2405_25071# vssd1 0.23fF $ **FLOATING
C2655 _0850_.A vssd1 23.23fF $ **FLOATING
C2656 _0842_.A0 vssd1 28.21fF $ **FLOATING
C2657 _0829_.A1 vssd1 21.34fF $ **FLOATING
C2658 a_4213_25223# vssd1 0.77fF $ **FLOATING
C2659 a_4035_25045# vssd1 0.83fF $ **FLOATING
C2660 a_2915_25437# vssd1 0.61fF $ **FLOATING
C2661 a_3083_25339# vssd1 0.82fF $ **FLOATING
C2662 a_2490_25437# vssd1 0.63fF $ **FLOATING
C2663 a_2658_25183# vssd1 0.58fF $ **FLOATING
C2664 a_2217_25071# vssd1 1.43fF $ **FLOATING
C2665 a_2051_25071# vssd1 1.81fF $ **FLOATING
C2666 a_25589_25615# vssd1 0.23fF $ **FLOATING
C2667 _1061_.Q vssd1 5.54fF $ **FLOATING
C2668 a_16123_25615# vssd1 0.25fF $ **FLOATING
C2669 a_10788_25615# vssd1 0.24fF $ **FLOATING
C2670 a_18689_25615# vssd1 0.23fF $ **FLOATING
C2671 _0861_.X vssd1 16.46fF $ **FLOATING
C2672 a_6809_25615# vssd1 0.20fF $ **FLOATING
C2673 a_13183_25615# vssd1 0.53fF $ **FLOATING
C2674 _0828_.Y vssd1 0.83fF $ **FLOATING
C2675 a_5547_25615# vssd1 0.39fF $ **FLOATING
C2676 io_out[5] vssd1 4.28fF
C2677 _0839_.Y vssd1 2.66fF $ **FLOATING
C2678 _1078_.Q vssd1 14.51fF $ **FLOATING
C2679 a_1591_25615# vssd1 0.39fF $ **FLOATING
C2680 a_2773_25615# vssd1 0.23fF $ **FLOATING
C2681 a_26099_25615# vssd1 0.61fF $ **FLOATING
C2682 a_26267_25589# vssd1 0.82fF $ **FLOATING
C2683 a_25674_25615# vssd1 0.63fF $ **FLOATING
C2684 a_25842_25589# vssd1 0.58fF $ **FLOATING
C2685 a_25401_25621# vssd1 1.43fF $ **FLOATING
C2686 _0993_.D vssd1 4.96fF $ **FLOATING
C2687 a_25235_25621# vssd1 1.81fF $ **FLOATING
C2688 a_19199_25615# vssd1 0.61fF $ **FLOATING
C2689 a_19367_25589# vssd1 0.82fF $ **FLOATING
C2690 a_18774_25615# vssd1 0.63fF $ **FLOATING
C2691 a_18942_25589# vssd1 0.58fF $ **FLOATING
C2692 a_18501_25621# vssd1 1.43fF $ **FLOATING
C2693 _1061_.D vssd1 5.10fF $ **FLOATING
C2694 a_18335_25621# vssd1 1.81fF $ **FLOATING
C2695 _0861_.A2 vssd1 1.51fF $ **FLOATING
C2696 _0861_.A1 vssd1 1.51fF $ **FLOATING
C2697 _0861_.B1 vssd1 20.11fF $ **FLOATING
C2698 a_15905_25589# vssd1 0.55fF $ **FLOATING
C2699 a_10515_25615# vssd1 0.57fF $ **FLOATING
C2700 _0789_.B1 vssd1 1.17fF $ **FLOATING
C2701 _0789_.A2 vssd1 2.87fF $ **FLOATING
C2702 a_6611_25589# vssd1 0.80fF $ **FLOATING
C2703 _0839_.B vssd1 2.63fF $ **FLOATING
C2704 _0840_.A1 vssd1 24.63fF $ **FLOATING
C2705 _0840_.A0 vssd1 15.37fF $ **FLOATING
C2706 a_4581_25847# vssd1 0.77fF $ **FLOATING
C2707 a_4403_25589# vssd1 0.83fF $ **FLOATING
C2708 a_3283_25615# vssd1 0.61fF $ **FLOATING
C2709 a_3451_25589# vssd1 0.97fF $ **FLOATING
C2710 a_2858_25615# vssd1 0.63fF $ **FLOATING
C2711 a_3026_25589# vssd1 0.58fF $ **FLOATING
C2712 a_2585_25621# vssd1 1.43fF $ **FLOATING
C2713 _1078_.D vssd1 1.18fF $ **FLOATING
C2714 a_2419_25621# vssd1 1.81fF $ **FLOATING
C2715 _0840_.X vssd1 1.83fF $ **FLOATING
C2716 a_25957_26159# vssd1 0.23fF $ **FLOATING
C2717 a_26467_26525# vssd1 0.61fF $ **FLOATING
C2718 a_26635_26427# vssd1 0.82fF $ **FLOATING
C2719 a_26042_26525# vssd1 0.63fF $ **FLOATING
C2720 a_26210_26271# vssd1 0.58fF $ **FLOATING
C2721 a_25769_26159# vssd1 1.43fF $ **FLOATING
C2722 _0994_.D vssd1 5.60fF $ **FLOATING
C2723 a_25603_26159# vssd1 1.81fF $ **FLOATING
C2724 _0994_.CLK vssd1 10.62fF $ **FLOATING
C2725 _1020_.Q vssd1 6.64fF $ **FLOATING
C2726 a_22185_26159# vssd1 0.23fF $ **FLOATING
C2727 a_22695_26525# vssd1 0.61fF $ **FLOATING
C2728 a_22863_26427# vssd1 0.82fF $ **FLOATING
C2729 a_22270_26525# vssd1 0.63fF $ **FLOATING
C2730 a_22438_26271# vssd1 0.58fF $ **FLOATING
C2731 a_21997_26159# vssd1 1.43fF $ **FLOATING
C2732 a_21831_26159# vssd1 1.81fF $ **FLOATING
C2733 a_16573_26159# vssd1 0.23fF $ **FLOATING
C2734 a_17083_26525# vssd1 0.61fF $ **FLOATING
C2735 a_17251_26427# vssd1 0.82fF $ **FLOATING
C2736 a_16658_26525# vssd1 0.63fF $ **FLOATING
C2737 a_16826_26271# vssd1 0.58fF $ **FLOATING
C2738 a_16385_26159# vssd1 1.43fF $ **FLOATING
C2739 _1052_.D vssd1 5.15fF $ **FLOATING
C2740 a_16219_26159# vssd1 1.81fF $ **FLOATING
C2741 a_10073_26133# vssd1 0.61fF $ **FLOATING
C2742 _0740_.X vssd1 3.06fF $ **FLOATING
C2743 _0819_.S vssd1 4.65fF $ **FLOATING
C2744 _1079_.Q vssd1 8.74fF $ **FLOATING
C2745 a_4337_26159# vssd1 0.23fF $ **FLOATING
C2746 a_13183_26159# vssd1 0.53fF $ **FLOATING
C2747 a_12355_26159# vssd1 0.53fF $ **FLOATING
C2748 a_9644_26311# vssd1 0.59fF $ **FLOATING
C2749 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 1.13fF $ **FLOATING
C2750 a_8215_26159# vssd1 0.53fF $ **FLOATING
C2751 _0817_.A vssd1 1.74fF $ **FLOATING
C2752 a_7435_26324# vssd1 0.52fF $ **FLOATING
C2753 a_6600_26409# vssd1 0.50fF $ **FLOATING
C2754 a_4847_26525# vssd1 0.61fF $ **FLOATING
C2755 a_5015_26427# vssd1 0.82fF $ **FLOATING
C2756 a_4422_26525# vssd1 0.63fF $ **FLOATING
C2757 a_4590_26271# vssd1 0.58fF $ **FLOATING
C2758 a_4149_26159# vssd1 1.43fF $ **FLOATING
C2759 a_3983_26159# vssd1 1.81fF $ **FLOATING
C2760 clkbuf_1_0__f_net57.X vssd1 4.02fF $ **FLOATING
C2761 a_1674_26159# vssd1 4.03fF $ **FLOATING
C2762 _0995_.Q vssd1 7.19fF $ **FLOATING
C2763 a_23381_26703# vssd1 0.23fF $ **FLOATING
C2764 a_19517_26703# vssd1 0.23fF $ **FLOATING
C2765 a_23891_26703# vssd1 0.61fF $ **FLOATING
C2766 a_24059_26677# vssd1 0.82fF $ **FLOATING
C2767 a_23466_26703# vssd1 0.63fF $ **FLOATING
C2768 a_23634_26677# vssd1 0.58fF $ **FLOATING
C2769 a_23193_26709# vssd1 1.43fF $ **FLOATING
C2770 _0994_.Q vssd1 6.77fF $ **FLOATING
C2771 a_23027_26709# vssd1 1.81fF $ **FLOATING
C2772 _0995_.CLK vssd1 16.19fF $ **FLOATING
C2773 a_20027_26703# vssd1 0.61fF $ **FLOATING
C2774 a_20195_26677# vssd1 0.82fF $ **FLOATING
C2775 a_19602_26703# vssd1 0.63fF $ **FLOATING
C2776 a_19770_26677# vssd1 0.58fF $ **FLOATING
C2777 a_19329_26709# vssd1 1.43fF $ **FLOATING
C2778 _1018_.D vssd1 7.14fF $ **FLOATING
C2779 a_19163_26709# vssd1 1.81fF $ **FLOATING
C2780 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.HI vssd1 0.42fF $ **FLOATING
C2781 a_14011_26703# vssd1 0.53fF $ **FLOATING
C2782 a_13183_26703# vssd1 0.53fF $ **FLOATING
C2783 a_4984_26703# vssd1 0.43fF $ **FLOATING
C2784 a_4729_26703# vssd1 0.32fF $ **FLOATING
C2785 temp1.capload\[2\].cap.Y vssd1 0.28fF $ **FLOATING
C2786 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 1.43fF $ **FLOATING
C2787 _0752_.Y vssd1 5.97fF $ **FLOATING
C2788 a_6559_27023# vssd1 0.28fF $ **FLOATING
C2789 a_5177_27023# vssd1 0.27fF $ **FLOATING
C2790 _1075_.Q vssd1 18.26fF $ **FLOATING
C2791 a_3141_26703# vssd1 0.23fF $ **FLOATING
C2792 a_12189_27001# vssd1 0.61fF $ **FLOATING
C2793 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 8.21fF $ **FLOATING
C2794 a_11760_26935# vssd1 0.59fF $ **FLOATING
C2795 _0835_.A1 vssd1 22.48fF $ **FLOATING
C2796 a_3651_26703# vssd1 0.61fF $ **FLOATING
C2797 a_3819_26677# vssd1 0.97fF $ **FLOATING
C2798 a_3226_26703# vssd1 0.63fF $ **FLOATING
C2799 a_3394_26677# vssd1 0.58fF $ **FLOATING
C2800 a_2953_26709# vssd1 1.43fF $ **FLOATING
C2801 _0835_.Y vssd1 1.65fF $ **FLOATING
C2802 a_2787_26709# vssd1 1.81fF $ **FLOATING
C2803 a_1757_26703# vssd1 0.85fF $ **FLOATING
C2804 _0831_.D vssd1 6.25fF $ **FLOATING
C2805 _0831_.B vssd1 1.79fF $ **FLOATING
C2806 a_1591_26703# vssd1 0.60fF $ **FLOATING
C2807 _1019_.Q vssd1 5.76fF $ **FLOATING
C2808 a_21081_27247# vssd1 0.23fF $ **FLOATING
C2809 a_21591_27613# vssd1 0.61fF $ **FLOATING
C2810 a_21759_27515# vssd1 0.82fF $ **FLOATING
C2811 a_21166_27613# vssd1 0.63fF $ **FLOATING
C2812 a_21334_27359# vssd1 0.58fF $ **FLOATING
C2813 a_20893_27247# vssd1 1.43fF $ **FLOATING
C2814 _1019_.D vssd1 4.85fF $ **FLOATING
C2815 a_20727_27247# vssd1 1.81fF $ **FLOATING
C2816 _1019_.CLK vssd1 13.01fF $ **FLOATING
C2817 a_18059_27247# vssd1 0.53fF $ **FLOATING
C2818 temp1.dac.vdac_single.einvp_batch\[0\].vref.TE vssd1 1.45fF $ **FLOATING
C2819 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.LO vssd1 0.48fF $ **FLOATING
C2820 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI vssd1 1.06fF $ **FLOATING
C2821 a_7385_27247# vssd1 0.27fF $ **FLOATING
C2822 temp1.capload\[10\].cap.Y vssd1 0.28fF $ **FLOATING
C2823 a_7192_27497# vssd1 0.43fF $ **FLOATING
C2824 a_6937_27497# vssd1 0.32fF $ **FLOATING
C2825 _1076_.Q vssd1 19.36fF $ **FLOATING
C2826 a_2313_27247# vssd1 0.23fF $ **FLOATING
C2827 a_11067_27247# vssd1 0.53fF $ **FLOATING
C2828 a_10239_27247# vssd1 0.53fF $ **FLOATING
C2829 temp1.capload\[10\].cap.A vssd1 5.24fF $ **FLOATING
C2830 _0837_.A1 vssd1 18.63fF $ **FLOATING
C2831 a_4802_27247# vssd1 4.03fF $ **FLOATING
C2832 clkbuf_0__0390_.A vssd1 1.35fF $ **FLOATING
C2833 a_4075_27247# vssd1 0.52fF $ **FLOATING
C2834 _0832_.A vssd1 1.67fF $ **FLOATING
C2835 a_2823_27613# vssd1 0.61fF $ **FLOATING
C2836 a_2991_27515# vssd1 0.97fF $ **FLOATING
C2837 a_2398_27613# vssd1 0.63fF $ **FLOATING
C2838 a_2566_27359# vssd1 0.58fF $ **FLOATING
C2839 a_2125_27247# vssd1 1.43fF $ **FLOATING
C2840 _0837_.Y vssd1 2.96fF $ **FLOATING
C2841 a_1959_27247# vssd1 1.81fF $ **FLOATING
C2842 _1053_.Q vssd1 5.35fF $ **FLOATING
C2843 a_15285_27791# vssd1 0.23fF $ **FLOATING
C2844 _0824_.Y vssd1 3.90fF $ **FLOATING
C2845 a_12525_27791# vssd1 0.23fF $ **FLOATING
C2846 _0815_.Y vssd1 2.54fF $ **FLOATING
C2847 a_9871_27791# vssd1 0.53fF $ **FLOATING
C2848 a_8583_27791# vssd1 0.53fF $ **FLOATING
C2849 a_4811_27791# vssd1 0.39fF $ **FLOATING
C2850 a_1775_27791# vssd1 0.39fF $ **FLOATING
C2851 a_7755_27791# vssd1 0.53fF $ **FLOATING
C2852 _0787_.X vssd1 1.55fF $ **FLOATING
C2853 _0843_.Y vssd1 2.52fF $ **FLOATING
C2854 a_15795_27791# vssd1 0.61fF $ **FLOATING
C2855 a_15963_27765# vssd1 0.82fF $ **FLOATING
C2856 a_15370_27791# vssd1 0.63fF $ **FLOATING
C2857 a_15538_27765# vssd1 0.58fF $ **FLOATING
C2858 a_15097_27797# vssd1 1.43fF $ **FLOATING
C2859 _1053_.D vssd1 6.13fF $ **FLOATING
C2860 a_14931_27797# vssd1 1.81fF $ **FLOATING
C2861 _1053_.CLK vssd1 14.50fF $ **FLOATING
C2862 a_12348_27791# vssd1 0.50fF $ **FLOATING
C2863 a_12242_27791# vssd1 0.58fF $ **FLOATING
C2864 a_12065_27791# vssd1 0.50fF $ **FLOATING
C2865 a_11746_27791# vssd1 0.54fF $ **FLOATING
C2866 _0823_.A vssd1 1.15fF $ **FLOATING
C2867 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 3.26fF $ **FLOATING
C2868 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 2.11fF $ **FLOATING
C2869 a_6600_27907# vssd1 0.50fF $ **FLOATING
C2870 _0844_.B vssd1 7.44fF $ **FLOATING
C2871 a_2686_27791# vssd1 4.03fF $ **FLOATING
C2872 _0843_.B vssd1 2.73fF $ **FLOATING
C2873 temp1.capload\[5\].cap.Y vssd1 0.28fF $ **FLOATING
C2874 temp1.capload\[12\].cap.Y vssd1 0.28fF $ **FLOATING
C2875 a_14287_28335# vssd1 0.53fF $ **FLOATING
C2876 a_13183_28335# vssd1 0.53fF $ **FLOATING
C2877 a_12355_28335# vssd1 0.53fF $ **FLOATING
C2878 a_11527_28335# vssd1 0.53fF $ **FLOATING
C2879 temp1.capload\[4\].cap_49.HI vssd1 0.42fF $ **FLOATING
C2880 _0821_.Y vssd1 2.07fF $ **FLOATING
C2881 _0820_.A vssd1 2.05fF $ **FLOATING
C2882 a_8079_28500# vssd1 0.52fF $ **FLOATING
C2883 _0821_.B vssd1 3.65fF $ **FLOATING
C2884 a_6651_28335# vssd1 0.65fF $ **FLOATING
C2885 _0833_.Y vssd1 1.96fF $ **FLOATING
C2886 a_5823_28585# vssd1 0.39fF $ **FLOATING
C2887 _1081_.Q vssd1 6.28fF $ **FLOATING
C2888 a_4337_28335# vssd1 0.23fF $ **FLOATING
C2889 _0833_.A vssd1 18.64fF $ **FLOATING
C2890 a_4847_28701# vssd1 0.61fF $ **FLOATING
C2891 a_5015_28603# vssd1 0.82fF $ **FLOATING
C2892 a_4422_28701# vssd1 0.63fF $ **FLOATING
C2893 a_4590_28447# vssd1 0.58fF $ **FLOATING
C2894 a_4149_28335# vssd1 1.43fF $ **FLOATING
C2895 a_3983_28335# vssd1 1.81fF $ **FLOATING
C2896 _1080_.Q vssd1 11.79fF $ **FLOATING
C2897 a_2405_28335# vssd1 0.23fF $ **FLOATING
C2898 a_2915_28701# vssd1 0.61fF $ **FLOATING
C2899 a_3083_28603# vssd1 0.82fF $ **FLOATING
C2900 a_2490_28701# vssd1 0.63fF $ **FLOATING
C2901 a_2658_28447# vssd1 0.58fF $ **FLOATING
C2902 a_2217_28335# vssd1 1.43fF $ **FLOATING
C2903 a_2051_28335# vssd1 1.81fF $ **FLOATING
C2904 a_14195_28879# vssd1 0.53fF $ **FLOATING
C2905 a_13367_28879# vssd1 0.53fF $ **FLOATING
C2906 a_12355_28879# vssd1 0.53fF $ **FLOATING
C2907 temp1.capload\[14\].cap.Y vssd1 0.28fF $ **FLOATING
C2908 a_10699_28879# vssd1 0.53fF $ **FLOATING
C2909 temp1.capload\[11\].cap_41.LO vssd1 5.31fF $ **FLOATING
C2910 a_15023_28887# vssd1 0.65fF $ **FLOATING
C2911 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 4.73fF $ **FLOATING
C2912 a_9779_28879# vssd1 0.52fF $ **FLOATING
C2913 temp1.capload\[11\].cap_41.HI vssd1 0.42fF $ **FLOATING
C2914 temp1.capload\[2\].cap_47.LO vssd1 2.09fF $ **FLOATING
C2915 temp1.capload\[0\].cap_39.HI vssd1 0.42fF $ **FLOATING
C2916 temp1.capload\[2\].cap_47.HI vssd1 0.42fF $ **FLOATING
C2917 a_1775_28879# vssd1 0.39fF $ **FLOATING
C2918 _0825_.X vssd1 0.92fF $ **FLOATING
C2919 a_5541_29199# vssd1 0.17fF $ **FLOATING
C2920 _0764_.X vssd1 4.22fF $ **FLOATING
C2921 _0836_.Y vssd1 3.87fF $ **FLOATING
C2922 a_7037_29177# vssd1 0.61fF $ **FLOATING
C2923 _0825_.A0 vssd1 9.88fF $ **FLOATING
C2924 _0825_.A1 vssd1 9.20fF $ **FLOATING
C2925 a_6608_29111# vssd1 0.59fF $ **FLOATING
C2926 _0764_.A1 vssd1 7.01fF $ **FLOATING
C2927 _0825_.S vssd1 7.27fF $ **FLOATING
C2928 a_5323_29111# vssd1 0.55fF $ **FLOATING
C2929 a_2686_28879# vssd1 4.03fF $ **FLOATING
C2930 clkbuf_1_1__f__0390_.A vssd1 7.55fF $ **FLOATING
C2931 _0836_.A vssd1 20.22fF $ **FLOATING
C2932 a_15667_29423# vssd1 0.53fF $ **FLOATING
C2933 a_14839_29423# vssd1 0.53fF $ **FLOATING
C2934 a_13367_29423# vssd1 0.53fF $ **FLOATING
C2935 a_12539_29423# vssd1 0.53fF $ **FLOATING
C2936 a_11619_29423# vssd1 0.70fF $ **FLOATING
C2937 fanout11.A vssd1 2.79fF $ **FLOATING
C2938 a_10791_29423# vssd1 0.53fF $ **FLOATING
C2939 a_9963_29423# vssd1 0.53fF $ **FLOATING
C2940 temp1.capload\[7\].cap_52.HI vssd1 0.42fF $ **FLOATING
C2941 a_7479_29673# vssd1 0.39fF $ **FLOATING
C2942 a_4441_29423# vssd1 0.27fF $ **FLOATING
C2943 _0445_.X vssd1 2.63fF $ **FLOATING
C2944 _0445_.A vssd1 12.69fF $ **FLOATING
C2945 a_6191_29423# vssd1 0.53fF $ **FLOATING
C2946 a_5273_29687# vssd1 0.76fF $ **FLOATING
C2947 _0445_.B vssd1 8.81fF $ **FLOATING
C2948 a_4248_29673# vssd1 0.43fF $ **FLOATING
C2949 _0845_.Y vssd1 2.13fF $ **FLOATING
C2950 a_3993_29673# vssd1 0.32fF $ **FLOATING
C2951 _0845_.A2 vssd1 8.88fF $ **FLOATING
C2952 _0845_.A1 vssd1 18.82fF $ **FLOATING
C2953 _0845_.B1 vssd1 1.83fF $ **FLOATING
C2954 a_1766_29423# vssd1 4.03fF $ **FLOATING
C2955 temp1.inv1_1.Y vssd1 4.15fF $ **FLOATING
C2956 a_15667_29967# vssd1 0.53fF $ **FLOATING
C2957 a_14839_29967# vssd1 0.53fF $ **FLOATING
C2958 a_14011_29967# vssd1 0.53fF $ **FLOATING
C2959 a_13183_29967# vssd1 0.53fF $ **FLOATING
C2960 a_12355_29967# vssd1 0.53fF $ **FLOATING
C2961 temp1.capload\[9\].cap.Y vssd1 0.28fF $ **FLOATING
C2962 a_10791_29967# vssd1 0.53fF $ **FLOATING
C2963 a_9963_29967# vssd1 0.53fF $ **FLOATING
C2964 a_8767_29967# vssd1 0.53fF $ **FLOATING
C2965 a_1975_29967# vssd1 0.22fF $ **FLOATING
C2966 a_7387_29967# vssd1 0.53fF $ **FLOATING
C2967 a_6559_29967# vssd1 0.53fF $ **FLOATING
C2968 a_5361_30287# vssd1 0.28fF $ **FLOATING
C2969 io_out[6] vssd1 2.62fF
C2970 _0847_.X vssd1 2.58fF $ **FLOATING
C2971 _0809_.A1 vssd1 4.55fF $ **FLOATING
C2972 _0809_.B2 vssd1 7.93fF $ **FLOATING
C2973 _0827_.A vssd1 15.60fF $ **FLOATING
C2974 a_5141_30199# vssd1 0.76fF $ **FLOATING
C2975 a_2962_29967# vssd1 4.03fF $ **FLOATING
C2976 clkbuf_0_temp1.i_precharge_n.A vssd1 4.61fF $ **FLOATING
C2977 _0845_.C1 vssd1 25.14fF $ **FLOATING
C2978 _0847_.B1 vssd1 6.39fF $ **FLOATING
C2979 _0847_.A1 vssd1 3.27fF $ **FLOATING
C2980 _0847_.A2 vssd1 16.60fF $ **FLOATING
C2981 _0847_.A3 vssd1 15.69fF $ **FLOATING
C2982 a_1735_29941# vssd1 1.12fF $ **FLOATING
C2983 a_15667_30511# vssd1 0.70fF $ **FLOATING
C2984 fanout13.A vssd1 7.82fF $ **FLOATING
C2985 a_14839_30511# vssd1 0.53fF $ **FLOATING
C2986 a_13367_30511# vssd1 0.53fF $ **FLOATING
C2987 a_12631_30511# vssd1 0.65fF $ **FLOATING
C2988 a_4342_30761# vssd1 0.22fF $ **FLOATING
C2989 _0798_.X vssd1 1.63fF $ **FLOATING
C2990 a_11803_30511# vssd1 0.53fF $ **FLOATING
C2991 a_10975_30511# vssd1 0.53fF $ **FLOATING
C2992 a_10147_30511# vssd1 0.53fF $ **FLOATING
C2993 a_9319_30511# vssd1 0.53fF $ **FLOATING
C2994 a_8215_30511# vssd1 0.53fF $ **FLOATING
C2995 a_7295_30511# vssd1 0.53fF $ **FLOATING
C2996 a_5078_30511# vssd1 4.03fF $ **FLOATING
C2997 _0798_.A2 vssd1 17.73fF $ **FLOATING
C2998 _0798_.A1 vssd1 3.63fF $ **FLOATING
C2999 a_4036_30663# vssd1 0.70fF $ **FLOATING
C3000 a_1766_30511# vssd1 4.03fF $ **FLOATING
C3001 a_14563_31055# vssd1 0.53fF $ **FLOATING
C3002 a_13735_31055# vssd1 0.53fF $ **FLOATING
C3003 a_11711_31055# vssd1 0.53fF $ **FLOATING
C3004 a_10791_31055# vssd1 0.53fF $ **FLOATING
C3005 a_9963_31055# vssd1 0.53fF $ **FLOATING
C3006 a_8767_31055# vssd1 0.53fF $ **FLOATING
C3007 a_7939_31055# vssd1 0.53fF $ **FLOATING
C3008 a_7111_31055# vssd1 0.53fF $ **FLOATING
C3009 a_5639_31055# vssd1 0.53fF $ **FLOATING
C3010 a_4811_31055# vssd1 0.53fF $ **FLOATING
C3011 _0444_.Y vssd1 3.03fF $ **FLOATING
C3012 a_1775_31375# vssd1 0.28fF $ **FLOATING
C3013 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.A vssd1 6.79fF $ **FLOATING
C3014 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd.TE vssd1 6.81fF $ **FLOATING
C3015 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.A vssd1 6.28fF $ **FLOATING
C3016 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd.TE vssd1 9.53fF $ **FLOATING
C3017 a_12999_31055# vssd1 0.70fF $ **FLOATING
C3018 fanout9.A vssd1 2.68fF $ **FLOATING
C3019 a_2686_31055# vssd1 4.03fF $ **FLOATING
C3020 clkbuf_1_0__f_temp1.dcdel_capnode_notouch_.A vssd1 6.13fF $ **FLOATING
C3021 _0444_.A vssd1 15.85fF $ **FLOATING
C3022 _0444_.B vssd1 15.94fF $ **FLOATING
C3023 temp1.capload\[0\].cap.Y vssd1 0.28fF $ **FLOATING
C3024 temp1.capload\[3\].cap.Y vssd1 0.28fF $ **FLOATING
C3025 temp1.capload\[15\].cap.Y vssd1 0.28fF $ **FLOATING
C3026 temp1.capload\[6\].cap.Y vssd1 0.28fF $ **FLOATING
C3027 temp1.capload\[0\].cap.A vssd1 5.23fF $ **FLOATING
C3028 temp1.capload\[15\].cap.B vssd1 16.89fF $ **FLOATING
C3029 temp1.capload\[3\].cap.A vssd1 1.90fF $ **FLOATING
C3030 temp1.capload\[3\].cap_48.HI vssd1 0.42fF $ **FLOATING
C3031 a_12355_31599# vssd1 0.65fF $ **FLOATING
C3032 a_11527_31599# vssd1 0.53fF $ **FLOATING
C3033 a_10699_31599# vssd1 0.53fF $ **FLOATING
C3034 a_9871_31599# vssd1 0.53fF $ **FLOATING
C3035 fanout10.A vssd1 7.56fF $ **FLOATING
C3036 temp1.capload\[9\].cap_54.LO vssd1 2.64fF $ **FLOATING
C3037 temp1.capload\[9\].cap_54.HI vssd1 0.42fF $ **FLOATING
C3038 a_8215_31599# vssd1 0.53fF $ **FLOATING
C3039 temp1.capload\[8\].cap_53.HI vssd1 0.42fF $ **FLOATING
C3040 temp1.capload\[12\].cap_42.LO vssd1 3.62fF $ **FLOATING
C3041 temp1.capload\[12\].cap_42.HI vssd1 0.42fF $ **FLOATING
C3042 io_out[7] vssd1 2.48fF
C3043 a_4065_31849# vssd1 0.21fF $ **FLOATING
C3044 a_5547_31599# vssd1 0.53fF $ **FLOATING
C3045 a_3983_31849# vssd1 1.01fF $ **FLOATING
C3046 _0814_.A2 vssd1 12.41fF $ **FLOATING
C3047 _0814_.A1 vssd1 4.50fF $ **FLOATING
C3048 _0814_.B1 vssd1 3.58fF $ **FLOATING
C3049 _0814_.B2 vssd1 4.88fF $ **FLOATING
C3050 a_1674_31599# vssd1 4.03fF $ **FLOATING
C3051 clkbuf_1_0__f_temp1.i_precharge_n.A vssd1 6.64fF $ **FLOATING
C3052 temp1.capload\[4\].cap.Y vssd1 0.28fF $ **FLOATING
C3053 temp1.capload\[13\].cap.Y vssd1 0.28fF $ **FLOATING
C3054 temp1.capload\[15\].cap_45.LO vssd1 1.87fF $ **FLOATING
C3055 temp1.capload\[7\].cap.Y vssd1 0.28fF $ **FLOATING
C3056 temp1.capload\[4\].cap.A vssd1 5.05fF $ **FLOATING
C3057 temp1.capload\[7\].cap.A vssd1 4.08fF $ **FLOATING
C3058 temp1.capload\[13\].cap.A vssd1 2.21fF $ **FLOATING
C3059 temp1.capload\[15\].cap_45.HI vssd1 0.42fF $ **FLOATING
C3060 temp1.capload\[8\].cap.Y vssd1 0.28fF $ **FLOATING
C3061 temp1.capload\[8\].cap.A vssd1 3.23fF $ **FLOATING
C3062 temp1.capload\[13\].cap.B vssd1 10.62fF $ **FLOATING
C3063 temp1.capload\[14\].cap_44.LO vssd1 2.94fF $ **FLOATING
C3064 temp1.capload\[13\].cap_43.HI vssd1 0.42fF $ **FLOATING
C3065 a_10699_32143# vssd1 0.53fF $ **FLOATING
C3066 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.TE vssd1 9.80fF $ **FLOATING
C3067 temp1.capload\[6\].cap_51.LO vssd1 4.17fF $ **FLOATING
C3068 temp1.capload\[14\].cap_44.HI vssd1 0.42fF $ **FLOATING
C3069 a_9135_32143# vssd1 0.53fF $ **FLOATING
C3070 a_8215_32143# vssd1 0.53fF $ **FLOATING
C3071 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref.TE vssd1 9.19fF $ **FLOATING
C3072 temp1.capload\[1\].cap_46.LO vssd1 4.90fF $ **FLOATING
C3073 temp1.capload\[6\].cap_51.HI vssd1 0.42fF $ **FLOATING
C3074 temp1.capload\[5\].cap_50.LO vssd1 4.31fF $ **FLOATING
C3075 temp1.capload\[1\].cap_46.HI vssd1 0.42fF $ **FLOATING
C3076 temp1.capload\[5\].cap_50.HI vssd1 0.42fF $ **FLOATING
C3077 a_4811_32143# vssd1 0.53fF $ **FLOATING
C3078 temp1.dcdc.Z vssd1 2.29fF $ **FLOATING
C3079 a_3983_32143# vssd1 0.53fF $ **FLOATING
C3080 clkbuf_1_1__f_net57.X vssd1 6.92fF $ **FLOATING
C3081 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.A vssd1 7.00fF $ **FLOATING
C3082 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd.TE vssd1 8.46fF $ **FLOATING
C3083 temp1.dcdc.A vssd1 3.13fF $ **FLOATING
C3084 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref.Z vssd1 62.60fF $ **FLOATING
C3085 a_1674_32143# vssd1 4.03fF $ **FLOATING
C3086 clkbuf_1_1__f_net57.A vssd1 7.01fF $ **FLOATING
C3087 vccd1 vssd1 3659.64fF
.ends

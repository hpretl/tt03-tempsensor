* PEX produced on Sat Dec 30 07:12:47 PM CET 2023 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from hpretl_tt03_temperature_sensor.ext - technology: sky130A

.subckt hpretl_tt03_temperature_sensor
+ io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] 
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
X0 a_5418_1653# a_5250_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1 a_6808_11177# a_6559_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X3 _044_ a_5864_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4 temp1.dcdel_capnode_notouch_ temp1.i_precharge_n a_6736_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X7 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11868_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X8 temp1.dac_vout_notouch_ net8 a_10764_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X9 a_3885_5737# _096_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X10 a_4541_10089# temp_delay_last vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9568_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X13 vssd1 _060_ a_4069_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X14 vccd1 net3 a_10423_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X16 vssd1 net4 a_11703_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X17 vssd1 net5 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 vssd1 net11 a_2511_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_5989_2767# ctr\[10\] a_5905_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X21 vssd1 a_3116_7637# _035_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X22 vssd1 _045_ _050_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 vssd1 _076_ a_7203_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 vssd1 _045_ a_5363_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 a_6706_4511# a_6538_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X26 a_6706_4511# a_6538_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X27 a_10764_3855# a_10515_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X28 a_2397_4399# a_1407_4399# a_2271_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X30 vccd1 ctr\[1\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X31 a_9224_5487# _080_ a_9034_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X34 temp1.dac_vout_notouch_ net7 a_11428_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X35 a_8164_4087# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X36 vssd1 a_2289_3829# _014_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X37 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11711_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X39 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11408_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X40 vccd1 a_7111_6031# _093_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X41 vccd1 ctr\[1\] a_5763_9867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X42 vccd1 net19 temp1.capload\[15\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X43 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_10028_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X44 vccd1 a_2106_5599# a_2033_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X45 a_2690_11837# a_2303_11703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X46 a_3245_7663# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X47 vccd1 a_2755_11689# a_2762_11593# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X48 vccd1 a_6503_9117# a_6671_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X49 a_6265_4399# a_6099_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X50 _070_ a_5324_7637# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X51 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 _087_ a_7295_5059# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X55 vccd1 a_6671_9019# ctr\[2\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X56 vccd1 _055_ a_2507_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X57 a_5849_9867# _070_ a_5763_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X58 a_3134_8207# a_2695_8213# a_3049_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X59 _057_ a_1427_3087# a_1665_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X60 a_12328_11177# a_12079_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X61 vssd1 a_1731_2388# _015_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X63 a_2104_8527# io_out[1] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X64 a_2033_5853# a_1499_5487# a_1938_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X66 vssd1 _070_ a_4259_8757# vssd1 sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X67 vccd1 a_4036_7637# _034_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X68 vssd1 a_7348_8725# temp1.dac.vdac_single.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X69 a_6541_6031# a_6375_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X70 a_11795_2223# net7 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X71 a_8951_6825# _095_ a_9034_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X72 a_12256_7439# net29 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X73 a_7072_10901# _073_ a_7201_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X74 a_2104_10703# a_1878_10499# a_1735_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X75 io_out[3] a_2442_10092# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X76 a_1846_1501# a_1573_1135# a_1761_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X77 a_1735_7093# a_1878_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X78 a_5207_8207# a_4425_8213# a_5123_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X79 vccd1 _026_ a_7564_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X80 net5 a_10239_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X81 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10415_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X82 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12236_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X83 a_9568_4943# a_9319_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X85 _045_ _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X86 vssd1 ctr\[8\] a_1509_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X87 a_8681_4649# _026_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R0 vccd1 temp1.capload\[6\].cap_25.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X88 a_4220_10927# io_out[5] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X89 a_3260_8585# a_2861_8213# a_3134_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X90 a_6553_2883# ctr\[12\] a_6457_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_7374_9839# _070_ a_7288_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X93 vccd1 net3 a_9871_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X94 a_6729_7119# _010_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X95 vssd1 ctr\[8\] _071_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X96 vccd1 a_7902_10357# a_7829_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X97 vccd1 ctr\[9\] a_5365_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X98 a_4165_7913# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X99 a_2861_8213# a_2695_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X100 a_3215_9813# _032_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X101 a_7477_8751# _078_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X103 vccd1 a_1959_1687# _032_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X104 temp1.dac_vout_notouch_ net7 a_11960_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X105 vssd1 a_2439_4667# a_2397_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X106 a_12236_6031# a_11987_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X108 a_4238_6941# a_3799_6575# a_4153_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X109 a_2471_11703# a_2755_11689# a_2690_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X110 a_2932_9269# _032_ a_3061_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X111 a_10255_9001# _026_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X112 vccd1 _080_ a_8951_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X113 a_4613_5487# _090_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X114 _083_ a_8307_7235# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X115 a_9588_9839# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X116 a_10968_3311# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X118 vssd1 a_3024_6005# _037_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X119 vccd1 _060_ _064_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X121 a_6009_3317# _049_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X122 a_3339_7663# ctr\[4\] a_3245_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X123 a_11612_10927# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X124 a_9033_8751# _093_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X125 a_7545_5059# _082_ a_7473_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X126 temp1.capload\[4\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X127 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10699_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X128 vccd1 net10 a_5639_6397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X129 a_9779_8751# _089_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X130 vccd1 io_in[1] a_1407_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X131 io_out[6] a_3215_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X132 a_1878_8323# _034_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X133 vccd1 _045_ a_6163_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X134 vccd1 _094_ a_7790_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X135 vssd1 _092_ a_7111_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X136 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_11251_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X137 vccd1 ctr\[1\] a_8101_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X138 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd _085_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X139 a_4364_6575# a_3965_6575# a_4238_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X140 a_5418_1653# a_5250_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X141 vccd1 net13 temp1.capload\[0\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X143 a_8285_2057# a_7295_1685# a_8159_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X144 a_12328_11471# a_12079_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X145 a_1665_5487# a_1499_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 a_5675_1679# a_4977_1685# a_5418_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X147 a_3153_6351# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X148 vssd1 a_8327_10357# ctr\[1\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R1 net14 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X149 vssd1 net12 a_3523_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X150 vccd1 _070_ a_7012_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X152 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_9034_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X153 a_10508_3311# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X155 a_2400_6575# a_1407_6575# a_2271_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X156 vccd1 net5 a_11159_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X157 io_out[4] a_2442_11180# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X158 vccd1 net11 a_3799_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X160 _026_ a_9319_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X161 vssd1 _048_ a_5904_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X162 a_1941_1501# a_1407_1135# a_1846_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X163 a_7741_2767# _020_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X164 a_7089_4399# a_6099_4399# a_6963_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X165 a_1855_11293# a_1407_10927# a_1761_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X166 a_5763_9867# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X167 vssd1 ctr\[7\] a_5169_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X169 a_7745_8323# _070_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X170 a_3061_9615# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X171 vssd1 a_4406_6687# a_4364_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X172 _076_ a_5283_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X173 vccd1 _005_ a_3309_11849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X174 a_4896_1135# _064_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X175 _091_ a_7203_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X177 vccd1 ctr\[3\] a_4165_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X178 a_9956_8527# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X179 a_3134_8207# a_2861_8213# a_3049_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X180 net7 a_10147_3863# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X181 vssd1 a_2014_1247# a_1972_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X182 vccd1 a_2442_10092# a_2355_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X184 vccd1 ctr\[2\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X185 vccd1 net12 a_2695_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X187 vccd1 a_3024_4373# _056_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X188 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10600_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X189 io_out[0] a_2442_6828# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X191 a_7012_10089# _082_ _042_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X192 a_3116_7637# _032_ a_3245_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X193 a_2400_10927# a_1407_10927# a_2271_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X195 a_2271_11293# a_1407_10927# a_2014_11063# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X196 _022_ a_3739_4193# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X197 io_out[5] a_2303_11703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X198 a_3516_5737# _051_ _012_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X200 a_8031_5737# _087_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
R2 temp1.dac.vdac_single.einvp_batch\[0\].vref_29.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X201 a_1573_7663# a_1407_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X202 vccd1 a_10924_8439# a_10875_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X204 a_5057_7439# ctr\[2\] a_4627_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X206 a_9033_9001# _080_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X207 ctr\[13\] a_8419_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 a_3481_4193# ctr\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X210 a_10049_5487# _091_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X211 a_2303_11703# a_2471_11703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X212 vssd1 _031_ a_4220_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X213 a_5911_9295# _040_ a_5693_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 vssd1 _054_ a_5363_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X215 a_3427_1385# _066_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X216 a_9955_4649# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
R3 vccd1 temp1.capload\[3\].cap_22.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X217 vccd1 a_6375_2883# _077_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X218 a_3153_4649# _021_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X219 vccd1 a_10239_5487# net5 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X220 vssd1 a_4319_11989# io_out[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X221 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10948_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X222 a_4897_3561# a_4709_3317# a_4815_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X223 a_2200_8207# _031_ a_1735_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X225 a_3247_6351# ctr\[6\] a_3153_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X226 vccd1 a_2014_11063# a_1948_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 a_10875_8207# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X229 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9864_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X230 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11980_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X231 a_4709_3317# _023_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X232 temp1.dac_vout_notouch_ net30 a_7820_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X233 vssd1 a_7131_4667# ctr\[4\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X234 a_2755_11689# net12 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 vssd1 a_6982_7093# a_6940_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X236 a_4153_6575# _012_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X237 a_8286_6031# a_8109_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X239 a_9660_10089# a_9411_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X241 vccd1 a_3302_8181# a_3229_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X242 a_10648_6263# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X243 a_1948_11293# a_1407_10927# a_1855_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X244 a_7461_10389# a_7295_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X245 a_3229_8207# a_2695_8213# a_3134_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X246 temp1.dac_vout_notouch_ net8 a_11980_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X247 vssd1 net11 a_3799_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X248 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_9034_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X250 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11612_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X251 ctr\[1\] a_8327_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 a_3155_9615# ctr\[5\] a_3061_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X253 a_5759_1679# a_4977_1685# a_5675_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X255 vccd1 _072_ a_6375_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X256 vssd1 temp1.dcdel_capnode_notouch_ a_5813_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X258 vssd1 a_7131_4667# a_7089_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X259 a_3233_5792# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
R4 temp1.capload\[4\].cap_23.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X260 a_10875_9839# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X261 a_3317_2057# a_2327_1685# a_3191_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X262 vccd1 _080_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X263 a_4747_6941# a_3965_6575# a_4663_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X264 a_2962_11748# a_2755_11689# a_3138_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X266 a_5829_5737# ctr\[9\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X267 a_7902_10357# a_7734_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X269 a_7820_9295# a_7571_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X270 vccd1 a_6395_1999# _067_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X271 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8951_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X272 vssd1 temp1.dcdel_capnode_notouch_ temp1.dcdel_out_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X275 a_5805_8751# a_5639_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X277 vssd1 net4 a_12079_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X278 a_2106_5599# a_1938_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X279 temp1.capload\[0\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X280 net4 a_10567_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X281 _045_ _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X282 a_8243_10383# a_7461_10389# a_8159_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X283 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9660_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X284 a_2355_1501# a_1573_1135# a_2271_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X285 a_2106_5599# a_1938_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X286 vssd1 a_1460_8725# net12 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X287 vssd1 a_2271_4765# a_2439_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X288 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9319_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X289 a_8114_5737# ctr\[4\] a_8031_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X290 a_6829_7663# _043_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X291 vssd1 _042_ a_7374_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X292 vccd1 net4 a_10975_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X293 vccd1 _027_ a_2939_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X294 _058_ a_2092_2883# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X295 vssd1 a_8327_10357# a_8285_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X296 vccd1 a_2442_10092# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X297 _082_ ctr\[1\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X298 a_7851_8323# _076_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X299 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd _026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X300 vccd1 net6 a_11987_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X302 a_10188_6263# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X303 ctr\[12\] a_8327_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X304 a_10785_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X305 a_5250_1679# a_4811_1685# a_5165_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X306 a_5819_4649# _040_ a_5601_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X307 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8031_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X308 vccd1 a_6429_6549# _010_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X310 temp1.capload\[1\].cap.Y net20 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X311 vssd1 a_5693_9269# _009_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X312 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12328_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X313 vssd1 _088_ a_8307_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X314 vccd1 _032_ a_7142_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X315 vccd1 a_4330_1135# a_4436_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X316 vssd1 net5 a_11159_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X319 vccd1 _096_ a_3153_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X320 vssd1 a_2563_10357# _031_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X321 a_2092_2883# _057_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X322 a_1761_6575# _000_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X323 vccd1 net6 a_11435_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X325 a_6982_7093# a_6814_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X327 a_7377_5059# _077_ a_7295_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X328 vssd1 a_8399_8215# _080_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 a_3689_10389# a_3523_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X330 a_4992_3561# _054_ a_4897_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X332 vssd1 net1 a_6375_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X333 vccd1 _090_ a_4365_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.105 ps=1.21 w=1 l=0.15
X334 _020_ a_7281_2528# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X335 temp_delay_last a_4555_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 vssd1 io_in[1] a_1407_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X339 a_5376_2057# a_4977_1685# a_5250_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X340 vssd1 a_4036_7093# _033_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X341 vccd1 _050_ a_3981_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X342 a_11796_7663# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X343 a_2014_7775# a_1846_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X344 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9411_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X345 a_2014_7775# a_1846_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X346 io_out[7] a_4319_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X347 a_8301_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X348 vssd1 a_4679_7637# _096_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X349 vccd1 _070_ a_4075_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X350 vssd1 _031_ a_2104_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X351 a_9660_10383# a_9411_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X352 a_9037_12015# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X354 a_3825_4193# ctr\[6\] a_3739_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X355 vccd1 temp1.dcdel_capnode_notouch_ temp1.capload\[2\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X356 a_4977_1685# a_4811_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X357 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10968_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X360 vssd1 _050_ a_4257_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X361 a_7381_5737# _076_ a_7285_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X363 a_2271_6941# a_1407_6575# a_2014_6711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X364 a_4036_7093# _032_ a_4165_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X365 vssd1 a_2303_11703# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X366 a_2865_2767# _016_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X367 vccd1 ctr\[9\] _059_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X368 vccd1 net11 a_7295_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X369 vccd1 a_8419_2741# a_8335_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X370 vssd1 a_3543_2741# a_3501_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X371 vccd1 _021_ a_4443_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X372 vssd1 temp_delay_last _027_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X374 vssd1 a_4555_10357# a_4513_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X375 a_7649_10383# _008_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X376 vssd1 temp1.dac.vdac_single.en_pupd a_7571_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
R5 vccd1 temp1.capload\[0\].cap_13.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X379 vccd1 a_7239_7119# a_7407_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X380 a_4165_7439# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X381 temp1.dac_vout_notouch_ net7 a_11888_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X382 vccd1 _080_ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X383 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9660_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X385 _077_ a_6375_2883# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X386 vssd1 a_2755_11689# a_2762_11593# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X387 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9411_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X388 a_5249_8585# a_4259_8213# a_5123_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X389 a_4404_9813# _040_ a_4796_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X390 a_2677_2773# a_2511_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X391 vssd1 _081_ a_8307_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X392 vssd1 net1 a_7387_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X393 a_4815_3561# _049_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_4982_1135# _063_ a_4896_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X396 vccd1 net12 a_7295_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X397 vccd1 _089_ a_9033_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X398 a_7348_8725# _093_ a_7477_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X399 vccd1 a_6963_4765# a_7131_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X401 vccd1 a_8159_10383# a_8327_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X402 vccd1 _045_ a_5065_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X403 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd _080_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X404 a_5613_3561# _049_ a_5541_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X405 a_4513_10761# a_3523_10389# a_4387_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X408 a_3131_7439# ctr\[7\] a_3035_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.107 ps=0.98 w=0.65 l=0.15
X409 a_11752_11703# net6 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X410 a_11776_10383# a_11527_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X411 a_6246_8863# a_6078_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X412 _023_ a_3983_3133# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X414 vccd1 net12 a_1407_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X415 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12328_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X416 _086_ ctr\[4\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X417 _069_ ctr\[12\] a_7102_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X418 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9955_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X419 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd a_10975_3863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X420 vccd1 ctr\[1\] a_6541_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X422 _045_ ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X423 a_8159_10383# a_7295_10389# a_7902_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X424 vssd1 _032_ a_4036_7637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X425 vccd1 _043_ a_5911_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X426 ctr\[11\] a_3359_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X427 vssd1 a_10975_3863# net3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 a_10047_7663# temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X429 vccd1 _045_ a_4985_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X430 _092_ a_5639_6397# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X431 vccd1 _093_ a_8951_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X432 temp1.dac_vout_notouch_ net7 a_10672_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X433 temp1.dac_vout_notouch_ net7 a_10580_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X435 vccd1 a_1735_9269# _003_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X436 a_11960_2767# a_11711_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X438 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11776_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X439 temp1.capload\[11\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X440 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11711_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X441 a_6645_6397# a_6375_6031# a_6541_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X442 _047_ ctr\[4\] a_5909_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X443 a_5415_7439# ctr\[3\] a_5057_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 _090_ ctr\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R6 vccd1 temp1.capload\[11\].cap_15.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X445 vccd1 _068_ a_7019_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X446 vccd1 net11 a_1407_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X447 vssd1 a_6963_4765# a_7131_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X448 _049_ ctr\[4\] a_5173_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 vccd1 _084_ _046_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X450 a_1952_10927# a_1573_10927# a_1855_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X451 vssd1 a_9319_2767# _026_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X452 a_10924_9991# net6 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X454 a_2271_8029# a_1407_7663# a_2014_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X455 vccd1 _079_ a_8399_8215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X456 vssd1 _072_ a_6375_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X457 a_10580_3561# a_10331_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X458 a_11704_6351# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X459 a_10672_2767# a_10423_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X460 a_4259_7439# ctr\[2\] a_4165_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X461 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8681_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X462 a_11868_5737# a_11619_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X466 vccd1 a_10648_6263# a_10599_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X467 a_3307_4087# ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X468 a_2014_11063# a_1855_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X469 vccd1 _050_ a_3516_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X471 a_6725_1679# ctr\[12\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X472 net3 a_10975_3863# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X474 vssd1 _084_ a_7663_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_6921_9839# a_6729_10144# _042_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X476 temp1.dac_vout_notouch_ net7 a_10120_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X477 vccd1 temp1.dcdel_out_n temp1.o_tempdelay vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X478 a_3685_8585# a_2695_8213# a_3559_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X479 vccd1 net11 a_2327_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X480 a_12163_4175# net7 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X482 a_3118_2741# a_2950_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X483 vccd1 a_2014_4511# a_1941_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X484 a_10004_4551# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X485 a_4215_5639# _050_ a_4613_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X486 a_8031_5737# _095_ a_8114_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X487 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd _026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X489 a_3118_2741# a_2950_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X490 a_4069_1999# a_3877_1740# _066_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X491 _027_ temp_delay_last vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X492 a_10120_3561# a_9871_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X493 a_4525_4399# _096_ a_4443_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X494 a_2104_9615# a_1878_9411# a_1735_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X495 a_11408_5737# a_11159_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X497 a_4897_3087# ctr\[8\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X498 a_6503_9117# a_5639_8751# a_6246_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X499 _032_ a_1959_1687# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X501 a_9037_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X502 vssd1 _076_ a_8307_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X503 vccd1 _024_ a_7019_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X504 a_5809_6397# ctr\[1\] a_5721_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X505 a_9344_6575# _085_ a_9224_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X506 _024_ a_4443_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X507 a_8569_6031# a_8392_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X508 vssd1 _026_ temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X509 _079_ a_7851_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X510 vccd1 a_3215_11989# io_out[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X511 vccd1 _032_ a_4533_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X512 vccd1 a_3375_2767# a_3543_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X513 vccd1 a_11752_4087# a_11703_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X514 ctr\[12\] a_8327_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X515 _052_ a_4215_5639# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.36 ps=2.72 w=1 l=0.15
X516 a_4789_6575# a_3799_6575# a_4663_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X517 a_6246_8863# a_6078_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X518 net8 a_11527_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X519 vccd1 net28 temp1.capload\[9\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X520 a_4259_3133# ctr\[11\] a_4153_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X521 vssd1 net11 a_1407_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_5515_10357# _028_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.28 ps=1.62 w=0.42 l=0.15
X523 a_3215_11989# in_measurement vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X524 vccd1 ctr\[11\] a_6625_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X525 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_11527_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X526 a_2397_1135# a_1407_1135# a_2271_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X527 vssd1 ctr\[5\] _088_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X530 a_11703_3855# net8 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X531 a_1878_9411# _036_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X532 a_3427_2473# _040_ a_3209_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X533 _025_ a_8859_2880# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X534 vccd1 a_2442_6828# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X535 vssd1 _054_ a_4815_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X536 a_6423_10615# ctr\[1\] a_6657_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X537 a_12212_4087# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X538 a_12072_8527# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X539 vccd1 _073_ _039_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X540 a_7203_5737# _077_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X541 a_3559_8207# a_2695_8213# a_3302_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X542 a_3209_1109# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X543 a_4627_7439# _070_ _045_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X544 vccd1 a_6671_9019# a_6587_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X545 vssd1 _076_ a_8307_7235# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X547 _042_ a_6729_10144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X548 vssd1 _029_ a_4404_9813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X549 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11803_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X550 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12236_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X551 a_9034_6575# ctr\[3\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X552 _084_ ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X553 vccd1 a_10004_4551# a_9955_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X555 a_10415_10703# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X557 _062_ ctr\[10\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X558 a_3739_4193# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X559 vssd1 a_7239_7119# a_7407_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X560 vssd1 a_1460_1653# net11 vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X561 a_1573_4399# a_1407_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X562 a_7461_10389# a_7295_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X563 a_1952_9839# a_1573_9839# a_1855_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X564 _060_ a_5363_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X565 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11980_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X566 vccd1 io_out[1] a_2200_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X567 a_5283_5737# ctr\[8\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X568 _094_ a_6541_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X569 vssd1 ctr\[2\] a_5864_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X570 a_12236_6825# a_11987_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X571 vssd1 _005_ a_3309_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X572 vccd1 ctr\[1\] a_5639_6397# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X573 _045_ ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X575 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd _089_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X576 temp1.dac_vout_notouch_ net8 a_10764_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X577 vssd1 a_4831_6843# a_4789_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X578 temp1.capload\[6\].cap.Y net25 a_5541_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 temp1.capload\[5\].cap.Y net24 a_10233_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X580 vccd1 a_3215_9813# _040_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X581 vssd1 a_6671_9019# ctr\[2\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X582 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11895_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X583 vssd1 a_2439_1403# a_2397_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X584 vssd1 a_2313_5175# _053_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X586 vccd1 a_3727_8181# a_3643_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X587 vccd1 net23 temp1.capload\[4\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X588 vccd1 ctr\[2\] a_5946_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X590 ctr\[11\] a_3359_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X591 a_10764_4649# a_10515_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X592 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8280_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X593 a_6477_1999# _065_ a_6395_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X594 ctr\[6\] a_2531_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X595 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_10239_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X596 a_9496_4175# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X597 a_8101_8323# _076_ a_8028_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X598 vssd1 a_2962_11748# a_2891_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X599 a_4425_8213# a_4259_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X600 a_6457_2883# ctr\[13\] a_6375_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X601 a_3375_2767# a_2677_2773# a_3118_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X602 vssd1 a_2934_1653# a_2892_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X603 vssd1 a_2442_6828# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X605 vssd1 _093_ a_9344_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X607 a_8859_2880# ctr\[13\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X608 a_2845_7119# net2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
R7 net21 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X609 a_5057_7439# ctr\[2\] a_4627_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X610 a_9033_9001# ctr\[5\] a_9233_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X614 a_3689_10389# a_3523_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X615 a_1757_2767# ctr\[8\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X616 _088_ ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X617 vssd1 _062_ a_4392_1795# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X618 vccd1 a_2442_11180# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X619 a_8280_4649# a_8031_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X620 vssd1 a_4404_9813# _006_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X621 a_3885_5737# ctr\[5\] _051_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X624 vssd1 _073_ a_7072_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X625 vccd1 _065_ a_3427_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X626 vssd1 _076_ a_7663_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X627 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9411_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X628 vssd1 net3 a_10791_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X629 a_5515_10357# _071_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X630 _063_ a_4392_1795# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X631 ctr\[0\] a_5291_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 ctr\[6\] a_2531_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 vssd1 net5 a_11987_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X634 vccd1 a_2007_5162# _013_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X635 vccd1 ctr\[2\] _043_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X637 a_3153_6031# _027_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X640 io_out[1] a_2439_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X641 _039_ _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X642 a_4982_1135# _040_ a_4813_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X644 vssd1 a_3852_4373# _061_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X645 temp1.dac_vout_notouch_ net8 a_12256_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X646 a_2355_11293# a_1573_10927# a_2271_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X647 net9 a_6191_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X648 io_out[5] a_2303_11703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X649 vccd1 a_2271_1501# a_2439_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X650 vssd1 a_2931_8903# _002_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X651 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9568_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X652 a_2014_4511# a_1846_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X653 a_7453_5737# _082_ a_7381_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X655 a_2014_4511# a_1846_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X656 _012_ a_3233_5792# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X657 temp1.dac_vout_notouch_ net7 a_11224_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X658 a_2681_1679# _018_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X659 a_4130_10357# a_3962_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X660 a_5165_1679# _017_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X661 vssd1 net12 a_7295_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X662 _040_ a_3215_9813# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X663 vccd1 _040_ a_3233_5792# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X664 vssd1 net6 a_11987_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X665 a_4153_6575# _012_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X666 a_8159_1679# a_7295_1685# a_7902_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X667 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9963_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X668 vssd1 net3 a_10331_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X669 a_10061_6825# _026_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X670 _040_ a_3215_9813# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X671 vccd1 _025_ a_9319_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X672 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8280_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X673 vssd1 a_2014_6711# a_1952_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X674 a_3981_4399# _022_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X676 vssd1 a_4130_10357# a_4088_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X677 a_9224_6575# _080_ a_9034_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X678 a_4387_10383# a_3689_10389# a_4130_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X680 a_11224_2767# a_10975_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X681 io_out[1] a_2439_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X682 io_out[7] a_4319_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X683 a_6963_4765# a_6099_4399# a_6706_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X684 a_6265_4399# a_6099_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X685 a_3459_2767# a_2677_2773# a_3375_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X686 a_7473_2223# _026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X687 vccd1 a_4831_6843# ctr\[5\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X688 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_10239_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X689 vccd1 net5 a_11619_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X690 a_10139_6351# temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X691 vccd1 net4 a_12079_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X692 net12 a_1460_8725# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X693 a_3245_7913# _027_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X694 vssd1 a_11251_9839# net6 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X695 a_8280_4943# a_8031_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X696 vccd1 net12 a_4259_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X697 a_11703_11791# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X698 vccd1 a_8327_10357# ctr\[1\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X699 net11 a_1460_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X700 a_4627_7439# _070_ _045_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X701 vssd1 _068_ a_7019_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X702 a_9773_5487# _087_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R8 net26 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X703 vssd1 a_2442_10092# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X704 a_4075_11471# _070_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X705 a_2931_8903# a_3074_8797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X706 io_out[4] a_2442_11180# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X707 vssd1 _031_ a_3300_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X708 temp1.capload\[12\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X709 temp1.capload\[3\].cap.Y net22 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X710 a_4859_8916# _041_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X711 _029_ a_5515_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
R9 vccd1 temp1.capload\[12\].cap_16.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X713 a_2104_9615# io_out[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X714 a_5363_3561# _059_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X715 a_10924_8439# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X716 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11704_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X719 net1 a_3834_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X720 _049_ ctr\[5\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X721 a_6732_6575# _045_ a_6429_6549# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X722 a_8951_7913# _095_ a_9034_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X723 io_out[4] a_2442_11180# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X725 vccd1 a_8327_1653# a_8243_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X726 a_1735_8181# a_1878_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X727 a_1761_6575# _000_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X729 a_2014_6711# a_1855_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X730 vssd1 ctr\[13\] _072_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X731 vccd1 a_8164_4087# a_8115_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X732 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12328_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X733 _045_ ctr\[3\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X735 a_12328_7913# a_12079_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
R10 vssd1 net23 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X736 temp1.capload\[14\].cap.Y net18 a_10785_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X737 vssd1 a_2271_1501# a_2439_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X739 ctr\[2\] a_6671_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X740 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9588_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X741 a_3994_10973# _038_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X743 vccd1 a_7407_7093# ctr\[3\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X744 _072_ ctr\[11\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X745 vssd1 net3 a_12163_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X746 vccd1 _084_ a_7913_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X747 vccd1 a_11251_9839# net6 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X748 vccd1 temp1.dcdel_capnode_notouch_ temp1.capload\[1\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X749 a_2271_11293# a_1573_10927# a_2014_11063# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X750 vccd1 a_11527_4943# net8 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X751 a_6817_6397# _071_ a_6717_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X752 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd _080_ a_9865_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X753 vccd1 _095_ a_8109_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X754 vssd1 net11 a_7295_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X755 a_4474_1795# _060_ a_4392_1795# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X756 _055_ a_6009_3317# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X757 a_4866_8181# a_4698_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X758 a_1855_10205# a_1573_9839# a_1761_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X761 vccd1 a_9233_8751# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X763 a_8115_3855# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X765 _072_ ctr\[12\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0894 ps=0.925 w=0.65 l=0.15
X766 _067_ _065_ a_6725_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X767 a_10705_5737# _026_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X768 a_11752_11703# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X769 a_3076_3145# a_2677_2773# a_2950_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X770 a_4330_1135# a_4153_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X771 a_10464_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X772 a_4624_9839# _039_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X773 net4 a_10567_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X774 a_4069_1999# _062_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X775 a_6729_7119# _010_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X776 temp1.dac_vout_notouch_ net7 a_11888_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X777 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9319_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X778 _069_ ctr\[13\] a_7019_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X779 a_2677_2773# a_2511_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X780 a_1938_5853# a_1499_5487# a_1853_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X782 temp1.capload\[13\].cap.Y net17 a_8301_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X783 a_7571_8751# _082_ a_7477_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X784 _050_ _049_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X785 a_11336_5487# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X786 a_2104_10703# io_out[4] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X787 a_11224_11177# a_10975_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X788 a_4859_8916# _041_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X789 vssd1 a_5601_4373# _011_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X791 a_2962_11748# a_2762_11593# a_3111_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X792 a_7203_5737# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X793 a_2289_3829# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X794 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9128_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X795 a_7209_8207# _076_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X796 a_9329_8751# _095_ a_9233_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.107 ps=0.98 w=0.65 l=0.15
X797 _045_ ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X798 a_1878_9411# _036_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X799 vssd1 _077_ _078_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X800 a_7994_2741# a_7826_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X801 vssd1 _060_ a_4985_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X802 vccd1 a_2439_4667# a_2355_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X803 a_9034_5737# _095_ a_9034_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X805 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9411_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X808 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8031_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X809 a_6423_10615# net9 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X811 vssd1 a_3375_2767# a_3543_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X812 vssd1 net4 a_10515_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X813 a_2313_5175# _032_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X814 temp1.dac_vout_notouch_ net8 a_11152_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X815 vccd1 ctr\[4\] a_3885_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X817 a_3138_11471# a_2891_11849# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X818 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11224_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X819 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9319_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X820 a_5415_7439# ctr\[1\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X821 vssd1 a_2007_5162# _013_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X823 a_1855_6941# a_1573_6575# a_1761_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X827 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_9034_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X828 _081_ ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X829 a_6541_7125# a_6375_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X830 vccd1 a_5675_1679# a_5843_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X831 ctr\[2\] a_6671_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 vssd1 ctr\[3\] _084_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X833 a_4971_7663# ctr\[3\] a_4875_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X834 vccd1 a_5324_7637# _070_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X835 a_1761_7663# _001_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X836 vssd1 net6 a_11703_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X837 a_10875_10089# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X838 a_3215_9813# _032_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X839 a_1573_9839# a_1407_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X840 _089_ a_8307_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X841 vccd1 ctr\[11\] a_3877_1740# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X843 a_1846_8029# a_1407_7663# a_1761_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X844 a_5065_3561# _049_ a_4992_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X845 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12072_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X846 vccd1 a_8251_2767# a_8419_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X847 vssd1 net5 a_11619_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X848 vccd1 temp1.dac_vout_notouch_ a_6559_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X849 vssd1 _051_ a_3425_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
R11 net13 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X850 vccd1 a_4555_10357# a_4471_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X852 vccd1 a_2271_6941# a_2442_6828# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X853 ctr\[0\] a_5291_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X854 vccd1 a_2932_9269# _036_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X855 vccd1 a_3359_1653# a_3275_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X856 vccd1 a_3209_1109# _018_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X857 net9 a_6191_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X858 a_7285_5737# _077_ a_7203_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X859 a_4165_7119# _027_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X860 vssd1 net29 a_12079_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X861 a_2563_10357# _030_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X862 vccd1 a_1735_7093# _000_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X863 vccd1 a_2289_3829# _014_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X864 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11684_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X865 a_4238_6941# a_3965_6575# a_4153_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X866 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12256_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X867 vccd1 a_10924_9991# a_10875_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X868 a_6814_7119# a_6375_7125# a_6729_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X869 vssd1 temp1.dcdel_capnode_notouch_ a_6457_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X870 vccd1 net11 a_1407_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X871 vssd1 a_3215_9813# _040_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X872 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_10140_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X873 vssd1 _024_ a_9013_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X874 _082_ ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X875 a_1665_3087# ctr\[8\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X877 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8115_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X879 a_1972_7663# a_1573_7663# a_1846_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X880 a_1761_9839# _003_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X881 vssd1 net11 a_2327_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X882 vccd1 net15 temp1.capload\[11\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X883 a_2271_10205# a_1573_9839# a_2014_9975# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X884 _087_ a_7295_5059# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X886 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd _026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X887 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11428_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X888 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_11059_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X889 net6 a_11251_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X890 a_11684_6825# a_11435_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X891 a_3427_2473# _061_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X892 a_7477_9001# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X893 a_5993_8751# _009_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X894 a_8251_2767# a_7387_2773# a_7994_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X896 vccd1 a_2271_10205# a_2442_10092# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X897 a_6940_7497# a_6541_7125# a_6814_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X898 a_3035_7439# _027_ a_2845_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X899 a_9779_8751# _080_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X900 vssd1 a_7994_2741# a_7952_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X901 _064_ _062_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 a_5794_10749# _028_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.175 ps=1.26 w=0.42 l=0.15
X905 a_10004_4551# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X906 a_8285_10761# a_7295_10389# a_8159_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X907 vssd1 _066_ a_3512_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X908 vssd1 net3 a_10975_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X909 a_6982_7093# a_6814_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X910 a_10255_9001# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X911 vssd1 _045_ a_6009_3317# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X912 vccd1 a_5283_5737# _076_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X913 vssd1 _046_ a_6732_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X914 a_4036_7637# _027_ a_4259_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
R12 vccd1 temp1.capload\[2\].cap_21.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X916 vccd1 ctr\[8\] a_1427_3087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X917 a_4443_4399# _096_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X918 a_7239_7119# a_6541_7125# a_6982_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X919 vssd1 a_1735_7093# _000_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X920 a_7826_2767# a_7387_2773# a_7741_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X921 a_11752_4087# net4 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X923 a_1853_5487# _013_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X925 vccd1 a_5418_1653# a_5345_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X926 a_8951_5737# _091_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X927 a_5541_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X928 vccd1 net6 a_12079_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X930 a_10233_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X931 vccd1 _080_ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X932 a_10875_10383# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X933 vccd1 a_4406_6687# a_4333_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X934 a_4451_9001# a_4259_8757# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X936 a_6091_3561# _054_ a_6009_3317# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X937 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd _083_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X938 a_8208_4399# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X939 a_3983_3133# ctr\[11\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X940 vccd1 _073_ a_4255_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X941 io_out[0] a_2442_6828# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X942 a_7851_8323# a_7745_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X943 vccd1 a_2014_1247# a_1941_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X944 _044_ a_5864_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X945 vssd1 a_2442_10092# a_2400_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X946 io_out[2] a_3727_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X947 vssd1 net2 a_3024_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X948 vssd1 ctr\[12\] a_6477_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X949 vssd1 a_9233_8751# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X950 a_5345_1679# a_4811_1685# a_5250_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X951 a_3965_6575# a_3799_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X952 vccd1 a_2442_6828# a_2355_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X953 a_7952_3145# a_7553_2773# a_7826_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X954 vccd1 a_2442_11180# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X955 a_11108_6727# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X956 a_3962_10383# a_3689_10389# a_3877_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X957 a_4333_6941# a_3799_6575# a_4238_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X958 a_2363_5853# a_1499_5487# a_2106_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X959 a_4675_11690# _074_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X960 vssd1 temp1.dcdel_capnode_notouch_ a_6089_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X961 vccd1 a_10924_10615# a_10875_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X962 a_6921_9839# _070_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X964 vccd1 net3 a_10791_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X965 vccd1 a_7072_10901# temp1.i_precharge_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X966 a_3302_8181# a_3134_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X967 vssd1 a_3215_11989# io_out[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X969 a_1573_1135# a_1407_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X970 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_10147_3863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X971 vssd1 _032_ a_2932_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X972 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9779_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X973 a_7841_6825# _076_ a_7745_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X975 vssd1 a_7407_7093# ctr\[3\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X976 vssd1 a_10147_3863# net7 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X977 a_10968_8751# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X979 a_4404_9813# temp_delay_last a_4624_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X980 a_1761_7663# _001_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X981 vssd1 a_3307_4087# _021_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X982 vssd1 _031_ a_2104_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X983 a_8113_12015# net20 temp1.capload\[1\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X984 a_1761_10927# _004_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X985 vccd1 a_5515_10357# _029_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.165 ps=1.33 w=1 l=0.15
X987 vssd1 _032_ a_7060_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X989 a_9034_5737# ctr\[6\] a_8951_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X991 a_11888_3087# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X993 a_7745_8323# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X994 a_6457_11791# net27 temp1.capload\[8\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X995 a_11061_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X996 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9687_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X997 vssd1 a_3302_8181# a_3260_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X999 a_3307_4087# ctr\[4\] a_3481_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1001 a_4065_3133# ctr\[9\] a_3983_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
R13 net30 vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1002 a_8307_9001# _077_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1003 vccd1 ctr\[7\] _054_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1004 vssd1 net3 a_11795_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1005 vccd1 net3 a_10331_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1006 a_7473_2223# a_7281_2528# _020_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1007 a_4815_3561# a_4709_3317# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X1008 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12256_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1009 vccd1 ctr\[0\] a_4679_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1010 _093_ a_7111_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1011 vssd1 a_7111_6031# _093_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1012 a_1460_1653# net1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1013 vccd1 a_8286_6031# a_8392_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1014 _065_ a_4815_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1015 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10875_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1016 ctr\[7\] a_2439_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1017 net7 a_10147_3863# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1018 a_3024_4373# ctr\[7\] a_3153_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1019 vccd1 a_2531_5755# a_2447_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1020 a_1846_8029# a_1573_7663# a_1761_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1021 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11868_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
R14 vccd1 temp1.capload\[7\].cap_26.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1023 a_6625_2883# ctr\[10\] a_6553_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1024 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_11527_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1025 _095_ a_7790_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1026 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_10061_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1027 a_5993_8751# _009_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1028 a_3965_6575# a_3799_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1029 a_3024_4373# ctr\[6\] a_3247_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1030 a_3852_4373# ctr\[9\] a_3981_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1031 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10875_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1032 vccd1 a_1427_3087# _057_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X1034 vccd1 net2 a_1959_1687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1035 vccd1 ctr\[7\] a_6375_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1036 _040_ a_3215_9813# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1037 vssd1 a_5675_1679# a_5843_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1039 _008_ a_7374_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X1040 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9588_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1041 a_1573_1135# a_1407_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1042 vssd1 a_2271_10205# a_2442_10092# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1043 vssd1 _029_ a_3131_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
R15 vccd1 temp1.capload\[14\].cap_18.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1045 a_6909_7119# a_6375_7125# a_6814_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1046 a_3852_4373# ctr\[8\] a_4075_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1047 ctr\[7\] a_2439_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1048 io_out[6] a_3215_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1049 vssd1 _077_ a_7851_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X1050 a_3049_8207# _002_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1051 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11408_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1052 a_8307_7235# _077_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1053 _071_ ctr\[9\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1054 a_6647_6825# _040_ a_6429_6549# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1055 vssd1 ctr\[1\] _082_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1056 a_3302_8181# a_3134_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1057 a_5693_9269# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1058 vccd1 a_3024_6005# _037_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1059 vssd1 net12 a_2695_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1060 a_11059_6825# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1061 vccd1 _093_ a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X1063 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10876_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1064 vccd1 net11 a_1499_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1065 a_6089_11791# net26 temp1.capload\[7\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1066 _038_ a_2845_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.112 ps=0.995 w=0.65 l=0.15
X1068 a_12256_7663# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1069 a_1855_10205# a_1407_9839# a_1761_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1070 temp1.dac_vout_notouch_ net30 a_7748_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1071 vccd1 net14 temp1.capload\[10\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1072 a_8304_5487# _080_ a_8114_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X1073 vssd1 _090_ a_4257_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1074 a_6423_10615# ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1076 temp1.dac_vout_notouch_ net7 a_10508_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1077 vccd1 _047_ a_5819_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1078 vssd1 _032_ a_2092_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1079 _085_ a_7663_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1082 a_6553_12015# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1083 vccd1 net10 a_6541_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1084 vssd1 net10 a_5915_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1085 a_3153_6031# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1086 a_7649_1679# _019_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1087 a_1941_8029# a_1407_7663# a_1846_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1088 vssd1 _094_ a_7790_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1089 vssd1 _073_ a_4617_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1090 _048_ _086_ a_6737_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1091 a_2713_11471# a_2303_11703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1092 a_6395_1999# _065_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X1093 _058_ a_2092_2883# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1094 vccd1 a_3559_8207# a_3727_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1095 io_out[6] a_3215_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1096 vccd1 _062_ a_4474_1795# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1100 vssd1 net6 a_10975_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1101 vssd1 ctr\[7\] a_3825_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd net5 a_10705_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1103 a_2355_6941# a_1573_6575# a_2271_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X1104 vccd1 ctr\[10\] a_3983_3133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1105 _041_ a_4451_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1106 vccd1 a_3116_7637# _035_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1108 temp1.dac_vout_notouch_ net7 a_10048_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1109 a_2950_2767# a_2677_2773# a_2865_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1110 io_out[3] a_2442_10092# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X1111 a_11704_10703# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1112 a_5169_4175# ctr\[6\] _054_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1114 a_10567_4917# temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1115 vccd1 _080_ a_8951_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X1117 a_4679_7637# ctr\[0\] a_5077_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1118 _019_ a_7019_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1119 a_6585_10749# net9 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1120 a_5639_6397# ctr\[7\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1122 io_out[2] a_3727_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1124 a_1573_9839# a_1407_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1125 vssd1 _045_ a_4815_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1126 a_4406_6687# a_4238_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1127 vssd1 a_4319_11989# io_out[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R16 vccd1 temp1.capload\[5\].cap_24.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1128 a_4406_6687# a_4238_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1129 a_9344_7663# _083_ a_9224_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X1130 a_5890_10749# net9 a_5794_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1131 _045_ ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X1132 ctr\[4\] a_7131_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1133 a_3245_7913# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1134 temp1.dac_vout_notouch_ net7 a_11040_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1135 a_2014_1247# a_1846_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1136 a_7663_6825# _077_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1137 a_8941_3133# ctr\[12\] a_8859_2880# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1138 a_2014_1247# a_1846_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1140 a_3851_11079# a_3994_10973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
R17 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd_30.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1141 vccd1 net12 a_5639_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1142 vssd1 _056_ a_2592_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1144 vssd1 net12 a_1407_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1145 vssd1 ctr\[4\] _086_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1146 io_out[7] a_4319_11989# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1147 a_8164_4087# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1148 vccd1 ctr\[6\] a_3153_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1149 a_10464_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1150 temp1.dac_vout_notouch_ net7 a_11960_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1151 vssd1 ctr\[12\] a_6375_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1152 vccd1 _081_ a_8557_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1154 a_11040_3561# a_10791_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1155 a_12164_6351# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
R18 net25 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1156 _077_ a_6375_2883# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X1157 net5 a_10239_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1158 vssd1 a_2442_11180# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X1159 vssd1 ctr\[6\] _090_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1160 vccd1 a_4319_11989# io_out[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1161 a_1846_4765# a_1407_4399# a_1761_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1162 vccd1 net16 temp1.capload\[12\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 vccd1 temp1.dcdel_capnode_notouch_ temp1.capload\[3\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1164 ctr\[4\] a_7131_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1165 a_10948_9295# a_10699_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1166 vssd1 net3 a_11711_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1167 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9588_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1168 a_6963_4765# a_6265_4399# a_6706_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1169 a_5415_7439# ctr\[3\] a_5057_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1170 a_2355_8029# a_1573_7663# a_2271_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1171 _071_ ctr\[8\] a_5829_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1172 vccd1 temp1.dcdel_capnode_notouch_ temp1.dcdel_out_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1173 a_7902_10357# a_7734_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1174 a_3209_2197# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1175 a_4259_8757# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X1176 a_10648_6263# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1178 a_7902_1653# a_7734_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1179 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8114_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X1180 _086_ ctr\[4\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1182 a_7019_2767# ctr\[12\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X1183 a_9034_7663# ctr\[2\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X1184 a_4679_7637# ctr\[1\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
R19 vccd1 temp1.capload\[15\].cap_19.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1185 a_10692_4175# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1186 vccd1 ctr\[4\] a_3307_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
R20 temp1.capload\[9\].cap_28.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1188 a_1731_2388# _058_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1190 vssd1 net3 a_10423_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1192 vccd1 a_10975_3863# net3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1193 a_4617_10927# _070_ _039_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1194 a_8159_10383# a_7461_10389# a_7902_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1195 vssd1 a_3215_9813# _040_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1196 a_1972_4399# a_1573_4399# a_1846_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1197 a_4215_5639# _090_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.365 ps=1.73 w=1 l=0.15
X1198 a_2174_2883# _057_ a_2092_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1200 vccd1 ctr\[4\] a_3245_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1201 temp1.capload\[14\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1203 a_6657_10749# _071_ a_6585_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1204 _062_ ctr\[10\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1205 vccd1 ctr\[4\] _047_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1206 _028_ a_5763_9867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1207 a_3061_9295# _027_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1208 a_5996_9615# _043_ a_5693_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1209 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11796_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1210 vssd1 _026_ temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1211 vssd1 _096_ a_3971_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1213 a_10096_7815# temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1214 vccd1 a_12212_4087# a_12163_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1215 vccd1 a_8159_1679# a_8327_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1216 a_10188_6263# temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1218 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11704_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1219 a_9785_7913# temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1221 a_2563_10357# _030_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1222 vssd1 a_7407_7093# a_7365_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1223 vccd1 a_8399_8215# _080_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1224 vssd1 ctr\[2\] _081_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1225 a_6587_9117# a_5805_8751# a_6503_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1226 a_10599_6351# temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X1227 a_8307_9001# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1228 a_6736_10927# temp1.dac_vout_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1229 vccd1 a_4036_7093# _033_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1230 a_6163_3561# _049_ a_6091_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1233 vccd1 a_6423_10615# _073_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1234 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_9034_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X1235 temp1.capload\[13\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1236 vccd1 net12 a_1407_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1237 _008_ a_7374_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1238 a_11844_2375# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1239 a_5819_4649# _048_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1240 vccd1 a_2962_11748# a_2891_11849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1241 ctr\[9\] a_3543_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1242 vccd1 a_5363_3561# _060_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1244 a_12163_3855# net7 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1245 _080_ a_8399_8215# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1246 a_9861_11791# net21 temp1.capload\[2\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1247 a_9496_5263# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1248 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10255_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1250 vssd1 a_11527_4943# net8 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1251 vssd1 _093_ a_9344_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X1252 _076_ a_5283_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X1254 a_6461_8527# _028_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1256 a_5801_2057# a_4811_1685# a_5675_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1257 vssd1 _086_ a_7295_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1258 vccd1 net5 a_11527_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1260 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11336_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1263 vccd1 a_2439_1403# a_2355_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1264 a_4165_7119# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1266 a_8208_5263# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1267 a_4257_5487# a_4215_5639# _052_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X1268 vccd1 a_7348_8725# temp1.dac.vdac_single.en_pupd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1269 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_10672_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1270 _070_ a_5324_7637# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1272 _059_ ctr\[8\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1274 a_11152_3087# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1276 io_out[0] a_2442_6828# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X1277 a_7741_2767# _020_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1278 vccd1 a_3851_11079# _005_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X1280 vssd1 a_8419_2741# a_8377_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1281 vssd1 a_4866_8181# a_4824_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1282 vccd1 a_2939_10615# _030_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1283 vssd1 a_3559_8207# a_3727_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1284 io_out[4] a_2442_11180# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X1285 vccd1 _060_ a_3427_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1287 vssd1 net5 a_11159_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1288 _074_ a_4255_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X1289 a_2934_1653# a_2766_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1290 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd _091_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1291 a_2271_10205# a_1407_9839# a_2014_9975# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1292 a_7734_1679# a_7295_1685# a_7649_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1294 vssd1 a_4036_7637# _034_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X1295 a_1761_4399# _014_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1296 a_2939_7119# ctr\[7\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1297 vccd1 net9 a_5515_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1298 a_8307_7235# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1299 a_10672_7913# a_10423_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1300 a_3512_1135# _065_ a_3209_1109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1301 a_7553_2773# a_7387_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1302 a_7477_9001# _078_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1303 a_12236_10383# a_11987_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1304 a_12256_10927# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1305 a_6633_1999# _065_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1306 vccd1 ctr\[10\] _062_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1307 vssd1 io_in[0] a_3834_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1308 vccd1 ctr\[7\] a_3739_4193# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1309 vccd1 ctr\[1\] _082_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1310 a_6717_6397# ctr\[1\] a_6645_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X1311 a_9233_8751# _080_ a_9117_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.14 ps=1.08 w=0.65 l=0.15
X1312 a_6538_4765# a_6099_4399# a_6453_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1314 a_11796_5487# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1315 vccd1 _075_ a_7201_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1316 vssd1 _040_ a_4982_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X1317 _092_ a_5639_6397# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
R21 vccd1 temp1.capload\[13\].cap_17.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1319 vssd1 a_2014_11063# a_1952_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X1320 vssd1 ctr\[9\] a_5283_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X1321 a_7860_2057# a_7461_1685# a_7734_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1322 a_4875_7663# ctr\[1\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X1323 a_4165_7663# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X1325 vccd1 a_2014_9975# a_1948_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X1326 a_9033_9001# _093_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1328 temp1.dac_vout_notouch_ net8 a_12052_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1329 a_2271_4765# a_1407_4399# a_2014_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1330 vccd1 ctr\[3\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1331 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10791_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1332 vccd1 _089_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1333 vccd1 a_3191_1679# a_3359_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1334 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12236_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1335 a_7902_1653# a_7734_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1336 vssd1 a_4831_6843# ctr\[5\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1337 a_8485_7235# _076_ a_8389_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1338 a_1853_5487# _013_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1340 a_9224_7663# _080_ a_9034_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
R22 net20 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1343 a_1948_10205# a_1407_9839# a_1855_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X1344 a_8159_1679# a_7461_1685# a_7902_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1345 a_6664_4399# a_6265_4399# a_6538_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1346 vccd1 ctr\[2\] a_4165_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1347 a_5909_4175# _096_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1348 vccd1 a_8327_10357# a_8243_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1349 a_4613_8207# _007_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1351 vssd1 net1 a_4153_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1352 vccd1 a_3118_2741# a_3045_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1353 _046_ _043_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1354 a_12052_4649# a_11803_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1355 _026_ a_9319_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
R23 net27 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1358 a_5911_9295# _044_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1359 a_10096_7815# temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1361 vccd1 a_2531_5755# ctr\[6\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1362 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11152_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1363 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10699_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1364 a_9773_6575# _085_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1367 a_11108_6727# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1368 vssd1 net5 a_11987_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1369 vssd1 net3 a_11251_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1370 vssd1 a_6706_4511# a_6664_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1371 a_4627_7439# ctr\[2\] a_5057_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1372 a_3045_2767# a_2511_2773# a_2950_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1373 vccd1 ctr\[3\] a_4679_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1374 a_1731_2388# _058_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1375 a_3191_1679# a_2327_1685# a_2934_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1376 vssd1 net4 a_11803_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1377 _066_ a_3877_1740# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X1378 vccd1 _040_ a_7281_2528# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X1379 a_7565_12015# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1380 a_4796_10089# _029_ a_4541_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1381 a_9936_9295# a_9687_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1382 a_2476_5059# _032_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X1383 vccd1 _071_ a_6423_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1384 a_5996_10749# _071_ a_5890_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X1387 vccd1 a_2313_5175# _053_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X1388 temp1.capload\[9\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1389 vccd1 a_2442_11180# a_2355_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X1390 net1 a_3834_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1391 a_11888_3311# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1393 _017_ a_4982_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1394 _091_ a_7203_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1395 a_10924_8439# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1397 a_2766_1679# a_2327_1685# a_2681_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1398 vssd1 net4 a_10515_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1399 a_4259_7663# ctr\[3\] a_4165_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1400 a_7994_2741# a_7826_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1401 _079_ a_7851_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1402 vccd1 a_4679_7637# _096_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X1403 vccd1 _088_ a_8557_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1405 a_5415_7439# ctr\[1\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1406 vccd1 a_2439_7931# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1407 vssd1 a_3024_4373# _056_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X1408 a_4319_11989# temp1.o_tempdelay vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1409 vssd1 _032_ a_3116_7637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X1410 vssd1 temp1.dcdel_capnode_notouch_ a_8113_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1411 a_9955_10383# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1412 a_7201_11177# _078_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1413 _019_ a_7019_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1414 a_10924_9991# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1416 a_2363_5853# a_1665_5487# a_2106_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1417 _055_ a_6009_3317# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1418 a_8424_5487# _087_ a_8304_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X1419 vssd1 ctr\[1\] a_5849_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1420 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8031_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1421 temp1.capload\[15\].cap.Y net19 a_11061_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1422 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9956_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1423 a_2892_2057# a_2493_1685# a_2766_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1424 vssd1 a_8159_1679# a_8327_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1426 a_4330_1135# a_4153_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1427 a_2200_9295# _031_ a_1735_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1428 a_4675_11690# _074_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1429 a_2400_9839# a_1407_9839# a_2271_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X1430 vssd1 _073_ a_4345_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1431 a_11428_3311# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1432 vssd1 _076_ a_7295_5059# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1433 vccd1 net5 a_12079_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1434 a_6453_4399# _011_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1435 a_9955_4399# temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X1436 a_5250_1679# a_4977_1685# a_5165_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1437 net2 a_1407_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1438 a_3153_4399# _021_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X1439 _088_ ctr\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1441 a_6737_5263# _045_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1442 vssd1 a_10239_5487# net5 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1443 a_9034_6825# _095_ a_9034_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X1444 a_7734_10383# a_7461_10389# a_7649_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1445 a_11980_9615# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1446 vccd1 net11 a_4811_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1447 a_7745_6825# _077_ a_7663_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1448 vccd1 _070_ _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
R24 net22 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1449 a_12164_6575# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1450 a_4866_8181# a_4698_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1452 vssd1 a_2439_7931# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1455 vssd1 a_7902_10357# a_7860_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1457 vccd1 _082_ a_7205_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1458 a_2104_7439# a_1878_7235# a_1735_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1459 a_7734_10383# a_7295_10389# a_7649_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1460 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_10791_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1461 a_11980_4399# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1462 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12164_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1463 vccd1 a_1460_8725# net12 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1464 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_9034_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X1466 a_1509_3087# _055_ a_1427_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1467 io_out[3] a_2442_10092# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X1469 vccd1 a_1460_1653# net11 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1470 vccd1 a_4663_6941# a_4831_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1471 _045_ _070_ a_4627_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1472 a_4036_7637# _032_ a_4165_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1473 vssd1 _093_ a_7348_8725# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X1474 a_9117_8751# _089_ a_9033_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X1475 vccd1 a_2931_8903# _002_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X1476 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd _080_ a_9773_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1477 a_2271_8029# a_1573_7663# a_2014_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1478 a_10047_7913# temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1479 a_1948_6941# a_1407_6575# a_1855_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
R25 net15 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1480 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd _080_ a_9779_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1481 vccd1 a_3215_9813# _040_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1483 vssd1 a_2442_11180# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X1484 a_10692_4399# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
R26 vssd1 net28 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1485 temp_delay_last a_4555_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1486 vssd1 a_1959_1687# _032_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1488 vssd1 net11 a_1407_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1489 a_8114_5487# ctr\[4\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X1490 _090_ ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1491 vccd1 a_3209_2197# _016_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1492 a_4255_11471# a_4075_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1493 vccd1 ctr\[4\] _049_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1494 vssd1 a_7072_10901# temp1.i_precharge_n vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X1495 vccd1 a_1735_8181# _001_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X1496 temp1.dac_vout_notouch_ net8 a_10692_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1497 vccd1 _092_ a_7111_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1499 _083_ a_8307_7235# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1500 vccd1 net25 temp1.capload\[6\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1501 vssd1 net6 a_11435_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1502 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9496_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1503 vccd1 _039_ a_4541_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1504 _068_ a_7060_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1505 vccd1 net24 temp1.capload\[5\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1506 vssd1 a_3209_1109# _018_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1507 vssd1 a_4675_11690# in_measurement vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1508 ctr\[8\] a_2439_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1509 a_1878_7235# _033_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1510 a_5601_4373# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1511 vssd1 a_4663_6941# a_4831_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1512 a_8761_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1514 vssd1 ctr\[10\] _072_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.0878 ps=0.92 w=0.65 l=0.15
X1515 a_1938_5853# a_1665_5487# a_1853_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1516 vssd1 a_6429_6549# _010_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1517 vccd1 net29 a_12079_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1518 a_3247_4399# _096_ a_3153_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1520 a_4160_1679# _060_ _066_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1521 a_5864_8323# _028_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1522 _057_ _055_ a_1757_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X1523 temp1.capload\[0\].cap.Y net13 a_10509_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1524 a_2865_2767# _016_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1525 vccd1 a_9319_2767# _026_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1527 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11040_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1528 a_2939_7119# net2 a_2845_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X1529 temp1.capload\[11\].cap.Y net15 a_6553_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1530 a_3962_10383# a_3523_10389# a_3877_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1531 a_6503_9117# a_5805_8751# a_6246_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1532 vccd1 ctr\[8\] a_3983_3133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1533 vccd1 a_7131_4667# a_7047_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1534 _045_ ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1535 vccd1 a_2271_11293# a_2442_11180# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X1536 vccd1 _032_ a_2174_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1539 a_4075_4399# _050_ a_3981_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1540 vssd1 _061_ a_3512_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1541 a_3074_8797# _035_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X1543 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd a_10975_3863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1544 a_4679_7637# ctr\[2\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1545 a_8251_2767# a_7553_2773# a_7994_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1546 a_6814_7119# a_6541_7125# a_6729_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1547 a_3994_10973# _038_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1548 _029_ a_5515_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X1549 _072_ ctr\[13\] a_6095_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.13 ps=1.26 w=1 l=0.15
X1551 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd _026_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1552 a_4985_2223# _062_ _064_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1553 a_9233_8751# _095_ a_9033_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1554 a_11844_2375# net3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1555 vssd1 _090_ a_7203_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1557 a_11040_9001# a_10791_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1558 vssd1 a_1735_8181# _001_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1559 a_2861_8213# a_2695_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1560 vssd1 _093_ a_8424_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X1561 a_8951_6825# _085_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X1562 a_1735_10357# a_1878_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1563 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11803_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1564 a_5905_2767# ctr\[11\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1566 _024_ a_4443_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1567 net10 a_6375_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1568 vssd1 net12 a_4259_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1569 vssd1 ctr\[11\] a_6375_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1570 a_2592_4175# _055_ a_2289_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1571 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd _026_ a_9785_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1572 a_7201_11177# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1573 a_5363_3561# _049_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1574 vccd1 ctr\[12\] a_8859_2880# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1575 ctr\[9\] a_3543_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1576 vccd1 net12 _075_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1578 a_4627_7439# ctr\[2\] a_5057_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1579 vccd1 temp1.dac.vdac_single.en_pupd a_7571_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1580 vssd1 net5 a_12079_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1581 vccd1 _045_ a_5613_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1582 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd _080_ a_10049_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1583 a_1761_9839# _003_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1584 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11888_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
R27 net18 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1585 a_4613_1135# a_4436_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1586 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref a_11251_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1589 a_5915_6397# _071_ a_5809_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1590 ctr\[10\] a_5843_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1591 a_8485_9001# _076_ a_8389_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1592 a_1952_6575# a_1573_6575# a_1855_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X1595 a_2064_5487# a_1665_5487# a_1938_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1596 a_10600_3087# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1597 a_4985_4943# _049_ _050_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1598 vccd1 a_2271_8029# a_2439_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1599 vccd1 net11 a_6099_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1601 a_2507_3855# _040_ a_2289_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1602 vccd1 a_5123_8207# a_5291_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1603 a_1665_3087# _055_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1606 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9411_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1607 vccd1 a_6982_7093# a_6909_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1609 vssd1 _031_ a_2104_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1610 vssd1 a_4387_10383# a_4555_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1611 a_10875_8527# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
R28 net17 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1612 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11803_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1613 vssd1 a_2106_5599# a_2064_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1614 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9779_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1615 a_10567_4917# temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1616 a_8286_6031# a_8109_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1617 a_5123_8207# a_4259_8213# a_4866_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1618 vccd1 a_11108_6727# a_11059_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1619 a_9034_6825# ctr\[3\] a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1620 a_10139_6031# temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1621 net2 a_1407_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1622 a_11703_11471# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
R29 vccd1 temp1.capload\[1\].cap_20.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1623 vccd1 a_10567_4917# net4 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1624 vccd1 _070_ _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1625 _046_ _084_ a_6829_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1626 vccd1 a_4130_10357# a_4057_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1627 vccd1 net5 a_12079_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1630 vccd1 a_10004_10615# a_9955_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1631 a_3559_8207# a_2861_8213# a_3302_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1632 a_12212_4087# net3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1633 a_9588_10703# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1634 a_8335_2767# a_7553_2773# a_8251_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1635 vssd1 ctr\[1\] a_7851_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1636 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1637 net6 a_11251_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1638 a_10509_11791# temp1.dcdel_capnode_notouch_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1639 _045_ _070_ a_4627_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1640 a_2014_11063# a_1855_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X1641 a_3061_9295# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1642 a_1846_1501# a_1407_1135# a_1761_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1643 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11776_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1645 vccd1 net10 a_6191_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1647 vccd1 a_11752_11703# a_11703_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1648 vccd1 _026_ a_10255_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1649 a_11960_3561# a_11711_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1650 vccd1 net6 a_11527_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1651 _065_ a_4815_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X1653 a_6729_10144# _032_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1654 a_8557_7235# _082_ a_8485_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1655 a_6375_2883# ctr\[13\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1656 vssd1 _054_ a_6009_3317# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1657 vssd1 a_2932_9269# _036_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X1658 a_6078_9117# a_5639_8751# a_5993_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1659 vccd1 net18 temp1.capload\[14\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1660 vssd1 a_2014_7775# a_1972_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1661 temp1.dac_vout_notouch_ net7 a_11500_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1663 a_6541_7125# a_6375_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1664 a_10876_9615# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1665 vssd1 _089_ a_9779_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1668 a_11776_6031# a_11527_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1669 vssd1 _032_ a_4451_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1670 vccd1 _080_ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1672 vccd1 net3 a_11251_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1673 vssd1 a_8327_1653# a_8285_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1674 a_1972_1135# a_1573_1135# a_1846_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1675 vccd1 a_5291_8181# a_5207_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1676 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_11435_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1677 vccd1 a_2442_6828# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X1678 vccd1 a_3727_8181# io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1679 _075_ net12 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1680 vccd1 a_11844_2375# a_11795_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X1682 vccd1 a_1735_10357# _004_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X1683 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11803_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1684 vssd1 net11 a_1499_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1685 a_7142_1385# _067_ a_7060_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1686 vssd1 _082_ a_6921_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X1687 a_6204_8751# a_5805_8751# a_6078_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1688 a_11500_3561# a_11251_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1689 _022_ a_3739_4193# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1690 vssd1 _095_ a_8109_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1691 a_4220_10927# a_3994_10973# a_3851_11079# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1692 a_10924_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1693 a_7461_1685# a_7295_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1694 a_2447_5853# a_1665_5487# a_2363_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1695 vccd1 net17 temp1.capload\[13\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1696 vccd1 _093_ a_8951_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X1697 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_9936_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1698 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12052_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1699 ctr\[3\] a_7407_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1700 vssd1 temp1.dcdel_capnode_notouch_ a_9861_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1701 a_3501_3145# a_2511_2773# a_3375_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1702 vssd1 a_2442_11180# a_2400_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X1704 vccd1 a_4859_8916# _007_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1705 a_3049_8207# _002_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1706 a_11795_2473# net7 temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X1707 _078_ _077_ a_7209_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1708 a_2313_5175# _052_ a_2476_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1709 vssd1 _032_ a_4036_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X1711 vssd1 a_6375_2883# _077_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X1712 a_2104_7439# io_out[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1713 a_7933_8323# a_7745_8323# a_7851_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1714 a_7553_2773# a_7387_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1715 vccd1 ctr\[5\] a_3061_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1717 vssd1 a_6246_8863# a_6204_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1718 net10 a_6375_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1719 temp1.capload\[10\].cap.Y net14 a_9037_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1720 a_8951_5737# _095_ a_9034_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X1721 vccd1 net5 a_11159_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1722 a_11868_7913# a_11619_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1723 a_12052_9295# a_11803_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1724 a_7323_7119# a_6541_7125# a_7239_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1725 vccd1 ctr\[1\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 _078_ _076_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1727 a_1761_4399# _014_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1729 a_10875_10703# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X1730 temp1.dac_vout_notouch_ net8 a_12328_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1731 a_9568_3855# a_9319_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1732 vccd1 a_3852_4373# _061_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1733 a_1573_7663# a_1407_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1735 a_12328_5737# a_12079_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1736 vssd1 a_2442_6828# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X1737 a_3877_10383# _006_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1739 vssd1 a_3851_11079# _005_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1741 a_1573_10927# a_1407_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1742 vssd1 a_8251_2767# a_8419_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1743 a_4088_10761# a_3689_10389# a_3962_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1744 temp1.dcdel_capnode_notouch_ temp1.i_precharge_n a_6808_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1745 vccd1 io_in[0] a_3834_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1746 vccd1 _062_ a_4160_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X1747 a_3111_11837# a_2891_11849# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1748 a_2355_10205# a_1573_9839# a_2271_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X1750 vccd1 a_2014_6711# a_1948_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X1752 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12052_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1753 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12144_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1756 vccd1 a_10147_3863# net7 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1757 vccd1 net1 a_6375_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1758 _031_ a_2563_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1759 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12164_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1761 _084_ ctr\[3\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1762 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12256_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1763 vccd1 io_out[3] a_2200_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X1764 vccd1 a_3307_4087# _021_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1765 a_11612_6575# temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1766 a_3309_11849# a_2762_11593# a_2962_11748# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1767 a_3981_4649# _022_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1768 vssd1 net12 a_1407_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1769 a_5541_3561# _054_ a_5445_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1770 vccd1 _080_ a_8951_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X1771 vssd1 ctr\[1\] a_5415_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1773 a_4613_4399# _021_ a_4525_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1774 vccd1 a_5693_9269# _009_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1775 a_1573_6575# a_1407_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1776 a_11408_7913# a_11159_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1777 a_1761_1135# _015_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1778 vccd1 temp1.dcdel_capnode_notouch_ temp1.capload\[8\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1779 a_11980_8751# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1781 vssd1 _023_ a_4719_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1782 a_1573_10927# a_1407_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1784 vssd1 a_4859_8916# _007_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1785 a_12052_9001# a_11803_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1786 a_12144_8207# a_11895_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1787 vccd1 temp1.o_tempdelay a_5515_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0746 ps=0.775 w=0.42 l=0.15
X1788 a_2681_1679# _018_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1789 a_4709_3317# _023_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1790 vssd1 a_3359_1653# a_3317_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1792 ctr\[10\] a_5843_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1793 a_8028_8323# _077_ a_7933_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X1794 vccd1 net1 a_4153_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1795 a_3113_10721# _029_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1796 a_5675_1679# a_4811_1685# a_5418_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1797 a_1878_7235# _033_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X1798 vssd1 a_5515_10357# _029_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.107 ps=0.98 w=0.65 l=0.15
X1799 temp1.dac_vout_notouch_ net8 a_10692_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
R30 net16 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1800 a_4404_9813# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X1801 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd _087_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1802 a_4663_6941# a_3799_6575# a_4406_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1803 vssd1 a_5418_1653# a_5376_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1804 vssd1 a_5123_8207# a_5291_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1805 a_2200_10383# _031_ a_1735_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1806 vssd1 net12 a_5639_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1807 a_2493_1685# a_2327_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1808 temp1.dac_vout_notouch_ net7 a_10968_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1809 vccd1 _027_ a_2939_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1811 a_2271_1501# a_1407_1135# a_2014_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1812 vccd1 net5 a_11987_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1814 net12 a_1460_8725# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1815 io_out[3] a_2442_10092# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1816 vccd1 _064_ a_4813_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1818 vccd1 _045_ a_6647_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1819 vccd1 _032_ a_6729_10144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X1820 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8208_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1821 vccd1 temp_delay_last _027_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1822 vccd1 net4 a_11803_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1823 a_3300_8751# a_3074_8797# a_2931_8903# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1824 a_2271_4765# a_1573_4399# a_2014_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1825 a_8114_5737# _095_ a_8114_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X1826 a_1665_5487# a_1499_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1828 vssd1 temp1.dcdel_out_n temp1.o_tempdelay vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1829 temp1.capload\[6\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1831 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9660_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1832 temp1.capload\[5\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1833 vssd1 net5 a_11619_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1834 a_6078_9117# a_5805_8751# a_5993_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1835 _059_ ctr\[9\] a_4897_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1836 a_3877_1740# ctr\[11\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1839 vssd1 net10 a_6191_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1840 vccd1 a_2014_7775# a_1941_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1841 vccd1 net4 a_10515_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1842 vssd1 a_3215_11989# io_out[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1843 a_1427_3087# _055_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X1844 a_8389_7235# _077_ a_8307_7235# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1846 temp1.capload\[12\].cap.Y net16 a_7565_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1847 _051_ ctr\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1848 a_3309_11849# a_2755_11689# a_2962_11748# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1849 vccd1 a_5843_1653# a_5759_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1850 a_3024_6005# net2 a_3153_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1851 vccd1 ctr\[12\] a_6395_1999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
R31 vccd1 temp1.capload\[8\].cap_27.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1853 a_7734_1679# a_7461_1685# a_7649_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1854 vssd1 a_1735_10357# _004_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1855 _032_ a_1959_1687# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1856 a_7913_6825# _082_ a_7841_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1857 vccd1 a_4831_6843# a_4747_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1858 a_9660_4649# a_9411_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1860 a_8569_6031# a_8392_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1861 a_1573_6575# a_1407_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1862 vccd1 temp1.dcdel_capnode_notouch_ temp1.capload\[7\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1863 a_5165_1679# _017_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1865 vccd1 _090_ a_7453_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1867 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8031_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1868 vccd1 a_5601_4373# _011_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1871 vssd1 net12 a_1407_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1872 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_9233_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.21 ps=1.29 w=0.65 l=0.15
X1873 vssd1 net11 a_4811_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1874 vssd1 _025_ a_9319_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1875 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_9200_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1876 a_7295_10927# _075_ a_7201_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1877 temp1.capload\[9\].cap.Y net28 a_9037_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1878 _023_ a_3983_3133# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1879 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd a_10047_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1880 vssd1 a_2442_10092# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X1882 a_6453_4399# _011_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1884 a_2200_7119# _031_ a_1735_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1885 a_10004_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X1886 a_4533_9001# a_4259_8757# a_4451_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1889 a_7748_9615# temp1.dac.vdac_single.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1890 a_9864_9615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1891 vccd1 net11 a_1407_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1892 a_3425_5487# a_3233_5792# _012_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1893 temp1.dac_vout_notouch_ net8 a_11224_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1894 vssd1 a_5291_8181# a_5249_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1895 vccd1 a_3215_11989# io_out[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1896 vssd1 a_3727_8181# io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1897 vccd1 _086_ _048_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1898 vccd1 a_6246_8863# a_6173_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1899 a_3643_8207# a_2861_8213# a_3559_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1900 vccd1 io_out[4] a_2200_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X1901 a_2271_6941# a_1573_6575# a_2014_6711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X1902 temp1.dac_vout_notouch_ net7 a_10600_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1904 a_9200_4649# a_8951_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1905 temp1.capload\[15\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1907 temp1.capload\[8\].cap.Y net27 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1909 vccd1 net11 a_2511_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1910 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_9034_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X1911 vccd1 a_7131_4667# ctr\[4\] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1912 vccd1 net12 a_1407_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1915 vccd1 ctr\[3\] _084_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1917 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12328_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1918 a_6095_2767# ctr\[12\] a_5989_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.19 ps=1.38 w=1 l=0.15
X1919 a_1846_4765# a_1573_4399# a_1761_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1920 a_12328_7119# a_12079_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1921 ctr\[3\] a_7407_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1922 vccd1 a_7902_1653# a_7829_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1923 vssd1 net3 a_11711_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1924 a_5805_8751# a_5639_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1926 a_11224_4649# a_10975_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1927 a_3396_9001# _031_ a_2931_8903# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1928 a_8557_9001# _082_ a_8485_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1930 a_6173_9117# a_5639_8751# a_6078_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1931 a_7829_1679# a_7295_1685# a_7734_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1932 vccd1 net4 a_10515_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1933 vssd1 a_5363_3561# _060_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X1934 _054_ ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1935 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd a_9319_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1936 a_6375_2883# ctr\[10\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1937 a_3116_7637# _027_ a_3339_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1938 a_7060_1385# _067_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1939 _095_ a_7790_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1940 _093_ a_7111_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1941 vccd1 _086_ a_7545_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1943 a_10048_3311# net3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X1944 a_2007_5162# _053_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1945 net3 a_10975_3863# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1946 vssd1 a_8286_6031# a_8392_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1947 vccd1 a_2271_4765# a_2439_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1948 a_2489_5487# a_1499_5487# a_2363_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1951 vssd1 net6 a_10875_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1952 _027_ temp_delay_last vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1953 _094_ a_6541_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X1954 a_1735_9269# a_1878_9411# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1955 a_7860_10761# a_7461_10389# a_7734_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1956 a_7295_5059# _077_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1957 a_5057_7439# ctr\[3\] a_5415_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1958 a_5173_4399# ctr\[5\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1959 vccd1 _029_ a_2939_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X1960 vssd1 a_2442_6828# a_2400_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X1961 vssd1 a_2014_9975# a_1952_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X1962 a_2507_3855# _056_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1963 a_3512_2223# _060_ a_3209_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1964 vccd1 ctr\[4\] _086_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1965 a_2766_1679# a_2493_1685# a_2681_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1966 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12256_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X1968 vssd1 ctr\[7\] a_6375_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1969 temp1.capload\[10\].cap.Y temp1.dcdel_capnode_notouch_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1970 a_1855_11293# a_1573_10927# a_1761_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X1971 vssd1 ctr\[5\] a_9329_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.29 as=0.115 ps=1 w=0.65 l=0.15
X1972 vssd1 net11 a_1407_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R32 vccd1 temp1.capload\[10\].cap_14.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1973 a_4316_11177# _031_ a_3851_11079# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1974 vccd1 _050_ a_4215_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X1976 a_7102_3087# _024_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X1977 a_2014_6711# a_1855_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1978 temp1.capload\[4\].cap.Y net23 a_8761_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1980 vssd1 a_3727_8181# a_3685_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1981 a_7201_10927# _078_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X1982 a_11684_11177# a_11435_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1983 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_10423_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X1984 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9955_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X1985 a_7663_6825# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1986 vccd1 _082_ a_7477_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1987 a_6647_6825# _046_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1988 a_4165_7913# _027_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1989 temp1.capload\[7\].cap.Y net26 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1990 vccd1 ctr\[5\] _088_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1991 a_7348_8725# _070_ a_7571_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1992 vssd1 ctr\[10\] _062_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1993 _038_ a_2845_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.172 ps=1.35 w=1 l=0.15
X1996 io_out[6] a_3215_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1997 a_1878_10499# _037_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1998 a_5946_8323# _028_ a_5864_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1999 a_2397_7663# a_1407_7663# a_2271_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2002 a_1941_4765# a_1407_4399# a_1846_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2003 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9411_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2004 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2007 a_4813_1385# _063_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2008 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11684_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X2009 vssd1 a_2531_5755# ctr\[6\] vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2010 vccd1 net5 a_11987_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2011 ctr\[1\] a_8327_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2012 vccd1 net3 a_10975_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2013 vccd1 _093_ a_8031_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X2016 a_7365_7497# a_6375_7125# a_7239_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2017 a_11703_4175# net8 temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2018 vccd1 a_4675_11690# in_measurement vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2019 a_10028_8207# a_9779_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2020 a_2014_9975# a_1855_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X2021 vssd1 a_2014_4511# a_1972_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2022 vssd1 _079_ a_8399_8215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2023 _025_ a_8859_2880# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2024 vccd1 a_2934_1653# a_2861_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2025 _063_ a_4392_1795# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2026 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2027 vssd1 a_2531_5755# a_2489_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2030 a_10415_10383# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X2031 ctr\[8\] a_2439_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2032 vssd1 net5 a_12079_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2033 a_11152_10927# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2034 a_4613_8207# _007_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2035 _043_ ctr\[2\] a_6461_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2036 a_3971_5487# ctr\[4\] _051_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2037 a_3024_6005# _027_ a_3247_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2038 _089_ a_8307_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2039 a_4443_4399# _022_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2040 a_7374_9839# _042_ a_7205_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X2041 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11960_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X2042 vssd1 temp1.dac_vout_notouch_ a_6559_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2044 a_7826_2767# a_7553_2773# a_7741_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2046 a_2934_1653# a_2766_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2048 a_8243_1679# a_7461_1685# a_8159_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2049 a_2861_1679# a_2327_1685# a_2766_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2050 vssd1 a_5324_7637# _070_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2051 a_2891_11849# a_2755_11689# a_2471_11703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2053 a_6629_8751# a_5639_8751# a_6503_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2054 a_12164_10703# net6 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2056 vssd1 net6 a_11527_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2057 a_2932_9269# _027_ a_3155_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2058 a_3191_1679# a_2493_1685# a_2934_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2059 a_4130_10357# a_3962_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2060 vccd1 a_10464_10615# a_10415_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X2061 a_4425_8213# a_4259_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2062 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9687_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2063 a_9013_3133# ctr\[13\] a_8941_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2064 vccd1 a_10096_7815# a_10047_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X2065 vccd1 _024_ a_8859_2880# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2066 a_6538_4765# a_6265_4399# a_6453_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2071 a_12256_5487# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2072 a_8377_3145# a_7387_2773# a_8251_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2073 vssd1 a_2271_6941# a_2442_6828# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2074 vccd1 io_out[5] a_4316_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2075 a_4471_10383# a_3689_10389# a_4387_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2076 a_1460_8725# net1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2077 a_2303_11703# a_2471_11703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2078 vssd1 net10 a_6817_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X2079 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11500_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X2080 _017_ a_4982_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X2081 a_5721_6397# ctr\[7\] a_5639_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X2083 a_1761_10927# _004_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X2084 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11612_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2085 vssd1 a_6423_10615# _073_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2086 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11251_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2087 vssd1 a_2439_7931# a_2397_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2088 vccd1 a_4319_11989# io_out[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2089 _067_ a_6395_1999# a_6633_1999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X2092 a_5365_5737# ctr\[8\] a_5283_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2093 a_3300_8751# io_out[2] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2095 vccd1 _080_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2096 _040_ a_3215_9813# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2097 a_2014_9975# a_1855_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2098 a_4698_8207# a_4259_8213# a_4613_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2099 _028_ a_5763_9867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2101 a_4319_11989# temp1.o_tempdelay vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2103 vssd1 a_2271_11293# a_2442_11180# vssd1 sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2104 a_11336_7663# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2105 net11 a_1460_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2107 a_10924_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2108 a_11500_9001# a_11251_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2109 a_8389_9001# _077_ a_8307_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2110 a_3983_3133# ctr\[9\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X2111 a_1855_6941# a_1407_6575# a_1761_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2112 a_11752_4087# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2113 vccd1 a_7994_2741# a_7921_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2115 a_5324_7637# ctr\[0\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2116 a_2355_4765# a_1573_4399# a_2271_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2117 a_7239_7119# a_6375_7125# a_6982_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2118 io_out[7] a_4319_11989# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2119 a_3153_4649# ctr\[6\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
R33 vssd1 net29 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2120 a_5813_11791# net22 temp1.capload\[3\].cap.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2121 a_7281_2528# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2122 vssd1 net3 a_9871_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2123 a_2007_5162# _053_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2124 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd a_10147_3863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2125 a_9034_7913# _095_ a_9034_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X2128 vssd1 net6 a_12079_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2129 vccd1 ctr\[3\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2130 a_2891_11849# a_2762_11593# a_2471_11703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2132 a_7473_5059# _076_ a_7377_5059# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2136 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref a_10423_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2137 vccd1 a_6706_4511# a_6633_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2138 a_4824_8585# a_4425_8213# a_4698_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2139 a_5077_7663# ctr\[2\] a_4971_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X2140 vssd1 a_2939_10615# _030_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2141 a_7072_10901# _070_ a_7295_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2142 vssd1 a_5283_5737# _076_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2143 a_6541_6031# _071_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X2144 a_2104_8527# a_1878_8323# a_1735_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2145 a_7921_2767# a_7387_2773# a_7826_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2146 a_7461_1685# a_7295_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2147 a_3981_4649# ctr\[8\] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2148 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref a_11435_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2149 a_10212_10089# a_9963_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2153 vssd1 net12 _075_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2154 a_2939_10615# _029_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X2157 a_5057_7439# ctr\[3\] a_5415_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2158 vssd1 a_8159_10383# a_8327_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2160 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_9233_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2161 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8951_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2162 a_9344_5487# _091_ a_9224_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X2163 a_5324_7637# ctr\[0\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2165 vssd1 a_6671_9019# a_6629_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2167 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd _080_ a_9773_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2168 a_1878_10499# _037_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X2169 a_3215_11989# in_measurement vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2170 a_3877_10383# _006_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2171 vssd1 a_3191_1679# a_3359_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2172 vssd1 a_10567_4917# net4 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2173 vccd1 a_2363_5853# a_2531_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2174 a_6633_4765# a_6099_4399# a_6538_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2175 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_10599_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X2177 vssd1 net4 a_10975_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2178 io_out[0] a_2442_6828# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X2179 a_3275_1679# a_2493_1685# a_3191_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2180 vccd1 _080_ a_8031_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X2181 vccd1 a_4404_9813# _006_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2182 a_1460_8725# net1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2183 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd a_10212_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X2185 _031_ a_2563_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2186 a_1460_1653# net1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2187 a_9588_4399# temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2188 _085_ a_7663_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2189 a_5123_8207# a_4425_8213# a_4866_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2191 temp1.dac_vout_notouch_ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd a_9496_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2192 vccd1 a_7407_7093# a_7323_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2193 a_7564_2473# _069_ _020_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X2194 a_4392_1795# _060_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2195 _047_ _096_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2196 vccd1 net12 a_3523_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2197 vccd1 ctr\[2\] _081_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2198 vssd1 a_3209_2197# _016_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2199 a_10599_6031# temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X2200 vccd1 a_4387_10383# a_4555_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2201 temp1.dac_vout_notouch_ net7 a_11152_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2202 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_12164_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2203 a_2471_11703# a_2762_11593# a_2713_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2204 a_1878_8323# _034_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X2205 vssd1 a_4330_1135# a_4436_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2206 a_3427_1385# _040_ a_3209_1109# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2207 vssd1 _052_ a_2313_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2208 a_5515_10357# temp1.o_tempdelay a_5996_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X2209 vssd1 ctr\[1\] a_5415_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2210 _068_ a_7060_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2211 _080_ a_8399_8215# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2212 temp1.capload\[2\].cap.Y net21 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2213 vssd1 net2 a_1959_1687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2214 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_8208_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2215 a_7829_10383# a_7295_10389# a_7734_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2216 vssd1 a_2363_5853# a_2531_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2218 a_4387_10383# a_3523_10389# a_4130_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2219 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd a_10139_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X2221 vccd1 a_2439_7931# a_2355_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2222 vccd1 a_2303_11703# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2223 _043_ _028_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2224 vssd1 _044_ a_5996_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2225 a_4057_10383# a_3523_10389# a_3962_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2226 a_9034_5487# ctr\[6\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X2227 a_9128_4399# temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2228 _060_ a_5363_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X2229 a_10600_7663# temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2230 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9963_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2231 vccd1 a_1731_2388# _015_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2232 a_11888_9839# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2233 vssd1 a_5843_1653# a_5801_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2234 ctr\[13\] a_8419_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2235 _081_ ctr\[2\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R34 net24 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2236 vccd1 net6 a_10975_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2238 vccd1 a_10188_6263# a_10139_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X2239 a_3425_5487# _050_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2240 a_4698_8207# a_4425_8213# a_4613_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2242 a_7295_5059# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2243 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11251_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2244 vssd1 a_7902_1653# a_7860_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2246 vssd1 net5 a_11527_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2247 vssd1 a_1735_9269# _003_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2248 vccd1 io_out[0] a_2200_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2249 _041_ a_4451_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X2250 a_1761_1135# _015_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2251 a_8951_7913# _083_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X2252 a_3074_8797# _035_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X2253 vccd1 _023_ a_4443_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2254 a_4977_1685# a_4811_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2255 vccd1 net3 a_11711_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2256 vssd1 ctr\[7\] a_3024_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X2257 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref a_11895_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2258 vccd1 a_2563_10357# _031_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2259 _074_ a_4255_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2260 a_1573_4399# a_1407_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2262 a_7288_9839# _082_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2263 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11796_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2264 a_4036_7093# _027_ a_4259_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2265 a_2493_1685# a_2327_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2266 a_12256_11791# net5 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2267 a_11152_4399# net4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2268 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2269 vssd1 a_2271_8029# a_2439_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2270 vssd1 net11 a_6099_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2271 a_4345_11837# a_4075_11471# a_4255_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X2272 vssd1 ctr\[9\] a_3852_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X2274 a_2755_11689# net12 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2275 a_3375_2767# a_2511_2773# a_3118_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2276 vssd1 _069_ a_7473_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2277 ctr\[5\] a_4831_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2278 a_7047_4765# a_6265_4399# a_6963_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2280 vssd1 a_3118_2741# a_3076_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2281 vccd1 io_out[2] a_3396_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2282 _075_ net12 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2283 a_2939_10615# _027_ a_3113_10721# vssd1 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2284 vccd1 net1 a_7387_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2285 a_9955_10703# temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2286 a_4613_1135# a_4436_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2287 _048_ _045_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2288 vssd1 _093_ a_9344_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X2289 a_5639_6397# _071_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2291 vccd1 ctr\[6\] _090_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2292 a_7649_10383# _008_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2294 a_2950_2767# a_2511_2773# a_2865_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2295 a_8115_4175# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2296 vccd1 a_4866_8181# a_4793_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2297 temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ a_11336_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X2298 a_6429_6549# _040_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
R35 net19 vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2299 vssd1 _031_ a_2104_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X2300 a_7205_10089# _070_ vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2301 a_11960_10089# a_11711_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X2302 vccd1 net5 a_11619_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2303 a_11428_8751# temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2304 a_10004_10615# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2305 a_7649_1679# _019_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2306 a_11059_6575# temp1.dac_vout_notouch_ temp1.dac_vout_notouch_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X2307 vccd1 a_2442_10092# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X2308 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref a_8114_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X2309 vssd1 ctr\[13\] _069_ vssd1 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2310 a_9034_7913# ctr\[2\] a_8951_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2311 a_5445_3561# _059_ a_5363_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2312 a_10140_9839# temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X2313 ctr\[5\] a_4831_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2314 a_4719_4399# _022_ a_4613_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2315 a_4663_6941# a_3965_6575# a_4406_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2316 a_4793_8207# a_4259_8213# a_4698_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2317 vssd1 a_6503_9117# a_6671_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2318 a_5904_4399# _047_ a_5601_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X2319 a_4153_3133# ctr\[8\] a_4065_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2320 a_4365_5737# _050_ _052_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X2321 a_6633_1999# ctr\[12\] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2322 vssd1 ctr\[10\] a_4259_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2323 net8 a_11527_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2324 vccd1 net3 a_11711_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X2325 a_9865_7439# _083_ vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2326 vccd1 a_3543_2741# a_3459_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2327 a_2271_1501# a_1573_1135# a_2014_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2328 vccd1 ctr\[2\] _045_ vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
C0 io_in[2] vssd1 0.228f
C1 io_in[3] vssd1 0.228f
C2 io_in[4] vssd1 0.228f
C3 io_in[5] vssd1 0.228f
C4 io_in[6] vssd1 0.228f
C5 io_in[7] vssd1 0.228f
C6 io_in[0] vssd1 2.51f
C7 io_in[1] vssd1 1.49f
C8 io_out[0] vssd1 2.56f
C9 io_out[1] vssd1 2.45f
C10 io_out[2] vssd1 2.83f
C11 io_out[3] vssd1 2.59f
C12 io_out[4] vssd1 2.62f
C13 io_out[5] vssd1 3.3f
C14 io_out[7] vssd1 2.75f
C15 io_out[6] vssd1 2.1f
C16 vccd1 vssd1 0.551p
C17 a_4813_1385# vssd1 0.253f  
C18 a_4613_1135# vssd1 0.227f  
C19 a_3427_1385# vssd1 0.253f  
C20 a_1761_1135# vssd1 0.23f  
C21 a_7060_1385# vssd1 0.502f  
C22 a_4982_1135# vssd1 0.55f  
C23 a_4436_1135# vssd1 0.498f  
C24 a_4330_1135# vssd1 0.578f  
C25 a_4153_1135# vssd1 0.5f  
C26 a_3834_1135# vssd1 0.535f  
C27 a_3209_1109# vssd1 0.55f  
C28 a_2271_1501# vssd1 0.609f  
C29 a_2439_1403# vssd1 0.817f  
C30 a_1846_1501# vssd1 0.626f  
C31 a_2014_1247# vssd1 0.581f  
C32 a_1573_1135# vssd1 1.43f  
C33 a_1407_1135# vssd1 1.81f  
C34 a_7649_1679# vssd1 0.23f  
C35 _067_ vssd1 0.967f  
C36 a_6633_1999# vssd1 0.211f  
C37 a_5165_1679# vssd1 0.23f  
C38 _063_ vssd1 1.02f  
C39 a_4069_1999# vssd1 0.21f  
C40 _066_ vssd1 1.04f  
C41 a_8159_1679# vssd1 0.609f  
C42 a_8327_1653# vssd1 0.817f  
C43 a_7734_1679# vssd1 0.626f  
C44 a_7902_1653# vssd1 0.581f  
C45 a_7461_1685# vssd1 1.43f  
C46 _019_ vssd1 0.87f  
C47 a_7295_1685# vssd1 1.81f  
C48 a_7019_1679# vssd1 0.524f  
C49 _068_ vssd1 1.06f  
C50 a_6395_1999# vssd1 0.706f  
C51 a_5675_1679# vssd1 0.609f  
C52 a_5843_1653# vssd1 0.817f  
C53 a_5250_1679# vssd1 0.626f  
C54 a_5418_1653# vssd1 0.581f  
C55 a_4977_1685# vssd1 1.43f  
C56 _017_ vssd1 1.28f  
C57 a_4811_1685# vssd1 1.81f  
C58 a_4392_1795# vssd1 0.502f  
C59 a_3877_1740# vssd1 0.446f  
C60 a_2681_1679# vssd1 0.23f  
C61 a_3191_1679# vssd1 0.609f  
C62 a_3359_1653# vssd1 0.817f  
C63 a_2766_1679# vssd1 0.626f  
C64 a_2934_1653# vssd1 0.581f  
C65 a_2493_1685# vssd1 1.43f  
C66 _018_ vssd1 1.2f  
C67 a_2327_1685# vssd1 1.81f  
C68 a_1959_1687# vssd1 0.648f  
C69 a_1460_1653# vssd1 0.648f  
C70 a_7473_2223# vssd1 0.21f  
C71 a_11844_2375# vssd1 0.525f  
C72 a_7281_2528# vssd1 0.446f  
C73 _064_ vssd1 1.1f  
C74 a_3427_2473# vssd1 0.253f  
C75 _015_ vssd1 1.19f  
C76 _062_ vssd1 1.66f  
C77 a_3209_2197# vssd1 0.55f  
C78 a_1731_2388# vssd1 0.524f  
C79 a_1407_2223# vssd1 0.524f  
C80 a_11711_2767# vssd1 0.525f  
C81 a_10975_2767# vssd1 0.525f  
C82 a_10423_2767# vssd1 0.525f  
C83 a_7019_2767# vssd1 0.238f  
C84 a_7741_2767# vssd1 0.23f  
C85 _069_ vssd1 0.895f  
C86 a_9319_2767# vssd1 0.698f  
C87 _025_ vssd1 0.688f  
C88 a_8859_2880# vssd1 0.619f  
C89 a_8251_2767# vssd1 0.609f  
C90 a_8419_2741# vssd1 0.817f  
C91 a_7826_2767# vssd1 0.626f  
C92 a_7994_2741# vssd1 0.581f  
C93 a_7553_2773# vssd1 1.43f  
C94 _020_ vssd1 1.06f  
C95 a_7387_2773# vssd1 1.81f  
C96 a_6375_2883# vssd1 0.858f  
C97 a_2865_2767# vssd1 0.23f  
C98 _058_ vssd1 1.15f  
C99 a_1665_3087# vssd1 0.211f  
C100 ctr\[13\] vssd1 2.85f  
C101 ctr\[12\] vssd1 4.61f  
C102 a_3983_3133# vssd1 0.729f  
C103 ctr\[10\] vssd1 3.83f  
C104 ctr\[11\] vssd1 3.66f  
C105 a_3375_2767# vssd1 0.609f  
C106 a_3543_2741# vssd1 0.817f  
C107 a_2950_2767# vssd1 0.626f  
C108 a_3118_2741# vssd1 0.581f  
C109 a_2677_2773# vssd1 1.43f  
C110 _016_ vssd1 1.12f  
C111 a_2511_2773# vssd1 1.81f  
C112 a_2092_2883# vssd1 0.502f  
C113 _057_ vssd1 0.704f  
C114 a_1427_3087# vssd1 0.706f  
C115 _060_ vssd1 3.51f  
C116 _059_ vssd1 1.01f  
C117 _065_ vssd1 3.55f  
C118 a_4709_3317# vssd1 0.432f  
C119 a_11711_3311# vssd1 0.525f  
C120 a_11251_3311# vssd1 0.525f  
C121 a_10791_3311# vssd1 0.525f  
C122 a_10331_3311# vssd1 0.525f  
C123 a_9871_3311# vssd1 0.525f  
C124 a_6009_3317# vssd1 0.665f  
C125 a_5363_3561# vssd1 0.858f  
C126 a_4815_3561# vssd1 0.697f  
C127 a_12212_4087# vssd1 0.525f  
C128 a_11752_4087# vssd1 0.525f  
C129 a_10515_3855# vssd1 0.525f  
C130 a_9319_3855# vssd1 0.525f  
C131 a_8164_4087# vssd1 0.525f  
C132 _054_ vssd1 2.44f  
C133 a_2507_3855# vssd1 0.253f  
C134 net3 vssd1 8.68f  
C135 net7 vssd1 5.95f  
C136 a_10975_3863# vssd1 0.648f  
C137 a_10147_3863# vssd1 0.648f  
C138 a_3739_4193# vssd1 0.56f  
C139 a_3307_4087# vssd1 0.56f  
C140 _055_ vssd1 4.38f  
C141 a_2289_3829# vssd1 0.55f  
C142 a_6453_4399# vssd1 0.23f  
C143 a_11803_4399# vssd1 0.525f  
C144 a_10975_4399# vssd1 0.525f  
C145 a_10515_4399# vssd1 0.525f  
C146 a_10004_4551# vssd1 0.525f  
C147 a_9411_4399# vssd1 0.525f  
C148 a_8951_4399# vssd1 0.525f  
C149 a_8031_4399# vssd1 0.525f  
C150 a_6963_4765# vssd1 0.609f  
C151 a_7131_4667# vssd1 0.97f  
C152 a_6538_4765# vssd1 0.626f  
C153 a_6706_4511# vssd1 0.581f  
C154 a_6265_4399# vssd1 1.43f  
C155 a_6099_4399# vssd1 1.81f  
C156 a_5819_4649# vssd1 0.253f  
C157 _011_ vssd1 1.03f  
C158 _024_ vssd1 3.59f  
C159 a_3981_4649# vssd1 0.203f  
C160 _061_ vssd1 1.52f  
C161 a_3153_4649# vssd1 0.203f  
C162 _056_ vssd1 0.896f  
C163 a_1761_4399# vssd1 0.23f  
C164 _047_ vssd1 0.822f  
C165 a_5601_4373# vssd1 0.55f  
C166 a_4443_4399# vssd1 0.729f  
C167 _023_ vssd1 1.86f  
C168 _022_ vssd1 1.87f  
C169 a_3852_4373# vssd1 0.655f  
C170 _021_ vssd1 2.01f  
C171 a_3024_4373# vssd1 0.655f  
C172 a_2271_4765# vssd1 0.609f  
C173 a_2439_4667# vssd1 0.817f  
C174 a_1846_4765# vssd1 0.626f  
C175 a_2014_4511# vssd1 0.581f  
C176 a_1573_4399# vssd1 1.43f  
C177 _014_ vssd1 1.14f  
C178 a_1407_4399# vssd1 1.81f  
C179 a_9319_4943# vssd1 0.525f  
C180 a_8031_4943# vssd1 0.525f  
C181 a_11527_4943# vssd1 0.698f  
C182 a_10567_4917# vssd1 0.698f  
C183 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vssd1 3.73f  
C184 a_7295_5059# vssd1 0.702f  
C185 _048_ vssd1 1.17f  
C186 _086_ vssd1 1.19f  
C187 a_6375_4943# vssd1 0.524f  
C188 _072_ vssd1 1.73f  
C189 _049_ vssd1 3.19f  
C190 a_2313_5175# vssd1 0.502f  
C191 _053_ vssd1 0.68f  
C192 a_2007_5162# vssd1 0.524f  
C193 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vssd1 1.92f  
C194 net8 vssd1 4.31f  
C195 a_12079_5487# vssd1 0.525f  
C196 net4 vssd1 5.48f  
C197 a_11619_5487# vssd1 0.525f  
C198 a_11159_5487# vssd1 0.525f  
C199 a_10239_5487# vssd1 0.648f  
C200 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd vssd1 2.34f  
C201 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd vssd1 2.92f  
C202 a_8951_5737# vssd1 0.333f  
C203 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref vssd1 4.32f  
C204 a_4257_5487# vssd1 0.211f  
C205 a_3425_5487# vssd1 0.21f  
C206 a_8031_5737# vssd1 0.333f  
C207 _052_ vssd1 1.6f  
C208 a_3885_5737# vssd1 0.238f  
C209 a_9034_5737# vssd1 0.723f  
C210 _091_ vssd1 2.6f  
C211 a_8114_5737# vssd1 0.723f  
C212 _087_ vssd1 2.18f  
C213 a_7203_5737# vssd1 0.702f  
C214 a_6191_5487# vssd1 0.524f  
C215 ctr\[8\] vssd1 6.7f  
C216 ctr\[9\] vssd1 4.32f  
C217 a_5283_5737# vssd1 0.642f  
C218 _090_ vssd1 2.34f  
C219 a_4215_5639# vssd1 0.706f  
C220 _050_ vssd1 2.9f  
C221 _051_ vssd1 0.768f  
C222 a_3233_5792# vssd1 0.446f  
C223 a_1853_5487# vssd1 0.23f  
C224 a_2363_5853# vssd1 0.609f  
C225 a_2531_5755# vssd1 0.97f  
C226 a_1938_5853# vssd1 0.626f  
C227 a_2106_5599# vssd1 0.581f  
C228 a_1665_5487# vssd1 1.43f  
C229 _013_ vssd1 0.994f  
C230 a_1499_5487# vssd1 1.81f  
C231 a_11987_6031# vssd1 0.525f  
C232 a_11527_6031# vssd1 0.525f  
C233 a_10648_6263# vssd1 0.525f  
C234 a_10188_6263# vssd1 0.525f  
C235 a_8569_6031# vssd1 0.227f  
C236 a_3153_6031# vssd1 0.203f  
C237 a_8392_6031# vssd1 0.498f  
C238 a_8286_6031# vssd1 0.578f  
C239 a_8109_6031# vssd1 0.5f  
C240 a_7790_6031# vssd1 0.535f  
C241 _094_ vssd1 1.04f  
C242 a_7111_6031# vssd1 0.698f  
C243 _092_ vssd1 1.01f  
C244 a_6541_6031# vssd1 0.673f  
C245 a_6375_6031# vssd1 0.641f  
C246 a_5639_6397# vssd1 0.729f  
C247 net10 vssd1 2.64f  
C248 ctr\[6\] vssd1 7.18f  
C249 a_3024_6005# vssd1 0.655f  
C250 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vssd1 1.98f  
C251 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd vssd1 1.47f  
C252 a_8951_6825# vssd1 0.333f  
C253 a_6647_6825# vssd1 0.253f  
C254 a_4153_6575# vssd1 0.23f  
C255 a_11987_6575# vssd1 0.525f  
C256 a_11435_6575# vssd1 0.525f  
C257 a_11108_6727# vssd1 0.525f  
C258 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref vssd1 2.39f  
C259 a_9034_6825# vssd1 0.723f  
C260 _085_ vssd1 1.58f  
C261 a_7663_6825# vssd1 0.702f  
C262 a_6429_6549# vssd1 0.55f  
C263 a_4663_6941# vssd1 0.609f  
C264 a_4831_6843# vssd1 0.97f  
C265 a_4238_6941# vssd1 0.626f  
C266 a_4406_6687# vssd1 0.581f  
C267 a_3965_6575# vssd1 1.43f  
C268 _012_ vssd1 1.41f  
C269 a_3799_6575# vssd1 1.81f  
C270 a_1761_6575# vssd1 0.216f  
C271 a_2271_6941# vssd1 0.599f  
C272 a_2442_6828# vssd1 1.41f  
C273 a_1855_6941# vssd1 0.627f  
C274 a_2014_6711# vssd1 0.587f  
C275 a_1573_6575# vssd1 1.39f  
C276 a_1407_6575# vssd1 1.77f  
C277 net11 vssd1 12.3f  
C278 a_12079_7119# vssd1 0.525f  
C279 net29 vssd1 1.08f  
C280 temp1.dac.vdac_single.einvp_batch\[0\].vref_29.HI vssd1 0.415f  
C281 a_8307_7235# vssd1 0.702f  
C282 _081_ vssd1 0.744f  
C283 a_4165_7119# vssd1 0.203f  
C284 a_2939_7119# vssd1 0.203f  
C285 a_6729_7119# vssd1 0.23f  
C286 a_5415_7439# vssd1 0.46f  
C287 a_5057_7439# vssd1 0.326f  
C288 _045_ vssd1 6.69f  
C289 a_4627_7439# vssd1 0.431f  
C290 a_2104_7439# vssd1 0.205f  
C291 _033_ vssd1 1.48f  
C292 _000_ vssd1 0.886f  
C293 a_7239_7119# vssd1 0.609f  
C294 a_7407_7093# vssd1 0.97f  
C295 a_6814_7119# vssd1 0.626f  
C296 a_6982_7093# vssd1 0.581f  
C297 a_6541_7125# vssd1 1.43f  
C298 _010_ vssd1 1.07f  
C299 a_6375_7125# vssd1 1.81f  
C300 a_4036_7093# vssd1 0.655f  
C301 a_2845_7119# vssd1 0.655f  
C302 ctr\[7\] vssd1 6.4f  
C303 net2 vssd1 4.7f  
C304 a_1878_7235# vssd1 0.443f  
C305 a_1735_7093# vssd1 0.65f  
C306 a_8951_7913# vssd1 0.333f  
C307 _046_ vssd1 1.23f  
C308 a_12079_7663# vssd1 0.525f  
C309 a_11619_7663# vssd1 0.525f  
C310 a_11159_7663# vssd1 0.525f  
C311 a_10423_7663# vssd1 0.525f  
C312 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vssd1 1.07f  
C313 a_10096_7815# vssd1 0.525f  
C314 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd vssd1 0.969f  
C315 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref vssd1 1.49f  
C316 a_9034_7913# vssd1 0.723f  
C317 _083_ vssd1 1.73f  
C318 _084_ vssd1 1.94f  
C319 _096_ vssd1 5.02f  
C320 a_4165_7913# vssd1 0.203f  
C321 a_3245_7913# vssd1 0.203f  
C322 a_1761_7663# vssd1 0.23f  
C323 a_5324_7637# vssd1 0.648f  
C324 a_4679_7637# vssd1 0.729f  
C325 ctr\[3\] vssd1 5.25f  
C326 a_4036_7637# vssd1 0.655f  
C327 ctr\[4\] vssd1 8.63f  
C328 a_3116_7637# vssd1 0.655f  
C329 a_2271_8029# vssd1 0.609f  
C330 a_2439_7931# vssd1 0.97f  
C331 a_1846_8029# vssd1 0.626f  
C332 a_2014_7775# vssd1 0.581f  
C333 a_1573_7663# vssd1 1.43f  
C334 a_1407_7663# vssd1 1.81f  
C335 a_11895_8207# vssd1 0.525f  
C336 a_10924_8439# vssd1 0.525f  
C337 a_9779_8207# vssd1 0.525f  
C338 a_8399_8215# vssd1 0.648f  
C339 _079_ vssd1 0.697f  
C340 a_7851_8323# vssd1 0.697f  
C341 a_7745_8323# vssd1 0.432f  
C342 ctr\[0\] vssd1 1.62f  
C343 a_4613_8207# vssd1 0.23f  
C344 a_3049_8207# vssd1 0.23f  
C345 a_2104_8527# vssd1 0.205f  
C346 _034_ vssd1 1.76f  
C347 _001_ vssd1 0.971f  
C348 a_5864_8323# vssd1 0.502f  
C349 a_5123_8207# vssd1 0.609f  
C350 a_5291_8181# vssd1 0.817f  
C351 a_4698_8207# vssd1 0.626f  
C352 a_4866_8181# vssd1 0.581f  
C353 a_4425_8213# vssd1 1.43f  
C354 a_4259_8213# vssd1 1.81f  
C355 a_3559_8207# vssd1 0.609f  
C356 a_3727_8181# vssd1 0.97f  
C357 a_3134_8207# vssd1 0.626f  
C358 a_3302_8181# vssd1 0.581f  
C359 a_2861_8213# vssd1 1.43f  
C360 a_2695_8213# vssd1 1.81f  
C361 a_1878_8323# vssd1 0.443f  
C362 a_1735_8181# vssd1 0.65f  
C363 a_9779_8751# vssd1 0.279f  
C364 a_10255_9001# vssd1 0.388f  
C365 a_9033_9001# vssd1 0.323f  
C366 _076_ vssd1 6.5f  
C367 _077_ vssd1 6.46f  
C368 a_7477_9001# vssd1 0.203f  
C369 ctr\[2\] vssd1 6.85f  
C370 a_5993_8751# vssd1 0.23f  
C371 a_11803_8751# vssd1 0.525f  
C372 a_11251_8751# vssd1 0.525f  
C373 a_10791_8751# vssd1 0.525f  
C374 _026_ vssd1 7.5f  
C375 a_9233_8751# vssd1 0.773f  
C376 _095_ vssd1 4.76f  
C377 _080_ vssd1 7.44f  
C378 _089_ vssd1 1.49f  
C379 a_8307_9001# vssd1 0.702f  
C380 _093_ vssd1 5.88f  
C381 a_7348_8725# vssd1 0.655f  
C382 a_6503_9117# vssd1 0.609f  
C383 a_6671_9019# vssd1 0.97f  
C384 a_6078_9117# vssd1 0.626f  
C385 a_6246_8863# vssd1 0.581f  
C386 a_5805_8751# vssd1 1.43f  
C387 a_5639_8751# vssd1 1.81f  
C388 a_3300_8751# vssd1 0.205f  
C389 _007_ vssd1 1.04f  
C390 a_4259_8757# vssd1 0.478f  
C391 _035_ vssd1 0.971f  
C392 _002_ vssd1 1.27f  
C393 _041_ vssd1 0.719f  
C394 a_4859_8916# vssd1 0.524f  
C395 a_4451_9001# vssd1 0.485f  
C396 a_3074_8797# vssd1 0.443f  
C397 a_2931_8903# vssd1 0.65f  
C398 net1 vssd1 10.9f  
C399 a_1460_8725# vssd1 0.648f  
C400 a_11803_9295# vssd1 0.525f  
C401 a_10699_9295# vssd1 0.525f  
C402 temp1.dac.vdac_single.einvp_batch\[0\].pupd_30.LO vssd1 0.479f  
C403 a_9687_9295# vssd1 0.525f  
C404 _088_ vssd1 0.872f  
C405 a_5911_9295# vssd1 0.253f  
C406 a_3061_9295# vssd1 0.203f  
C407 a_7571_9295# vssd1 0.525f  
C408 _009_ vssd1 1.07f  
C409 a_2104_9615# vssd1 0.205f  
C410 _036_ vssd1 0.985f  
C411 net30 vssd1 0.816f  
C412 temp1.dac.vdac_single.en_pupd vssd1 1.16f  
C413 _044_ vssd1 1.11f  
C414 _043_ vssd1 2.09f  
C415 a_5693_9269# vssd1 0.55f  
C416 ctr\[5\] vssd1 10f  
C417 a_2932_9269# vssd1 0.655f  
C418 a_1878_9411# vssd1 0.443f  
C419 a_1735_9269# vssd1 0.65f  
C420 a_6921_9839# vssd1 0.21f  
C421 a_7205_10089# vssd1 0.253f  
C422 a_11711_9839# vssd1 0.525f  
C423 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref vssd1 7.63f  
C424 a_11251_9839# vssd1 0.698f  
C425 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref vssd1 3.68f  
C426 a_10924_9991# vssd1 0.525f  
C427 a_9963_9839# vssd1 0.525f  
C428 a_9411_9839# vssd1 0.525f  
C429 a_7374_9839# vssd1 0.55f  
C430 _042_ vssd1 0.873f  
C431 _082_ vssd1 7.31f  
C432 a_6729_10144# vssd1 0.446f  
C433 a_4541_10089# vssd1 0.191f  
C434 a_1761_9839# vssd1 0.216f  
C435 a_5763_9867# vssd1 0.56f  
C436 _040_ vssd1 14.3f  
C437 a_4404_9813# vssd1 0.847f  
C438 _032_ vssd1 13f  
C439 a_3215_9813# vssd1 1.2f  
C440 a_2271_10205# vssd1 0.599f  
C441 a_2442_10092# vssd1 1.41f  
C442 a_1855_10205# vssd1 0.627f  
C443 a_2014_9975# vssd1 0.587f  
C444 a_1573_9839# vssd1 1.39f  
C445 _003_ vssd1 0.888f  
C446 a_1407_9839# vssd1 1.77f  
C447 a_11987_10383# vssd1 0.525f  
C448 a_11527_10383# vssd1 0.525f  
C449 a_10924_10615# vssd1 0.525f  
C450 a_10464_10615# vssd1 0.525f  
C451 a_10004_10615# vssd1 0.525f  
C452 a_9411_10383# vssd1 0.525f  
C453 a_7649_10383# vssd1 0.23f  
C454 a_3877_10383# vssd1 0.23f  
C455 _027_ vssd1 6.4f  
C456 _029_ vssd1 7.54f  
C457 a_2104_10703# vssd1 0.205f  
C458 _037_ vssd1 2.8f  
C459 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd vssd1 4.91f  
C460 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vssd1 7.27f  
C461 a_8159_10383# vssd1 0.609f  
C462 a_8327_10357# vssd1 0.97f  
C463 a_7734_10383# vssd1 0.626f  
C464 a_7902_10357# vssd1 0.581f  
C465 a_7461_10389# vssd1 1.43f  
C466 _008_ vssd1 0.999f  
C467 a_7295_10389# vssd1 1.81f  
C468 ctr\[1\] vssd1 10f  
C469 a_6423_10615# vssd1 0.619f  
C470 _071_ vssd1 4.61f  
C471 net9 vssd1 3.32f  
C472 _028_ vssd1 2.74f  
C473 a_5515_10357# vssd1 0.887f  
C474 temp_delay_last vssd1 1.49f  
C475 a_4387_10383# vssd1 0.609f  
C476 a_4555_10357# vssd1 0.817f  
C477 a_3962_10383# vssd1 0.626f  
C478 a_4130_10357# vssd1 0.581f  
C479 a_3689_10389# vssd1 1.43f  
C480 _006_ vssd1 1.21f  
C481 a_3523_10389# vssd1 1.81f  
C482 a_2939_10615# vssd1 0.56f  
C483 _030_ vssd1 0.7f  
C484 a_2563_10357# vssd1 0.698f  
C485 a_1878_10499# vssd1 0.443f  
C486 a_1735_10357# vssd1 0.65f  
C487 a_4220_10927# vssd1 0.205f  
C488 a_7201_11177# vssd1 0.203f  
C489 _039_ vssd1 1.06f  
C490 _038_ vssd1 2.43f  
C491 a_1761_10927# vssd1 0.216f  
C492 a_12079_10927# vssd1 0.525f  
C493 a_11435_10927# vssd1 0.525f  
C494 a_10975_10927# vssd1 0.525f  
C495 _075_ vssd1 0.745f  
C496 _078_ vssd1 2.11f  
C497 a_7072_10901# vssd1 0.655f  
C498 temp1.i_precharge_n vssd1 0.634f  
C499 a_6559_10927# vssd1 0.525f  
C500 _031_ vssd1 5.3f  
C501 a_3994_10973# vssd1 0.443f  
C502 a_3851_11079# vssd1 0.65f  
C503 a_2271_11293# vssd1 0.599f  
C504 a_2442_11180# vssd1 1.41f  
C505 a_1855_11293# vssd1 0.627f  
C506 a_2014_11063# vssd1 0.587f  
C507 a_1573_10927# vssd1 1.39f  
C508 _004_ vssd1 0.888f  
C509 a_1407_10927# vssd1 1.77f  
C510 a_12079_11471# vssd1 0.525f  
C511 a_11752_11703# vssd1 0.525f  
C512 temp1.capload\[15\].cap.Y vssd1 0.281f  
C513 temp1.capload\[14\].cap.Y vssd1 0.281f  
C514 temp1.capload\[0\].cap.Y vssd1 0.281f  
C515 temp1.capload\[5\].cap.Y vssd1 0.281f  
C516 temp1.capload\[2\].cap.Y vssd1 0.281f  
C517 net5 vssd1 9.17f  
C518 net6 vssd1 5.68f  
C519 temp1.dac_vout_notouch_ vssd1 55.2f  
C520 temp1.capload\[9\].cap_28.HI vssd1 0.415f  
C521 temp1.capload\[4\].cap_23.HI vssd1 0.415f  
C522 temp1.capload\[9\].cap.Y vssd1 0.281f  
C523 temp1.capload\[4\].cap.Y vssd1 0.281f  
C524 temp1.capload\[13\].cap.Y vssd1 0.281f  
C525 temp1.capload\[8\].cap.Y vssd1 0.281f  
C526 temp1.capload\[7\].cap.Y vssd1 0.281f  
C527 temp1.capload\[3\].cap.Y vssd1 0.281f  
C528 temp1.capload\[6\].cap.Y vssd1 0.281f  
C529 a_3309_11849# vssd1 0.23f  
C530 net28 vssd1 0.938f  
C531 net23 vssd1 1.13f  
C532 temp1.dcdel_out_n vssd1 0.613f  
C533 _074_ vssd1 0.725f  
C534 a_4675_11690# vssd1 0.524f  
C535 a_4255_11471# vssd1 0.508f  
C536 _073_ vssd1 3.47f  
C537 a_4075_11471# vssd1 0.604f  
C538 _070_ vssd1 9.95f  
C539 net12 vssd1 11.7f  
C540 _005_ vssd1 1.11f  
C541 a_2891_11849# vssd1 0.581f  
C542 a_2962_11748# vssd1 0.626f  
C543 a_2762_11593# vssd1 1.43f  
C544 a_2755_11689# vssd1 1.81f  
C545 a_2471_11703# vssd1 0.609f  
C546 a_2303_11703# vssd1 0.97f  
C547 temp1.capload\[15\].cap_19.HI vssd1 0.415f  
C548 net19 vssd1 1.09f  
C549 temp1.capload\[14\].cap_18.HI vssd1 0.415f  
C550 net18 vssd1 1.09f  
C551 temp1.capload\[0\].cap_13.HI vssd1 0.415f  
C552 net13 vssd1 1.09f  
C553 temp1.capload\[5\].cap_24.HI vssd1 0.415f  
C554 net24 vssd1 1.09f  
C555 net21 vssd1 1.37f  
C556 temp1.capload\[2\].cap_21.HI vssd1 0.415f  
C557 temp1.capload\[10\].cap_14.HI vssd1 0.415f  
C558 temp1.capload\[13\].cap_17.HI vssd1 0.415f  
C559 temp1.capload\[10\].cap.Y vssd1 0.281f  
C560 net14 vssd1 0.821f  
C561 temp1.capload\[12\].cap_16.HI vssd1 0.415f  
C562 net17 vssd1 1.09f  
C563 temp1.capload\[1\].cap.Y vssd1 0.281f  
C564 temp1.capload\[12\].cap.Y vssd1 0.281f  
C565 net16 vssd1 0.821f  
C566 net20 vssd1 1.09f  
C567 temp1.capload\[1\].cap_20.HI vssd1 0.415f  
C568 temp1.capload\[11\].cap_15.HI vssd1 0.415f  
C569 temp1.capload\[11\].cap.Y vssd1 0.281f  
C570 net15 vssd1 0.821f  
C571 temp1.dcdel_capnode_notouch_ vssd1 9.5f  
C572 net27 vssd1 1.16f  
C573 temp1.capload\[8\].cap_27.HI vssd1 0.415f  
C574 temp1.capload\[6\].cap_25.HI vssd1 0.415f  
C575 net25 vssd1 1.21f  
C576 net22 vssd1 1.12f  
C577 temp1.capload\[3\].cap_22.HI vssd1 0.415f  
C578 net26 vssd1 1.39f  
C579 temp1.capload\[7\].cap_26.HI vssd1 0.415f  
C580 temp1.o_tempdelay vssd1 2.92f  
C581 a_4319_11989# vssd1 1.2f  
C582 in_measurement vssd1 1.25f  
C583 a_3215_11989# vssd1 1.2f  
.ends

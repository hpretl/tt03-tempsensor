magic
tech sky130A
magscale 1 2
timestamp 1703959959
<< viali >>
rect 4353 12393 4387 12427
rect 5365 12257 5399 12291
rect 7389 12257 7423 12291
rect 5641 12189 5675 12223
rect 5733 12189 5767 12223
rect 6193 12189 6227 12223
rect 6475 12189 6509 12223
rect 6653 12189 6687 12223
rect 6745 12189 6779 12223
rect 7487 12189 7521 12223
rect 7665 12189 7699 12223
rect 7757 12189 7791 12223
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9689 12189 9723 12223
rect 10333 12189 10367 12223
rect 10609 12189 10643 12223
rect 10885 12189 10919 12223
rect 11161 12189 11195 12223
rect 3157 12121 3191 12155
rect 3525 12121 3559 12155
rect 4629 12121 4663 12155
rect 4629 11849 4663 11883
rect 3453 11713 3487 11747
rect 4813 11713 4847 11747
rect 5054 11713 5088 11747
rect 5227 11713 5261 11747
rect 5330 11713 5364 11747
rect 5457 11713 5491 11747
rect 5641 11713 5675 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 8217 11713 8251 11747
rect 8401 11713 8435 11747
rect 8677 11713 8711 11747
rect 8861 11711 8895 11745
rect 8976 11713 9010 11747
rect 9137 11713 9171 11747
rect 9505 11713 9539 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10149 11713 10183 11747
rect 10333 11713 10367 11747
rect 10425 11713 10459 11747
rect 10609 11713 10643 11747
rect 10701 11713 10735 11747
rect 10885 11713 10919 11747
rect 10977 11713 11011 11747
rect 11161 11713 11195 11747
rect 3709 11645 3743 11679
rect 4077 11645 4111 11679
rect 4537 11645 4571 11679
rect 11621 11645 11655 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 12449 11645 12483 11679
rect 4445 11577 4479 11611
rect 2329 11509 2363 11543
rect 4951 11509 4985 11543
rect 9229 11509 9263 11543
rect 11621 11509 11655 11543
rect 12449 11509 12483 11543
rect 3801 11305 3835 11339
rect 6929 11305 6963 11339
rect 6929 11169 6963 11203
rect 7021 11169 7055 11203
rect 7297 11169 7331 11203
rect 7757 11169 7791 11203
rect 10977 11169 11011 11203
rect 11437 11169 11471 11203
rect 12081 11169 12115 11203
rect 1409 11101 1443 11135
rect 1685 11101 1719 11135
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 6561 11101 6595 11135
rect 7205 11101 7239 11135
rect 7389 11101 7423 11135
rect 7481 11101 7515 11135
rect 7665 11101 7699 11135
rect 11345 11101 11379 11135
rect 11805 11101 11839 11135
rect 12449 11101 12483 11135
rect 2789 10965 2823 10999
rect 4537 10965 4571 10999
rect 11345 10965 11379 10999
rect 11805 10965 11839 10999
rect 12449 10965 12483 10999
rect 1685 10761 1719 10795
rect 2605 10761 2639 10795
rect 5825 10761 5859 10795
rect 6535 10761 6569 10795
rect 9781 10761 9815 10795
rect 11897 10761 11931 10795
rect 5089 10693 5123 10727
rect 6101 10693 6135 10727
rect 6745 10693 6779 10727
rect 1869 10625 1903 10659
rect 2145 10625 2179 10659
rect 2329 10625 2363 10659
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 3249 10625 3283 10659
rect 3792 10625 3826 10659
rect 4997 10625 5031 10659
rect 5733 10625 5767 10659
rect 5917 10625 5951 10659
rect 7564 10625 7598 10659
rect 9413 10625 9447 10659
rect 10333 10625 10367 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 11989 10625 12023 10659
rect 3525 10557 3559 10591
rect 7297 10557 7331 10591
rect 9873 10557 9907 10591
rect 10241 10557 10275 10591
rect 10701 10557 10735 10591
rect 11161 10557 11195 10591
rect 11897 10557 11931 10591
rect 12357 10557 12391 10591
rect 6377 10489 6411 10523
rect 9781 10489 9815 10523
rect 4905 10421 4939 10455
rect 5549 10421 5583 10455
rect 6561 10421 6595 10455
rect 8677 10421 8711 10455
rect 9873 10421 9907 10455
rect 10333 10421 10367 10455
rect 10793 10421 10827 10455
rect 12357 10421 12391 10455
rect 4353 10217 4387 10251
rect 6101 10217 6135 10251
rect 7665 10217 7699 10251
rect 11437 10217 11471 10251
rect 12081 10217 12115 10251
rect 6653 10149 6687 10183
rect 6929 10149 6963 10183
rect 9781 10081 9815 10115
rect 11161 10081 11195 10115
rect 12081 10081 12115 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 6929 10013 6963 10047
rect 7113 10013 7147 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 8493 10013 8527 10047
rect 9413 10013 9447 10047
rect 9965 10013 9999 10047
rect 10333 10013 10367 10047
rect 10793 10013 10827 10047
rect 11713 10013 11747 10047
rect 3525 9945 3559 9979
rect 11345 9945 11379 9979
rect 2789 9877 2823 9911
rect 3433 9877 3467 9911
rect 7297 9877 7331 9911
rect 8401 9877 8435 9911
rect 9781 9877 9815 9911
rect 10333 9877 10367 9911
rect 10793 9877 10827 9911
rect 1685 9673 1719 9707
rect 10057 9673 10091 9707
rect 11069 9673 11103 9707
rect 12173 9673 12207 9707
rect 1869 9537 1903 9571
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 3065 9537 3099 9571
rect 3249 9537 3283 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6101 9537 6135 9571
rect 8769 9537 8803 9571
rect 9689 9537 9723 9571
rect 10701 9537 10735 9571
rect 11805 9537 11839 9571
rect 2881 9469 2915 9503
rect 3157 9469 3191 9503
rect 3341 9469 3375 9503
rect 7573 9469 7607 9503
rect 7941 9469 7975 9503
rect 8033 9469 8067 9503
rect 10057 9401 10091 9435
rect 11069 9401 11103 9435
rect 12173 9401 12207 9435
rect 5641 9333 5675 9367
rect 7941 9333 7975 9367
rect 8677 9333 8711 9367
rect 4445 9129 4479 9163
rect 7297 9129 7331 9163
rect 8309 9129 8343 9163
rect 11161 9129 11195 9163
rect 8769 9061 8803 9095
rect 9689 9061 9723 9095
rect 10333 9061 10367 9095
rect 4721 8993 4755 9027
rect 5641 8993 5675 9027
rect 7481 8993 7515 9027
rect 7665 8993 7699 9027
rect 8401 8993 8435 9027
rect 8953 8993 8987 9027
rect 9045 8993 9079 9027
rect 10793 8993 10827 9027
rect 11253 8993 11287 9027
rect 11805 8993 11839 9027
rect 1685 8925 1719 8959
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3525 8925 3559 8959
rect 4261 8925 4295 8959
rect 4997 8925 5031 8959
rect 5897 8925 5931 8959
rect 7573 8925 7607 8959
rect 7757 8925 7791 8959
rect 8585 8925 8619 8959
rect 9249 8925 9283 8959
rect 9505 8925 9539 8959
rect 9781 8925 9815 8959
rect 9965 8925 9999 8959
rect 10333 8925 10367 8959
rect 10517 8925 10551 8959
rect 11161 8925 11195 8959
rect 11621 8925 11655 8959
rect 12173 8925 12207 8959
rect 8309 8857 8343 8891
rect 10149 8857 10183 8891
rect 1501 8789 1535 8823
rect 2881 8789 2915 8823
rect 4813 8789 4847 8823
rect 7021 8789 7055 8823
rect 9137 8789 9171 8823
rect 11621 8789 11655 8823
rect 12173 8789 12207 8823
rect 4077 8585 4111 8619
rect 6193 8585 6227 8619
rect 7205 8585 7239 8619
rect 8309 8585 8343 8619
rect 8585 8585 8619 8619
rect 10149 8585 10183 8619
rect 10793 8585 10827 8619
rect 12265 8585 12299 8619
rect 2964 8517 2998 8551
rect 4528 8517 4562 8551
rect 5825 8517 5859 8551
rect 6009 8517 6043 8551
rect 7665 8517 7699 8551
rect 1869 8449 1903 8483
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 2697 8449 2731 8483
rect 4261 8449 4295 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 8125 8449 8159 8483
rect 8401 8449 8435 8483
rect 9781 8449 9815 8483
rect 10149 8449 10183 8483
rect 10793 8449 10827 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 12265 8449 12299 8483
rect 7941 8381 7975 8415
rect 6469 8313 6503 8347
rect 1685 8245 1719 8279
rect 5641 8245 5675 8279
rect 7757 8245 7791 8279
rect 2789 8041 2823 8075
rect 3065 8041 3099 8075
rect 3985 8041 4019 8075
rect 5365 8041 5399 8075
rect 9965 8041 9999 8075
rect 10793 8041 10827 8075
rect 11529 7973 11563 8007
rect 11989 7973 12023 8007
rect 3433 7905 3467 7939
rect 4353 7905 4387 7939
rect 9781 7905 9815 7939
rect 10333 7905 10367 7939
rect 10793 7905 10827 7939
rect 11161 7905 11195 7939
rect 11621 7905 11655 7939
rect 12081 7905 12115 7939
rect 1409 7837 1443 7871
rect 1676 7837 1710 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3525 7837 3559 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 4445 7837 4479 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5549 7837 5583 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 8953 7837 8987 7871
rect 9111 7837 9145 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10425 7837 10459 7871
rect 12449 7837 12483 7871
rect 4905 7769 4939 7803
rect 9321 7769 9355 7803
rect 9597 7769 9631 7803
rect 4629 7701 4663 7735
rect 4813 7701 4847 7735
rect 6837 7701 6871 7735
rect 11529 7701 11563 7735
rect 11989 7701 12023 7735
rect 12449 7701 12483 7735
rect 3985 7497 4019 7531
rect 7757 7497 7791 7531
rect 8769 7497 8803 7531
rect 9965 7497 9999 7531
rect 12449 7497 12483 7531
rect 1869 7361 1903 7395
rect 2145 7361 2179 7395
rect 2329 7361 2363 7395
rect 2973 7361 3007 7395
rect 4169 7361 4203 7395
rect 4261 7361 4295 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5457 7361 5491 7395
rect 6101 7361 6135 7395
rect 6633 7361 6667 7395
rect 8309 7361 8343 7395
rect 8585 7361 8619 7395
rect 8861 7361 8895 7395
rect 9781 7361 9815 7395
rect 9965 7361 9999 7395
rect 12449 7361 12483 7395
rect 2881 7293 2915 7327
rect 3065 7293 3099 7327
rect 3157 7293 3191 7327
rect 4353 7293 4387 7327
rect 4445 7293 4479 7327
rect 6377 7293 6411 7327
rect 8401 7293 8435 7327
rect 8953 7293 8987 7327
rect 11989 7293 12023 7327
rect 12081 7293 12115 7327
rect 3341 7225 3375 7259
rect 1685 7157 1719 7191
rect 6009 7157 6043 7191
rect 8309 7157 8343 7191
rect 2789 6953 2823 6987
rect 6377 6953 6411 6987
rect 7665 6953 7699 6987
rect 10977 6953 11011 6987
rect 11805 6953 11839 6987
rect 12357 6953 12391 6987
rect 1685 6817 1719 6851
rect 7757 6817 7791 6851
rect 9597 6817 9631 6851
rect 11345 6817 11379 6851
rect 11437 6817 11471 6851
rect 11805 6817 11839 6851
rect 11989 6817 12023 6851
rect 12357 6817 12391 6851
rect 1409 6749 1443 6783
rect 3801 6749 3835 6783
rect 6561 6749 6595 6783
rect 6837 6749 6871 6783
rect 7941 6749 7975 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 8953 6749 8987 6783
rect 9111 6749 9145 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 9873 6749 9907 6783
rect 9965 6749 9999 6783
rect 10149 6749 10183 6783
rect 10977 6749 11011 6783
rect 4046 6681 4080 6715
rect 6745 6681 6779 6715
rect 7665 6681 7699 6715
rect 9321 6681 9355 6715
rect 5181 6613 5215 6647
rect 8125 6613 8159 6647
rect 9873 6613 9907 6647
rect 10057 6613 10091 6647
rect 2973 6409 3007 6443
rect 5917 6409 5951 6443
rect 6745 6409 6779 6443
rect 7297 6409 7331 6443
rect 10057 6409 10091 6443
rect 10517 6409 10551 6443
rect 11897 6409 11931 6443
rect 12357 6409 12391 6443
rect 5641 6341 5675 6375
rect 6862 6341 6896 6375
rect 3157 6273 3191 6307
rect 3341 6273 3375 6307
rect 5825 6273 5859 6307
rect 6009 6273 6043 6307
rect 6193 6273 6227 6307
rect 7205 6273 7239 6307
rect 10057 6273 10091 6307
rect 10517 6273 10551 6307
rect 11529 6273 11563 6307
rect 11989 6273 12023 6307
rect 12357 6273 12391 6307
rect 3249 6205 3283 6239
rect 3433 6205 3467 6239
rect 6377 6205 6411 6239
rect 6653 6205 6687 6239
rect 7757 6205 7791 6239
rect 8033 6205 8067 6239
rect 10425 6205 10459 6239
rect 10885 6205 10919 6239
rect 11897 6205 11931 6239
rect 7021 6137 7055 6171
rect 3433 5865 3467 5899
rect 5917 5865 5951 5899
rect 6377 5865 6411 5899
rect 7481 5865 7515 5899
rect 9597 5865 9631 5899
rect 11989 5865 12023 5899
rect 3801 5797 3835 5831
rect 5641 5797 5675 5831
rect 7665 5797 7699 5831
rect 4445 5729 4479 5763
rect 6561 5729 6595 5763
rect 7297 5729 7331 5763
rect 11621 5729 11655 5763
rect 11989 5729 12023 5763
rect 1501 5661 1535 5695
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 3617 5661 3651 5695
rect 4077 5661 4111 5695
rect 4537 5661 4571 5695
rect 5457 5661 5491 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6193 5661 6227 5695
rect 6653 5661 6687 5695
rect 7481 5661 7515 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9412 5661 9446 5695
rect 9689 5661 9723 5695
rect 9873 5661 9907 5695
rect 9965 5661 9999 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11161 5661 11195 5695
rect 11529 5661 11563 5695
rect 12081 5661 12115 5695
rect 12449 5661 12483 5695
rect 1768 5593 1802 5627
rect 3801 5593 3835 5627
rect 5273 5593 5307 5627
rect 7205 5593 7239 5627
rect 8191 5593 8225 5627
rect 8401 5593 8435 5627
rect 9091 5593 9125 5627
rect 9229 5593 9263 5627
rect 9321 5593 9355 5627
rect 2881 5525 2915 5559
rect 3985 5525 4019 5559
rect 4169 5525 4203 5559
rect 8677 5525 8711 5559
rect 9873 5525 9907 5559
rect 10149 5525 10183 5559
rect 10425 5525 10459 5559
rect 10701 5525 10735 5559
rect 11529 5525 11563 5559
rect 12449 5525 12483 5559
rect 1961 5321 1995 5355
rect 4997 5321 5031 5355
rect 6561 5321 6595 5355
rect 7757 5321 7791 5355
rect 8401 5321 8435 5355
rect 9689 5321 9723 5355
rect 11713 5321 11747 5355
rect 2605 5253 2639 5287
rect 7113 5253 7147 5287
rect 11621 5253 11655 5287
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 6377 5185 6411 5219
rect 6653 5175 6687 5209
rect 6837 5185 6871 5219
rect 7205 5185 7239 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 8033 5185 8067 5219
rect 9689 5185 9723 5219
rect 10701 5185 10735 5219
rect 8401 5117 8435 5151
rect 9321 5117 9355 5151
rect 6745 4981 6779 5015
rect 7481 4981 7515 5015
rect 10609 4981 10643 5015
rect 2789 4777 2823 4811
rect 7481 4777 7515 4811
rect 4445 4709 4479 4743
rect 8401 4709 8435 4743
rect 9873 4709 9907 4743
rect 10885 4709 10919 4743
rect 11345 4709 11379 4743
rect 12173 4709 12207 4743
rect 3157 4641 3191 4675
rect 3249 4641 3283 4675
rect 3341 4641 3375 4675
rect 3985 4641 4019 4675
rect 4997 4641 5031 4675
rect 8033 4641 8067 4675
rect 9321 4641 9355 4675
rect 9781 4641 9815 4675
rect 10517 4641 10551 4675
rect 10977 4641 11011 4675
rect 11805 4641 11839 4675
rect 1409 4573 1443 4607
rect 3433 4573 3467 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4261 4573 4295 4607
rect 4721 4573 4755 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 6101 4573 6135 4607
rect 8585 4573 8619 4607
rect 8769 4573 8803 4607
rect 8953 4573 8987 4607
rect 9413 4573 9447 4607
rect 10241 4573 10275 4607
rect 1676 4505 1710 4539
rect 5549 4505 5583 4539
rect 6346 4505 6380 4539
rect 8677 4505 8711 4539
rect 2973 4437 3007 4471
rect 3801 4437 3835 4471
rect 4629 4437 4663 4471
rect 4813 4437 4847 4471
rect 5181 4437 5215 4471
rect 5917 4437 5951 4471
rect 8401 4437 8435 4471
rect 9321 4437 9355 4471
rect 9735 4437 9769 4471
rect 9873 4437 9907 4471
rect 10885 4437 10919 4471
rect 11345 4437 11379 4471
rect 12173 4437 12207 4471
rect 2237 4233 2271 4267
rect 3249 4233 3283 4267
rect 4077 4233 4111 4267
rect 5917 4233 5951 4267
rect 9689 4233 9723 4267
rect 10885 4233 10919 4267
rect 11621 4233 11655 4267
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 2697 4097 2731 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 5089 4097 5123 4131
rect 5273 4097 5307 4131
rect 5825 4097 5859 4131
rect 6009 4097 6043 4131
rect 8033 4097 8067 4131
rect 8401 4097 8435 4131
rect 9321 4097 9355 4131
rect 9689 4097 9723 4131
rect 10149 4097 10183 4131
rect 10517 4097 10551 4131
rect 10885 4097 10919 4131
rect 10977 4097 11011 4131
rect 11989 4097 12023 4131
rect 3617 4029 3651 4063
rect 11621 4029 11655 4063
rect 12081 4029 12115 4063
rect 12449 4029 12483 4063
rect 11161 3961 11195 3995
rect 5181 3893 5215 3927
rect 8033 3893 8067 3927
rect 10333 3893 10367 3927
rect 12081 3893 12115 3927
rect 5089 3689 5123 3723
rect 5641 3689 5675 3723
rect 6009 3689 6043 3723
rect 10241 3621 10275 3655
rect 10701 3621 10735 3655
rect 11161 3621 11195 3655
rect 11621 3621 11655 3655
rect 12081 3621 12115 3655
rect 4997 3553 5031 3587
rect 5457 3553 5491 3587
rect 6101 3553 6135 3587
rect 9873 3553 9907 3587
rect 10333 3553 10367 3587
rect 10793 3553 10827 3587
rect 11253 3553 11287 3587
rect 11713 3553 11747 3587
rect 4629 3485 4663 3519
rect 5089 3485 5123 3519
rect 5641 3485 5675 3519
rect 6009 3485 6043 3519
rect 5365 3417 5399 3451
rect 5273 3349 5307 3383
rect 5825 3349 5859 3383
rect 6377 3349 6411 3383
rect 10241 3349 10275 3383
rect 10701 3349 10735 3383
rect 11161 3349 11195 3383
rect 11621 3349 11655 3383
rect 12081 3349 12115 3383
rect 1961 3145 1995 3179
rect 3893 3145 3927 3179
rect 4537 3145 4571 3179
rect 4997 3145 5031 3179
rect 6101 3145 6135 3179
rect 9061 3145 9095 3179
rect 9229 3145 9263 3179
rect 10793 3145 10827 3179
rect 11345 3145 11379 3179
rect 12081 3145 12115 3179
rect 2053 3077 2087 3111
rect 3985 3077 4019 3111
rect 4261 3077 4295 3111
rect 5825 3077 5859 3111
rect 7113 3077 7147 3111
rect 8861 3077 8895 3111
rect 9413 3077 9447 3111
rect 1593 3009 1627 3043
rect 2237 3009 2271 3043
rect 2780 3009 2814 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4813 3009 4847 3043
rect 4997 3009 5031 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 7645 3009 7679 3043
rect 10793 3009 10827 3043
rect 11345 3009 11379 3043
rect 12081 3009 12115 3043
rect 1685 2941 1719 2975
rect 2513 2941 2547 2975
rect 6009 2941 6043 2975
rect 6469 2941 6503 2975
rect 10425 2941 10459 2975
rect 10977 2941 11011 2975
rect 11713 2941 11747 2975
rect 5917 2873 5951 2907
rect 6837 2873 6871 2907
rect 2421 2805 2455 2839
rect 6377 2805 6411 2839
rect 7297 2805 7331 2839
rect 8769 2805 8803 2839
rect 9045 2805 9079 2839
rect 9505 2805 9539 2839
rect 1593 2601 1627 2635
rect 3157 2601 3191 2635
rect 7481 2601 7515 2635
rect 7205 2533 7239 2567
rect 11713 2533 11747 2567
rect 12081 2465 12115 2499
rect 1409 2397 1443 2431
rect 1869 2397 1903 2431
rect 3341 2397 3375 2431
rect 3617 2397 3651 2431
rect 4813 2397 4847 2431
rect 4905 2397 4939 2431
rect 5089 2397 5123 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 4721 2329 4755 2363
rect 1685 2261 1719 2295
rect 3525 2261 3559 2295
rect 4905 2261 4939 2295
rect 11713 2261 11747 2295
rect 3709 2057 3743 2091
rect 6193 2057 6227 2091
rect 7205 2057 7239 2091
rect 8677 2057 8711 2091
rect 4537 1989 4571 2023
rect 5080 1989 5114 2023
rect 7542 1989 7576 2023
rect 1685 1921 1719 1955
rect 1961 1921 1995 1955
rect 2329 1921 2363 1955
rect 2596 1921 2630 1955
rect 4077 1921 4111 1955
rect 4261 1921 4295 1955
rect 4353 1921 4387 1955
rect 4813 1921 4847 1955
rect 6561 1921 6595 1955
rect 7021 1921 7055 1955
rect 7297 1921 7331 1955
rect 3801 1853 3835 1887
rect 6469 1853 6503 1887
rect 1501 1785 1535 1819
rect 6929 1785 6963 1819
rect 2145 1717 2179 1751
rect 4077 1717 4111 1751
rect 4721 1717 4755 1751
rect 2789 1513 2823 1547
rect 3157 1513 3191 1547
rect 5273 1513 5307 1547
rect 7389 1513 7423 1547
rect 1409 1377 1443 1411
rect 1676 1309 1710 1343
rect 3341 1309 3375 1343
rect 3617 1309 3651 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4813 1309 4847 1343
rect 5089 1309 5123 1343
rect 7021 1309 7055 1343
rect 7205 1309 7239 1343
rect 4905 1241 4939 1275
rect 3525 1173 3559 1207
<< metal1 >>
rect 1104 12538 12788 12560
rect 1104 12486 2410 12538
rect 2462 12486 2474 12538
rect 2526 12486 2538 12538
rect 2590 12486 2602 12538
rect 2654 12486 2666 12538
rect 2718 12486 5331 12538
rect 5383 12486 5395 12538
rect 5447 12486 5459 12538
rect 5511 12486 5523 12538
rect 5575 12486 5587 12538
rect 5639 12486 8252 12538
rect 8304 12486 8316 12538
rect 8368 12486 8380 12538
rect 8432 12486 8444 12538
rect 8496 12486 8508 12538
rect 8560 12486 11173 12538
rect 11225 12486 11237 12538
rect 11289 12486 11301 12538
rect 11353 12486 11365 12538
rect 11417 12486 11429 12538
rect 11481 12486 12788 12538
rect 1104 12464 12788 12486
rect 4338 12384 4344 12436
rect 4396 12384 4402 12436
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12288 5411 12291
rect 5810 12288 5816 12300
rect 5399 12260 5816 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7423 12260 8064 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 5626 12180 5632 12232
rect 5684 12180 5690 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 1302 12112 1308 12164
rect 1360 12152 1366 12164
rect 3145 12155 3203 12161
rect 3145 12152 3157 12155
rect 1360 12124 3157 12152
rect 1360 12112 1366 12124
rect 3145 12121 3157 12124
rect 3191 12121 3203 12155
rect 3145 12115 3203 12121
rect 3510 12112 3516 12164
rect 3568 12112 3574 12164
rect 4617 12155 4675 12161
rect 4617 12121 4629 12155
rect 4663 12121 4675 12155
rect 4617 12115 4675 12121
rect 4632 12084 4660 12115
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 5736 12152 5764 12183
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 6454 12180 6460 12232
rect 6512 12229 6518 12232
rect 8036 12229 8064 12260
rect 6512 12220 6521 12229
rect 6641 12223 6699 12229
rect 6512 12192 6557 12220
rect 6512 12183 6521 12192
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6687 12192 6745 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7475 12223 7533 12229
rect 7475 12189 7487 12223
rect 7521 12220 7533 12223
rect 7653 12223 7711 12229
rect 7521 12192 7595 12220
rect 7521 12189 7533 12192
rect 7475 12183 7533 12189
rect 6512 12180 6518 12183
rect 5592 12124 5764 12152
rect 5592 12112 5598 12124
rect 6086 12112 6092 12164
rect 6144 12112 6150 12164
rect 7567 12152 7595 12192
rect 7653 12189 7665 12223
rect 7699 12220 7711 12223
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7699 12192 7757 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8220 12152 8248 12183
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 9171 12192 9229 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9217 12189 9229 12192
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 10042 12220 10048 12232
rect 9723 12192 10048 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 8956 12152 8984 12183
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10318 12180 10324 12232
rect 10376 12180 10382 12232
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 7567 12124 8984 12152
rect 6104 12084 6132 12112
rect 8956 12096 8984 12124
rect 4632 12056 6132 12084
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 1104 11994 12947 12016
rect 1104 11942 3870 11994
rect 3922 11942 3934 11994
rect 3986 11942 3998 11994
rect 4050 11942 4062 11994
rect 4114 11942 4126 11994
rect 4178 11942 6791 11994
rect 6843 11942 6855 11994
rect 6907 11942 6919 11994
rect 6971 11942 6983 11994
rect 7035 11942 7047 11994
rect 7099 11942 9712 11994
rect 9764 11942 9776 11994
rect 9828 11942 9840 11994
rect 9892 11942 9904 11994
rect 9956 11942 9968 11994
rect 10020 11942 12633 11994
rect 12685 11942 12697 11994
rect 12749 11942 12761 11994
rect 12813 11942 12825 11994
rect 12877 11942 12889 11994
rect 12941 11942 12947 11994
rect 1104 11920 12947 11942
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 3568 11852 4629 11880
rect 3568 11840 3574 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 5534 11840 5540 11892
rect 5592 11840 5598 11892
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 5810 11840 5816 11892
rect 5868 11840 5874 11892
rect 6178 11840 6184 11892
rect 6236 11840 6242 11892
rect 8386 11840 8392 11892
rect 8444 11840 8450 11892
rect 10042 11840 10048 11892
rect 10100 11840 10106 11892
rect 10318 11840 10324 11892
rect 10376 11840 10382 11892
rect 10594 11840 10600 11892
rect 10652 11840 10658 11892
rect 10870 11840 10876 11892
rect 10928 11840 10934 11892
rect 11146 11840 11152 11892
rect 11204 11840 11210 11892
rect 3441 11747 3499 11753
rect 3441 11713 3453 11747
rect 3487 11744 3499 11747
rect 3786 11744 3792 11756
rect 3487 11716 3792 11744
rect 3487 11713 3499 11716
rect 3441 11707 3499 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4540 11716 4813 11744
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4338 11676 4344 11688
rect 4111 11648 4344 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1360 11512 2329 11540
rect 1360 11500 1366 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2317 11503 2375 11509
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 3712 11540 3740 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4540 11685 4568 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 5042 11747 5100 11753
rect 5042 11713 5054 11747
rect 5088 11744 5100 11747
rect 5215 11747 5273 11753
rect 5215 11744 5227 11747
rect 5088 11716 5227 11744
rect 5088 11713 5100 11716
rect 5042 11707 5100 11713
rect 5215 11713 5227 11716
rect 5261 11713 5273 11747
rect 5215 11707 5273 11713
rect 5318 11747 5376 11753
rect 5318 11713 5330 11747
rect 5364 11744 5376 11747
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5364 11716 5457 11744
rect 5364 11713 5376 11716
rect 5318 11707 5376 11713
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5552 11744 5580 11840
rect 5644 11812 5672 11840
rect 5828 11812 5856 11840
rect 6196 11812 6224 11840
rect 5644 11784 5764 11812
rect 5828 11784 6040 11812
rect 6196 11784 6408 11812
rect 5736 11753 5764 11784
rect 6012 11753 6040 11784
rect 6380 11753 6408 11784
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5552 11716 5641 11744
rect 5445 11707 5503 11713
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11713 6239 11747
rect 6181 11707 6239 11713
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6730 11744 6736 11756
rect 6595 11716 6736 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11645 4583 11679
rect 5460 11676 5488 11707
rect 5920 11676 5948 11707
rect 6196 11676 6224 11707
rect 6454 11676 6460 11688
rect 5460 11648 6460 11676
rect 4525 11639 4583 11645
rect 6454 11636 6460 11648
rect 6512 11676 6518 11688
rect 6564 11676 6592 11707
rect 6730 11704 6736 11716
rect 6788 11744 6794 11756
rect 8404 11753 8432 11840
rect 10060 11812 10088 11840
rect 9784 11784 10088 11812
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 6788 11716 8217 11744
rect 6788 11704 6794 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 6512 11648 6592 11676
rect 8220 11676 8248 11707
rect 8680 11676 8708 11707
rect 8846 11704 8852 11756
rect 8904 11704 8910 11756
rect 8938 11704 8944 11756
rect 8996 11753 9002 11756
rect 9784 11753 9812 11784
rect 10336 11753 10364 11840
rect 10612 11753 10640 11840
rect 10888 11753 10916 11840
rect 11164 11753 11192 11840
rect 8996 11747 9022 11753
rect 9010 11713 9022 11747
rect 8996 11707 9022 11713
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9171 11716 9505 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 9999 11716 10149 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 8996 11704 9002 11707
rect 10152 11676 10180 11707
rect 10428 11676 10456 11707
rect 10704 11676 10732 11707
rect 10980 11676 11008 11707
rect 8220 11648 8708 11676
rect 6512 11636 6518 11648
rect 4430 11568 4436 11620
rect 4488 11568 4494 11620
rect 8680 11608 8708 11648
rect 9646 11648 11008 11676
rect 11609 11679 11667 11685
rect 8938 11608 8944 11620
rect 8680 11580 8944 11608
rect 8938 11568 8944 11580
rect 8996 11608 9002 11620
rect 9646 11608 9674 11648
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 8996 11580 9674 11608
rect 8996 11568 9002 11580
rect 3568 11512 3740 11540
rect 4939 11543 4997 11549
rect 3568 11500 3574 11512
rect 4939 11509 4951 11543
rect 4985 11540 4997 11543
rect 6086 11540 6092 11552
rect 4985 11512 6092 11540
rect 4985 11509 4997 11512
rect 4939 11503 4997 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 11624 11549 11652 11639
rect 11974 11636 11980 11688
rect 12032 11636 12038 11688
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8904 11512 9229 11540
rect 8904 11500 8910 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9217 11503 9275 11509
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 11882 11540 11888 11552
rect 11655 11512 11888 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 11882 11500 11888 11512
rect 11940 11540 11946 11552
rect 12452 11549 12480 11639
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 11940 11512 12449 11540
rect 11940 11500 11946 11512
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 1104 11450 12788 11472
rect 1104 11398 2410 11450
rect 2462 11398 2474 11450
rect 2526 11398 2538 11450
rect 2590 11398 2602 11450
rect 2654 11398 2666 11450
rect 2718 11398 5331 11450
rect 5383 11398 5395 11450
rect 5447 11398 5459 11450
rect 5511 11398 5523 11450
rect 5575 11398 5587 11450
rect 5639 11398 8252 11450
rect 8304 11398 8316 11450
rect 8368 11398 8380 11450
rect 8432 11398 8444 11450
rect 8496 11398 8508 11450
rect 8560 11398 11173 11450
rect 11225 11398 11237 11450
rect 11289 11398 11301 11450
rect 11353 11398 11365 11450
rect 11417 11398 11429 11450
rect 11481 11398 12788 11450
rect 1104 11376 12788 11398
rect 3786 11296 3792 11348
rect 3844 11296 3850 11348
rect 4430 11296 4436 11348
rect 4488 11296 4494 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6788 11308 6929 11336
rect 6788 11296 6794 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 4448 11268 4476 11296
rect 4448 11240 4752 11268
rect 1320 11172 4476 11200
rect 1320 11144 1348 11172
rect 1302 11092 1308 11144
rect 1360 11092 1366 11144
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1486 11132 1492 11144
rect 1443 11104 1492 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3844 11104 3985 11132
rect 3844 11092 3850 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 2590 11024 2596 11076
rect 2648 11064 2654 11076
rect 4264 11064 4292 11095
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4448 11141 4476 11172
rect 4724 11141 4752 11240
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 6963 11172 7021 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7009 11169 7021 11172
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7331 11172 7757 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11011 11172 11437 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11425 11169 11437 11172
rect 11471 11200 11483 11203
rect 11514 11200 11520 11212
rect 11471 11172 11520 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11514 11160 11520 11172
rect 11572 11200 11578 11212
rect 11974 11200 11980 11212
rect 11572 11172 11980 11200
rect 11572 11160 11578 11172
rect 11974 11160 11980 11172
rect 12032 11200 12038 11212
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 12032 11172 12081 11200
rect 12032 11160 12038 11172
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5810 11132 5816 11144
rect 4755 11104 5816 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 2648 11036 4292 11064
rect 4356 11064 4384 11092
rect 4540 11064 4568 11095
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 5166 11064 5172 11076
rect 4356 11036 5172 11064
rect 2648 11024 2654 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 5828 11064 5856 11092
rect 7484 11064 7512 11095
rect 5828 11036 7512 11064
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2777 10999 2835 11005
rect 2777 10996 2789 10999
rect 2372 10968 2789 10996
rect 2372 10956 2378 10968
rect 2777 10965 2789 10968
rect 2823 10965 2835 10999
rect 2777 10959 2835 10965
rect 4522 10956 4528 11008
rect 4580 10956 4586 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 7668 10996 7696 11095
rect 7340 10968 7696 10996
rect 7340 10956 7346 10968
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 11348 11005 11376 11095
rect 11808 11005 11836 11095
rect 11333 10999 11391 11005
rect 11333 10996 11345 10999
rect 10284 10968 11345 10996
rect 10284 10956 10290 10968
rect 11333 10965 11345 10968
rect 11379 10996 11391 10999
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11379 10968 11805 10996
rect 11379 10965 11391 10968
rect 11333 10959 11391 10965
rect 11793 10965 11805 10968
rect 11839 10996 11851 10999
rect 11882 10996 11888 11008
rect 11839 10968 11888 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 11882 10956 11888 10968
rect 11940 10996 11946 11008
rect 12452 11005 12480 11095
rect 12437 10999 12495 11005
rect 12437 10996 12449 10999
rect 11940 10968 12449 10996
rect 11940 10956 11946 10968
rect 12437 10965 12449 10968
rect 12483 10965 12495 10999
rect 12437 10959 12495 10965
rect 1104 10906 12947 10928
rect 1104 10854 3870 10906
rect 3922 10854 3934 10906
rect 3986 10854 3998 10906
rect 4050 10854 4062 10906
rect 4114 10854 4126 10906
rect 4178 10854 6791 10906
rect 6843 10854 6855 10906
rect 6907 10854 6919 10906
rect 6971 10854 6983 10906
rect 7035 10854 7047 10906
rect 7099 10854 9712 10906
rect 9764 10854 9776 10906
rect 9828 10854 9840 10906
rect 9892 10854 9904 10906
rect 9956 10854 9968 10906
rect 10020 10854 12633 10906
rect 12685 10854 12697 10906
rect 12749 10854 12761 10906
rect 12813 10854 12825 10906
rect 12877 10854 12889 10906
rect 12941 10854 12947 10906
rect 1104 10832 12947 10854
rect 1670 10752 1676 10804
rect 1728 10752 1734 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2590 10792 2596 10804
rect 2280 10764 2596 10792
rect 2280 10752 2286 10764
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6362 10792 6368 10804
rect 5859 10764 6368 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6362 10752 6368 10764
rect 6420 10792 6426 10804
rect 6523 10795 6581 10801
rect 6523 10792 6535 10795
rect 6420 10764 6535 10792
rect 6420 10752 6426 10764
rect 6523 10761 6535 10764
rect 6569 10761 6581 10795
rect 6523 10755 6581 10761
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 9815 10764 10272 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10244 10736 10272 10764
rect 11882 10752 11888 10804
rect 11940 10752 11946 10804
rect 2958 10724 2964 10736
rect 1872 10696 2964 10724
rect 1762 10616 1768 10668
rect 1820 10616 1826 10668
rect 1872 10665 1900 10696
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 3252 10696 5089 10724
rect 3252 10668 3280 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 6086 10684 6092 10736
rect 6144 10684 6150 10736
rect 6733 10727 6791 10733
rect 6733 10693 6745 10727
rect 6779 10724 6791 10727
rect 6914 10724 6920 10736
rect 6779 10696 6920 10724
rect 6779 10693 6791 10696
rect 6733 10687 6791 10693
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 10042 10724 10048 10736
rect 6972 10696 8708 10724
rect 6972 10684 6978 10696
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10656 2191 10659
rect 2222 10656 2228 10668
rect 2179 10628 2228 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2314 10616 2320 10668
rect 2372 10616 2378 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2731 10628 2881 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3142 10656 3148 10668
rect 3099 10628 3148 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3780 10659 3838 10665
rect 3780 10625 3792 10659
rect 3826 10656 3838 10659
rect 4338 10656 4344 10668
rect 3826 10628 4344 10656
rect 3826 10625 3838 10628
rect 3780 10619 3838 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4908 10628 4997 10656
rect 1780 10588 1808 10616
rect 2332 10588 2360 10616
rect 1780 10560 2360 10588
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10557 3571 10591
rect 3513 10551 3571 10557
rect 3528 10464 3556 10551
rect 3510 10412 3516 10464
rect 3568 10412 3574 10464
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 4908 10461 4936 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 7558 10665 7564 10668
rect 5960 10628 6592 10656
rect 5960 10616 5966 10628
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 5868 10560 6408 10588
rect 5868 10548 5874 10560
rect 6380 10529 6408 10560
rect 6365 10523 6423 10529
rect 6365 10489 6377 10523
rect 6411 10489 6423 10523
rect 6365 10483 6423 10489
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4672 10424 4905 10452
rect 4672 10412 4678 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 4893 10415 4951 10421
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 6564 10461 6592 10628
rect 7552 10619 7564 10665
rect 7558 10616 7564 10619
rect 7616 10616 7622 10668
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 8680 10464 8708 10696
rect 9416 10696 10048 10724
rect 9416 10665 9444 10696
rect 10042 10684 10048 10696
rect 10100 10684 10106 10736
rect 10226 10684 10232 10736
rect 10284 10684 10290 10736
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 9401 10619 9459 10625
rect 9876 10628 10333 10656
rect 9876 10597 9904 10628
rect 10321 10625 10333 10628
rect 10367 10656 10379 10659
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10367 10628 10793 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11572 10628 11989 10656
rect 11572 10616 11578 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9784 10560 9873 10588
rect 9784 10532 9812 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10100 10560 10241 10588
rect 10100 10548 10106 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 10275 10560 10701 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10689 10557 10701 10560
rect 10735 10588 10747 10591
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10735 10560 11161 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12345 10591 12403 10597
rect 12345 10588 12357 10591
rect 11940 10560 12357 10588
rect 11940 10548 11946 10560
rect 12345 10557 12357 10560
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 9766 10480 9772 10532
rect 9824 10480 9830 10532
rect 5537 10455 5595 10461
rect 5537 10452 5549 10455
rect 5040 10424 5549 10452
rect 5040 10412 5046 10424
rect 5537 10421 5549 10424
rect 5583 10421 5595 10455
rect 5537 10415 5595 10421
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 8662 10412 8668 10464
rect 8720 10412 8726 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 10226 10452 10232 10464
rect 9907 10424 10232 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10226 10412 10232 10424
rect 10284 10452 10290 10464
rect 12360 10461 12388 10551
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 10284 10424 10333 10452
rect 10284 10412 10290 10424
rect 10321 10421 10333 10424
rect 10367 10452 10379 10455
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10367 10424 10793 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 12345 10455 12403 10461
rect 12345 10421 12357 10455
rect 12391 10421 12403 10455
rect 12345 10415 12403 10421
rect 1104 10362 12788 10384
rect 1104 10310 2410 10362
rect 2462 10310 2474 10362
rect 2526 10310 2538 10362
rect 2590 10310 2602 10362
rect 2654 10310 2666 10362
rect 2718 10310 5331 10362
rect 5383 10310 5395 10362
rect 5447 10310 5459 10362
rect 5511 10310 5523 10362
rect 5575 10310 5587 10362
rect 5639 10310 8252 10362
rect 8304 10310 8316 10362
rect 8368 10310 8380 10362
rect 8432 10310 8444 10362
rect 8496 10310 8508 10362
rect 8560 10310 11173 10362
rect 11225 10310 11237 10362
rect 11289 10310 11301 10362
rect 11353 10310 11365 10362
rect 11417 10310 11429 10362
rect 11481 10310 12788 10362
rect 1104 10288 12788 10310
rect 4338 10208 4344 10260
rect 4396 10208 4402 10260
rect 4982 10208 4988 10260
rect 5040 10208 5046 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 5776 10220 6101 10248
rect 5776 10208 5782 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7616 10220 7665 10248
rect 7616 10208 7622 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 8662 10208 8668 10260
rect 8720 10208 8726 10260
rect 11425 10251 11483 10257
rect 11425 10217 11437 10251
rect 11471 10248 11483 10251
rect 11514 10248 11520 10260
rect 11471 10220 11520 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 5000 10112 5028 10208
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 3200 10084 5028 10112
rect 5092 10152 6653 10180
rect 3200 10072 3206 10084
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 1486 10044 1492 10056
rect 1443 10016 1492 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 4522 10004 4528 10056
rect 4580 10004 4586 10056
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4816 10053 4844 10084
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 3513 9979 3571 9985
rect 3513 9945 3525 9979
rect 3559 9976 3571 9979
rect 3602 9976 3608 9988
rect 3559 9948 3608 9976
rect 3559 9945 3571 9948
rect 3513 9939 3571 9945
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 2314 9908 2320 9920
rect 1820 9880 2320 9908
rect 1820 9868 1826 9880
rect 2314 9868 2320 9880
rect 2372 9908 2378 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2372 9880 2789 9908
rect 2372 9868 2378 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 4908 9908 4936 10007
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5092 10044 5120 10152
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 6917 10183 6975 10189
rect 6917 10149 6929 10183
rect 6963 10149 6975 10183
rect 6917 10143 6975 10149
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 6822 10112 6828 10124
rect 5224 10084 5764 10112
rect 5224 10072 5230 10084
rect 5736 10053 5764 10084
rect 5920 10084 6828 10112
rect 5920 10053 5948 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 6932 10112 6960 10143
rect 6932 10084 7512 10112
rect 5040 10016 5120 10044
rect 5721 10047 5779 10053
rect 5040 10004 5046 10016
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 5534 9908 5540 9920
rect 3467 9880 5540 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5736 9908 5764 10007
rect 6932 9976 6960 10007
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 7484 10053 7512 10084
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7208 9976 7236 10007
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 8168 10016 8493 10044
rect 8168 10004 8174 10016
rect 8481 10013 8493 10016
rect 8527 10044 8539 10047
rect 8680 10044 8708 10208
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 11149 10115 11207 10121
rect 9824 10084 10180 10112
rect 9824 10072 9830 10084
rect 10152 10056 10180 10084
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11440 10112 11468 10211
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11940 10220 12081 10248
rect 11940 10208 11946 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 12084 10121 12112 10211
rect 11195 10084 11468 10112
rect 12069 10115 12127 10121
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 12069 10081 12081 10115
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 8527 10016 8708 10044
rect 9401 10047 9459 10053
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9447 10016 9965 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9953 10013 9965 10016
rect 9999 10044 10011 10047
rect 10042 10044 10048 10056
rect 9999 10016 10048 10044
rect 9999 10013 10011 10016
rect 9953 10007 10011 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10134 10004 10140 10056
rect 10192 10044 10198 10056
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 10192 10016 10333 10044
rect 10192 10004 10198 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 6932 9948 8432 9976
rect 7098 9908 7104 9920
rect 5736 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9908 7162 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7156 9880 7297 9908
rect 7156 9868 7162 9880
rect 7285 9877 7297 9880
rect 7331 9908 7343 9911
rect 7374 9908 7380 9920
rect 7331 9880 7380 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7374 9868 7380 9880
rect 7432 9908 7438 9920
rect 7650 9908 7656 9920
rect 7432 9880 7656 9908
rect 7432 9868 7438 9880
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 8404 9917 8432 9948
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8570 9908 8576 9920
rect 8435 9880 8576 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 10226 9908 10232 9920
rect 9815 9880 10232 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 10226 9868 10232 9880
rect 10284 9908 10290 9920
rect 10796 9917 10824 10007
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11333 9979 11391 9985
rect 11333 9945 11345 9979
rect 11379 9976 11391 9979
rect 11514 9976 11520 9988
rect 11379 9948 11520 9976
rect 11379 9945 11391 9948
rect 11333 9939 11391 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10284 9880 10333 9908
rect 10284 9868 10290 9880
rect 10321 9877 10333 9880
rect 10367 9908 10379 9911
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10367 9880 10793 9908
rect 10367 9877 10379 9880
rect 10321 9871 10379 9877
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 10781 9871 10839 9877
rect 1104 9818 12947 9840
rect 1104 9766 3870 9818
rect 3922 9766 3934 9818
rect 3986 9766 3998 9818
rect 4050 9766 4062 9818
rect 4114 9766 4126 9818
rect 4178 9766 6791 9818
rect 6843 9766 6855 9818
rect 6907 9766 6919 9818
rect 6971 9766 6983 9818
rect 7035 9766 7047 9818
rect 7099 9766 9712 9818
rect 9764 9766 9776 9818
rect 9828 9766 9840 9818
rect 9892 9766 9904 9818
rect 9956 9766 9968 9818
rect 10020 9766 12633 9818
rect 12685 9766 12697 9818
rect 12749 9766 12761 9818
rect 12813 9766 12825 9818
rect 12877 9766 12889 9818
rect 12941 9766 12947 9818
rect 1104 9744 12947 9766
rect 1670 9664 1676 9716
rect 1728 9664 1734 9716
rect 10045 9707 10103 9713
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10226 9704 10232 9716
rect 10091 9676 10232 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 3142 9636 3148 9648
rect 3068 9608 3148 9636
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2222 9568 2228 9580
rect 2179 9540 2228 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 1872 9500 1900 9531
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 3068 9577 3096 9608
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 10060 9636 10088 9667
rect 10226 9664 10232 9676
rect 10284 9704 10290 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 10284 9676 11069 9704
rect 10284 9664 10290 9676
rect 5592 9608 6224 9636
rect 5592 9596 5598 9608
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 5828 9577 5856 9608
rect 6196 9580 6224 9608
rect 9600 9608 10088 9636
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6086 9528 6092 9580
rect 6144 9528 6150 9580
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 6288 9540 8769 9568
rect 2869 9503 2927 9509
rect 2869 9500 2881 9503
rect 1872 9472 2881 9500
rect 2869 9469 2881 9472
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3602 9500 3608 9512
rect 3375 9472 3608 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 3160 9432 3188 9463
rect 3602 9460 3608 9472
rect 3660 9500 3666 9512
rect 4430 9500 4436 9512
rect 3660 9472 4436 9500
rect 3660 9460 3666 9472
rect 4430 9460 4436 9472
rect 4488 9500 4494 9512
rect 4982 9500 4988 9512
rect 4488 9472 4988 9500
rect 4488 9460 4494 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 6288 9500 6316 9540
rect 8757 9537 8769 9540
rect 8803 9568 8815 9571
rect 9490 9568 9496 9580
rect 8803 9540 9496 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 5224 9472 6316 9500
rect 5224 9460 5230 9472
rect 6546 9460 6552 9512
rect 6604 9460 6610 9512
rect 7558 9460 7564 9512
rect 7616 9460 7622 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7975 9472 8033 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 9600 9500 9628 9608
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 10042 9568 10048 9580
rect 9723 9540 10048 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 8021 9463 8079 9469
rect 9416 9472 9628 9500
rect 5184 9432 5212 9460
rect 3160 9404 5212 9432
rect 5629 9367 5687 9373
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 5718 9364 5724 9376
rect 5675 9336 5724 9364
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6564 9364 6592 9460
rect 9416 9432 9444 9472
rect 7944 9404 9444 9432
rect 10045 9435 10103 9441
rect 7944 9373 7972 9404
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 10134 9432 10140 9444
rect 10091 9404 10140 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 10612 9432 10640 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 12161 9707 12219 9713
rect 12161 9673 12173 9707
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 11054 9568 11060 9580
rect 10735 9540 11060 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11054 9528 11060 9540
rect 11112 9568 11118 9580
rect 11698 9568 11704 9580
rect 11112 9540 11704 9568
rect 11112 9528 11118 9540
rect 11698 9528 11704 9540
rect 11756 9568 11762 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11756 9540 11805 9568
rect 11756 9528 11762 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 10962 9432 10968 9444
rect 10612 9404 10968 9432
rect 10962 9392 10968 9404
rect 11020 9432 11026 9444
rect 12176 9441 12204 9667
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 11020 9404 11069 9432
rect 11020 9392 11026 9404
rect 11057 9401 11069 9404
rect 11103 9432 11115 9435
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 11103 9404 12173 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 12161 9401 12173 9404
rect 12207 9401 12219 9435
rect 12161 9395 12219 9401
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 6564 9336 7941 9364
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 7929 9327 7987 9333
rect 8662 9324 8668 9376
rect 8720 9324 8726 9376
rect 1104 9274 12788 9296
rect 1104 9222 2410 9274
rect 2462 9222 2474 9274
rect 2526 9222 2538 9274
rect 2590 9222 2602 9274
rect 2654 9222 2666 9274
rect 2718 9222 5331 9274
rect 5383 9222 5395 9274
rect 5447 9222 5459 9274
rect 5511 9222 5523 9274
rect 5575 9222 5587 9274
rect 5639 9222 8252 9274
rect 8304 9222 8316 9274
rect 8368 9222 8380 9274
rect 8432 9222 8444 9274
rect 8496 9222 8508 9274
rect 8560 9222 11173 9274
rect 11225 9222 11237 9274
rect 11289 9222 11301 9274
rect 11353 9222 11365 9274
rect 11417 9222 11429 9274
rect 11481 9222 12788 9274
rect 1104 9200 12788 9222
rect 4430 9120 4436 9172
rect 4488 9120 4494 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7558 9160 7564 9172
rect 7331 9132 7564 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8570 9160 8576 9172
rect 8343 9132 8576 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8312 9092 8340 9123
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 8662 9120 8668 9172
rect 8720 9120 8726 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11020 9132 11161 9160
rect 11020 9120 11026 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 7576 9064 8340 9092
rect 4709 9027 4767 9033
rect 1320 8996 3556 9024
rect 1320 8968 1348 8996
rect 1302 8916 1308 8968
rect 1360 8916 1366 8968
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2038 8956 2044 8968
rect 1719 8928 2044 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 3528 8965 3556 8996
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 4755 8996 5028 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 3559 8928 3648 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 2240 8888 2268 8916
rect 3344 8888 3372 8919
rect 2240 8860 3372 8888
rect 3620 8832 3648 8928
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 5000 8965 5028 8996
rect 5552 8996 5641 9024
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5552 8900 5580 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7248 8996 7481 9024
rect 7248 8984 7254 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 5885 8959 5943 8965
rect 5885 8956 5897 8959
rect 5776 8928 5897 8956
rect 5776 8916 5782 8928
rect 5885 8925 5897 8928
rect 5931 8925 5943 8959
rect 5885 8919 5943 8925
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 7576 8965 7604 9064
rect 7650 8984 7656 9036
rect 7708 8984 7714 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 7892 8996 8401 9024
rect 7892 8984 7898 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7484 8928 7573 8956
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 7300 8888 7328 8916
rect 7484 8900 7512 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 8573 8959 8631 8965
rect 7791 8928 8524 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 5592 8860 7328 8888
rect 5592 8848 5598 8860
rect 7466 8848 7472 8900
rect 7524 8848 7530 8900
rect 8294 8848 8300 8900
rect 8352 8848 8358 8900
rect 8496 8888 8524 8928
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8680 8956 8708 9120
rect 8757 9095 8815 9101
rect 8757 9061 8769 9095
rect 8803 9092 8815 9095
rect 9677 9095 9735 9101
rect 8803 9064 9076 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 8938 9024 8944 9036
rect 8619 8928 8708 8956
rect 8772 8996 8944 9024
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8772 8888 8800 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9048 9033 9076 9064
rect 9677 9061 9689 9095
rect 9723 9092 9735 9095
rect 9723 9064 9996 9092
rect 9723 9061 9735 9064
rect 9677 9055 9735 9061
rect 9033 9027 9091 9033
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9968 9024 9996 9064
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 10100 9064 10333 9092
rect 10100 9052 10106 9064
rect 10321 9061 10333 9064
rect 10367 9061 10379 9095
rect 10321 9055 10379 9061
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 9079 8996 9812 9024
rect 9968 8996 10793 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9237 8959 9295 8965
rect 9237 8956 9249 8959
rect 9180 8928 9249 8956
rect 9180 8916 9186 8928
rect 9237 8925 9249 8928
rect 9283 8925 9295 8959
rect 9237 8919 9295 8925
rect 9490 8916 9496 8968
rect 9548 8916 9554 8968
rect 9784 8965 9812 8996
rect 10336 8965 10364 8996
rect 10781 8993 10793 8996
rect 10827 9024 10839 9027
rect 11054 9024 11060 9036
rect 10827 8996 11060 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 11112 8996 11253 9024
rect 11112 8984 11118 8996
rect 11241 8993 11253 8996
rect 11287 9024 11299 9027
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11287 8996 11805 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 8496 8860 8800 8888
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 2682 8820 2688 8832
rect 1544 8792 2688 8820
rect 1544 8780 1550 8792
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 3326 8820 3332 8832
rect 2915 8792 3332 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3602 8780 3608 8832
rect 3660 8780 3666 8832
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6696 8792 7021 8820
rect 6696 8780 6702 8792
rect 7009 8789 7021 8792
rect 7055 8820 7067 8823
rect 8846 8820 8852 8832
rect 7055 8792 8852 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 9088 8792 9137 8820
rect 9088 8780 9094 8792
rect 9125 8789 9137 8792
rect 9171 8820 9183 8823
rect 9968 8820 9996 8919
rect 10134 8848 10140 8900
rect 10192 8848 10198 8900
rect 10520 8888 10548 8919
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 11020 8928 11161 8956
rect 11020 8916 11026 8928
rect 11149 8925 11161 8928
rect 11195 8956 11207 8959
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11195 8928 11621 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 10244 8860 10548 8888
rect 10244 8832 10272 8860
rect 9171 8792 9996 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 11624 8829 11652 8919
rect 12176 8829 12204 8919
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 12161 8823 12219 8829
rect 12161 8820 12173 8823
rect 11655 8792 12173 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 12161 8789 12173 8792
rect 12207 8789 12219 8823
rect 12161 8783 12219 8789
rect 1104 8730 12947 8752
rect 1104 8678 3870 8730
rect 3922 8678 3934 8730
rect 3986 8678 3998 8730
rect 4050 8678 4062 8730
rect 4114 8678 4126 8730
rect 4178 8678 6791 8730
rect 6843 8678 6855 8730
rect 6907 8678 6919 8730
rect 6971 8678 6983 8730
rect 7035 8678 7047 8730
rect 7099 8678 9712 8730
rect 9764 8678 9776 8730
rect 9828 8678 9840 8730
rect 9892 8678 9904 8730
rect 9956 8678 9968 8730
rect 10020 8678 12633 8730
rect 12685 8678 12697 8730
rect 12749 8678 12761 8730
rect 12813 8678 12825 8730
rect 12877 8678 12889 8730
rect 12941 8678 12947 8730
rect 1104 8656 12947 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 2740 8588 3556 8616
rect 2740 8576 2746 8588
rect 1872 8520 2636 8548
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 1872 8489 1900 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2222 8480 2228 8492
rect 2179 8452 2228 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 1780 8412 1808 8440
rect 2332 8412 2360 8443
rect 1780 8384 2360 8412
rect 2608 8344 2636 8520
rect 2700 8489 2728 8576
rect 2952 8551 3010 8557
rect 2952 8517 2964 8551
rect 2998 8548 3010 8551
rect 3326 8548 3332 8560
rect 2998 8520 3332 8548
rect 2998 8517 3010 8520
rect 2952 8511 3010 8517
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 3528 8492 3556 8588
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3660 8588 4077 8616
rect 3660 8576 3666 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4798 8576 4804 8628
rect 4856 8576 4862 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5132 8588 6040 8616
rect 5132 8576 5138 8588
rect 4516 8551 4574 8557
rect 4516 8517 4528 8551
rect 4562 8548 4574 8551
rect 4816 8548 4844 8576
rect 4562 8520 4844 8548
rect 4562 8517 4574 8520
rect 4516 8511 4574 8517
rect 5810 8508 5816 8560
rect 5868 8508 5874 8560
rect 6012 8557 6040 8588
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6144 8588 6193 8616
rect 6144 8576 6150 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6181 8579 6239 8585
rect 7190 8576 7196 8628
rect 7248 8576 7254 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 9030 8616 9036 8628
rect 8619 8588 9036 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 5997 8551 6055 8557
rect 5997 8517 6009 8551
rect 6043 8548 6055 8551
rect 6638 8548 6644 8560
rect 6043 8520 6644 8548
rect 6043 8517 6055 8520
rect 5997 8511 6055 8517
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 7650 8508 7656 8560
rect 7708 8508 7714 8560
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3568 8452 4261 8480
rect 3568 8440 3574 8452
rect 4249 8449 4261 8452
rect 4295 8480 4307 8483
rect 5534 8480 5540 8492
rect 4295 8452 5540 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5828 8480 5856 8508
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5828 8478 6040 8480
rect 6196 8478 6377 8480
rect 5828 8452 6377 8478
rect 6012 8450 6224 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6656 8480 6684 8508
rect 6595 8452 6684 8480
rect 7101 8483 7159 8489
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 2608 8316 2728 8344
rect 1670 8236 1676 8288
rect 1728 8236 1734 8288
rect 2700 8276 2728 8316
rect 5994 8304 6000 8356
rect 6052 8344 6058 8356
rect 6454 8344 6460 8356
rect 6052 8316 6460 8344
rect 6052 8304 6058 8316
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 7116 8344 7144 8443
rect 7300 8412 7328 8443
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8312 8480 8340 8579
rect 9030 8576 9036 8588
rect 9088 8616 9094 8628
rect 9214 8616 9220 8628
rect 9088 8588 9220 8616
rect 9088 8576 9094 8588
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10137 8619 10195 8625
rect 10137 8616 10149 8619
rect 10008 8588 10149 8616
rect 10008 8576 10014 8588
rect 10137 8585 10149 8588
rect 10183 8616 10195 8619
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10183 8588 10793 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10781 8585 10793 8588
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 8312 8452 8401 8480
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 10042 8480 10048 8492
rect 9815 8452 10048 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10796 8489 10824 8579
rect 10962 8576 10968 8588
rect 11020 8616 11026 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 11020 8588 12265 8616
rect 11020 8576 11026 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 12268 8489 12296 8579
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 11112 8452 11161 8480
rect 11112 8440 11118 8452
rect 11149 8449 11161 8452
rect 11195 8480 11207 8483
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11195 8452 11897 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7300 8384 7941 8412
rect 7929 8381 7941 8384
rect 7975 8412 7987 8415
rect 8294 8412 8300 8424
rect 7975 8384 8300 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 8036 8356 8064 8384
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 7116 8316 7788 8344
rect 7760 8288 7788 8316
rect 8018 8304 8024 8356
rect 8076 8304 8082 8356
rect 3970 8276 3976 8288
rect 2700 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 5718 8276 5724 8288
rect 5675 8248 5724 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 1104 8186 12788 8208
rect 1104 8134 2410 8186
rect 2462 8134 2474 8186
rect 2526 8134 2538 8186
rect 2590 8134 2602 8186
rect 2654 8134 2666 8186
rect 2718 8134 5331 8186
rect 5383 8134 5395 8186
rect 5447 8134 5459 8186
rect 5511 8134 5523 8186
rect 5575 8134 5587 8186
rect 5639 8134 8252 8186
rect 8304 8134 8316 8186
rect 8368 8134 8380 8186
rect 8432 8134 8444 8186
rect 8496 8134 8508 8186
rect 8560 8134 11173 8186
rect 11225 8134 11237 8186
rect 11289 8134 11301 8186
rect 11353 8134 11365 8186
rect 11417 8134 11429 8186
rect 11481 8134 12788 8186
rect 1104 8112 12788 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 1820 8044 2789 8072
rect 1820 8032 1826 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 3970 8032 3976 8084
rect 4028 8032 4034 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4798 8072 4804 8084
rect 4304 8044 4804 8072
rect 4304 8032 4310 8044
rect 4798 8032 4804 8044
rect 4856 8072 4862 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 4856 8044 5365 8072
rect 4856 8032 4862 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10008 8044 10793 8072
rect 10008 8032 10014 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3252 7936 3280 8032
rect 8938 7964 8944 8016
rect 8996 7964 9002 8016
rect 10796 8004 10824 8035
rect 11517 8007 11575 8013
rect 11517 8004 11529 8007
rect 10796 7976 11529 8004
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 3252 7908 3433 7936
rect 3421 7905 3433 7908
rect 3467 7936 3479 7939
rect 3694 7936 3700 7948
rect 3467 7908 3700 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 3694 7896 3700 7908
rect 3752 7936 3758 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3752 7908 4353 7936
rect 3752 7896 3758 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 8956 7936 8984 7964
rect 10796 7945 10824 7976
rect 9769 7939 9827 7945
rect 8956 7908 9444 7936
rect 4341 7899 4399 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 1486 7868 1492 7880
rect 1443 7840 1492 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 1670 7877 1676 7880
rect 1664 7868 1676 7877
rect 1631 7840 1676 7868
rect 1664 7831 1676 7840
rect 1670 7828 1676 7831
rect 1728 7828 1734 7880
rect 3160 7868 3188 7896
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3160 7840 3249 7868
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3252 7800 3280 7831
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 3510 7828 3516 7880
rect 3568 7828 3574 7880
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4172 7800 4200 7831
rect 3252 7772 4200 7800
rect 4264 7800 4292 7831
rect 4430 7828 4436 7880
rect 4488 7828 4494 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5074 7868 5080 7880
rect 5031 7840 5080 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5215 7840 5549 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5537 7837 5549 7840
rect 5583 7868 5595 7871
rect 5718 7868 5724 7880
rect 5583 7840 5724 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6512 7840 6745 7868
rect 6512 7828 6518 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7834 7868 7840 7880
rect 6963 7840 7840 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 9122 7877 9128 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9099 7871 9128 7877
rect 9099 7837 9111 7871
rect 9099 7831 9128 7837
rect 9122 7828 9128 7831
rect 9180 7828 9186 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9416 7877 9444 7908
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 9815 7908 10333 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 10321 7905 10333 7908
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 4893 7803 4951 7809
rect 4893 7800 4905 7803
rect 4264 7772 4905 7800
rect 4893 7769 4905 7772
rect 4939 7800 4951 7803
rect 5442 7800 5448 7812
rect 4939 7772 5448 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 9309 7803 9367 7809
rect 9309 7769 9321 7803
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 9585 7803 9643 7809
rect 9585 7769 9597 7803
rect 9631 7800 9643 7803
rect 9692 7800 9720 7831
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10042 7868 10048 7880
rect 9999 7840 10048 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10428 7800 10456 7831
rect 9631 7772 10456 7800
rect 9631 7769 9643 7772
rect 9585 7763 9643 7769
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 3660 7704 4629 7732
rect 3660 7692 3666 7704
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 4617 7695 4675 7701
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 6270 7732 6276 7744
rect 4847 7704 6276 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 6696 7704 6837 7732
rect 6696 7692 6702 7704
rect 6825 7701 6837 7704
rect 6871 7701 6883 7735
rect 6825 7695 6883 7701
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9324 7732 9352 7763
rect 11072 7744 11100 7976
rect 11517 7973 11529 7976
rect 11563 8004 11575 8007
rect 11977 8007 12035 8013
rect 11977 8004 11989 8007
rect 11563 7976 11989 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 11977 7973 11989 7976
rect 12023 7973 12035 8007
rect 11977 7967 12035 7973
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11195 7908 11621 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11609 7905 11621 7908
rect 11655 7936 11667 7939
rect 12066 7936 12072 7948
rect 11655 7908 12072 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 12452 7744 12480 7831
rect 8812 7704 9352 7732
rect 8812 7692 8818 7704
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 11112 7704 11529 7732
rect 11112 7692 11118 7704
rect 11517 7701 11529 7704
rect 11563 7732 11575 7735
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 11563 7704 11989 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 11977 7701 11989 7704
rect 12023 7732 12035 7735
rect 12434 7732 12440 7744
rect 12023 7704 12440 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 1104 7642 12947 7664
rect 1104 7590 3870 7642
rect 3922 7590 3934 7642
rect 3986 7590 3998 7642
rect 4050 7590 4062 7642
rect 4114 7590 4126 7642
rect 4178 7590 6791 7642
rect 6843 7590 6855 7642
rect 6907 7590 6919 7642
rect 6971 7590 6983 7642
rect 7035 7590 7047 7642
rect 7099 7590 9712 7642
rect 9764 7590 9776 7642
rect 9828 7590 9840 7642
rect 9892 7590 9904 7642
rect 9956 7590 9968 7642
rect 10020 7590 12633 7642
rect 12685 7590 12697 7642
rect 12749 7590 12761 7642
rect 12813 7590 12825 7642
rect 12877 7590 12889 7642
rect 12941 7590 12947 7642
rect 1104 7568 12947 7590
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 2746 7500 3985 7528
rect 2746 7460 2774 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 5500 7500 7757 7528
rect 5500 7488 5506 7500
rect 7745 7497 7757 7500
rect 7791 7528 7803 7531
rect 8570 7528 8576 7540
rect 7791 7500 8576 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8754 7488 8760 7540
rect 8812 7488 8818 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10042 7528 10048 7540
rect 9999 7500 10048 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 12434 7488 12440 7540
rect 12492 7488 12498 7540
rect 1872 7432 2774 7460
rect 1872 7401 1900 7432
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3142 7460 3148 7472
rect 2924 7432 3148 7460
rect 2924 7420 2930 7432
rect 3142 7420 3148 7432
rect 3200 7460 3206 7472
rect 3200 7432 4200 7460
rect 3200 7420 3206 7432
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2222 7392 2228 7404
rect 2179 7364 2228 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2314 7352 2320 7404
rect 2372 7352 2378 7404
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3694 7392 3700 7404
rect 3007 7364 3700 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3694 7352 3700 7364
rect 3752 7392 3758 7404
rect 4172 7401 4200 7432
rect 4264 7432 5120 7460
rect 4264 7401 4292 7432
rect 5092 7404 5120 7432
rect 4157 7395 4215 7401
rect 3752 7364 3924 7392
rect 3752 7352 3758 7364
rect 2866 7284 2872 7336
rect 2924 7284 2930 7336
rect 3050 7284 3056 7336
rect 3108 7284 3114 7336
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 3786 7284 3792 7336
rect 3844 7284 3850 7336
rect 3329 7259 3387 7265
rect 3329 7225 3341 7259
rect 3375 7256 3387 7259
rect 3804 7256 3832 7284
rect 3375 7228 3832 7256
rect 3896 7256 3924 7364
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5460 7401 5488 7488
rect 6270 7460 6276 7472
rect 6104 7432 6276 7460
rect 6104 7401 6132 7432
rect 6270 7420 6276 7432
rect 6328 7460 6334 7472
rect 8110 7460 8116 7472
rect 6328 7432 8116 7460
rect 6328 7420 6334 7432
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8772 7460 8800 7488
rect 8772 7432 9812 7460
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 6512 7364 6633 7392
rect 6512 7352 6518 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 6621 7355 6679 7361
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8297 7395 8355 7401
rect 8297 7392 8309 7395
rect 8076 7364 8309 7392
rect 8076 7352 8082 7364
rect 8297 7361 8309 7364
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 4356 7256 4384 7287
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 3896 7228 4384 7256
rect 3375 7225 3387 7228
rect 3329 7219 3387 7225
rect 1670 7148 1676 7200
rect 1728 7148 1734 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4448 7188 4476 7284
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 6380 7256 6408 7287
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 7800 7296 8401 7324
rect 7800 7284 7806 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8588 7324 8616 7355
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 9784 7401 9812 7432
rect 12452 7401 12480 7488
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8588 7296 8953 7324
rect 8389 7287 8447 7293
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9858 7324 9864 7336
rect 9272 7296 9864 7324
rect 9272 7284 9278 7296
rect 9858 7284 9864 7296
rect 9916 7324 9922 7336
rect 9968 7324 9996 7355
rect 9916 7296 9996 7324
rect 11977 7327 12035 7333
rect 9916 7284 9922 7296
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 12023 7296 12081 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 5592 7228 6408 7256
rect 5592 7216 5598 7228
rect 3568 7160 4476 7188
rect 3568 7148 3574 7160
rect 5994 7148 6000 7200
rect 6052 7148 6058 7200
rect 6380 7188 6408 7228
rect 6546 7188 6552 7200
rect 6380 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7524 7160 8309 7188
rect 7524 7148 7530 7160
rect 8297 7157 8309 7160
rect 8343 7157 8355 7191
rect 8297 7151 8355 7157
rect 1104 7098 12788 7120
rect 1104 7046 2410 7098
rect 2462 7046 2474 7098
rect 2526 7046 2538 7098
rect 2590 7046 2602 7098
rect 2654 7046 2666 7098
rect 2718 7046 5331 7098
rect 5383 7046 5395 7098
rect 5447 7046 5459 7098
rect 5511 7046 5523 7098
rect 5575 7046 5587 7098
rect 5639 7046 8252 7098
rect 8304 7046 8316 7098
rect 8368 7046 8380 7098
rect 8432 7046 8444 7098
rect 8496 7046 8508 7098
rect 8560 7046 11173 7098
rect 11225 7046 11237 7098
rect 11289 7046 11301 7098
rect 11353 7046 11365 7098
rect 11417 7046 11429 7098
rect 11481 7046 12788 7098
rect 1104 7024 12788 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2314 6984 2320 6996
rect 1820 6956 2320 6984
rect 1820 6944 1826 6956
rect 2314 6944 2320 6956
rect 2372 6984 2378 6996
rect 2777 6987 2835 6993
rect 2777 6984 2789 6987
rect 2372 6956 2789 6984
rect 2372 6944 2378 6956
rect 2777 6953 2789 6956
rect 2823 6953 2835 6987
rect 2777 6947 2835 6953
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 6454 6984 6460 6996
rect 6411 6956 6460 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7524 6956 7665 6984
rect 7524 6944 7530 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 10965 6987 11023 6993
rect 10965 6953 10977 6987
rect 11011 6984 11023 6987
rect 11054 6984 11060 6996
rect 11011 6956 11060 6984
rect 11011 6953 11023 6956
rect 10965 6947 11023 6953
rect 11054 6944 11060 6956
rect 11112 6984 11118 6996
rect 11793 6987 11851 6993
rect 11793 6984 11805 6987
rect 11112 6956 11805 6984
rect 11112 6944 11118 6956
rect 11793 6953 11805 6956
rect 11839 6984 11851 6987
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 11839 6956 12357 6984
rect 11839 6953 11851 6956
rect 11793 6947 11851 6953
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 3142 6916 3148 6928
rect 2740 6888 3148 6916
rect 2740 6876 2746 6888
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 8938 6876 8944 6928
rect 8996 6876 9002 6928
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 6178 6848 6184 6860
rect 5736 6820 6184 6848
rect 5736 6792 5764 6820
rect 6178 6808 6184 6820
rect 6236 6848 6242 6860
rect 7742 6848 7748 6860
rect 6236 6820 6592 6848
rect 6236 6808 6242 6820
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 1452 6752 3801 6780
rect 1452 6740 1458 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6564 6789 6592 6820
rect 7392 6820 7748 6848
rect 7392 6792 7420 6820
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8956 6848 8984 6876
rect 11808 6857 11836 6947
rect 9585 6851 9643 6857
rect 8956 6820 9444 6848
rect 9416 6792 9444 6820
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 9631 6820 11345 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6696 6752 6837 6780
rect 6696 6740 6702 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7892 6752 7941 6780
rect 7892 6740 7898 6752
rect 7929 6749 7941 6752
rect 7975 6780 7987 6783
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7975 6752 8309 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8570 6780 8576 6792
rect 8435 6752 8576 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 9122 6789 9128 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8628 6752 8953 6780
rect 8628 6740 8634 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9099 6783 9128 6789
rect 9099 6749 9111 6783
rect 9099 6743 9128 6749
rect 9122 6740 9128 6743
rect 9180 6740 9186 6792
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 4034 6715 4092 6721
rect 4034 6712 4046 6715
rect 3476 6684 4046 6712
rect 3476 6672 3482 6684
rect 4034 6681 4046 6684
rect 4080 6681 4092 6715
rect 6012 6712 6040 6740
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 6012 6684 6745 6712
rect 4034 6675 4092 6681
rect 6656 6656 6684 6684
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7653 6715 7711 6721
rect 7653 6712 7665 6715
rect 7248 6684 7665 6712
rect 7248 6672 7254 6684
rect 7653 6681 7665 6684
rect 7699 6712 7711 6715
rect 8018 6712 8024 6724
rect 7699 6684 8024 6712
rect 7699 6681 7711 6684
rect 7653 6675 7711 6681
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 9309 6715 9367 6721
rect 8128 6684 8984 6712
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4890 6644 4896 6656
rect 3844 6616 4896 6644
rect 3844 6604 3850 6616
rect 4890 6604 4896 6616
rect 4948 6644 4954 6656
rect 5166 6644 5172 6656
rect 4948 6616 5172 6644
rect 4948 6604 4954 6616
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 6638 6604 6644 6656
rect 6696 6604 6702 6656
rect 8128 6653 8156 6684
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6613 8171 6647
rect 8956 6644 8984 6684
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 9692 6712 9720 6743
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 10152 6789 10180 6820
rect 11333 6817 11345 6820
rect 11379 6848 11391 6851
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 11379 6820 11437 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11425 6817 11437 6820
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 11793 6851 11851 6857
rect 11793 6817 11805 6851
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12066 6848 12072 6860
rect 12023 6820 12072 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12360 6857 12388 6947
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 9355 6684 9720 6712
rect 9968 6712 9996 6743
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11054 6780 11060 6792
rect 11011 6752 11060 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 10244 6712 10272 6740
rect 9968 6684 10272 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 9324 6644 9352 6675
rect 8956 6616 9352 6644
rect 9861 6647 9919 6653
rect 8113 6607 8171 6613
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 9950 6644 9956 6656
rect 9907 6616 9956 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10318 6644 10324 6656
rect 10091 6616 10324 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 1104 6554 12947 6576
rect 1104 6502 3870 6554
rect 3922 6502 3934 6554
rect 3986 6502 3998 6554
rect 4050 6502 4062 6554
rect 4114 6502 4126 6554
rect 4178 6502 6791 6554
rect 6843 6502 6855 6554
rect 6907 6502 6919 6554
rect 6971 6502 6983 6554
rect 7035 6502 7047 6554
rect 7099 6502 9712 6554
rect 9764 6502 9776 6554
rect 9828 6502 9840 6554
rect 9892 6502 9904 6554
rect 9956 6502 9968 6554
rect 10020 6502 12633 6554
rect 12685 6502 12697 6554
rect 12749 6502 12761 6554
rect 12813 6502 12825 6554
rect 12877 6502 12889 6554
rect 12941 6502 12947 6554
rect 1104 6480 12947 6502
rect 2958 6400 2964 6452
rect 3016 6400 3022 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 5960 6412 6745 6440
rect 5960 6400 5966 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6440 7343 6443
rect 8662 6440 8668 6452
rect 7331 6412 8668 6440
rect 7331 6409 7343 6412
rect 7285 6403 7343 6409
rect 8662 6400 8668 6412
rect 8720 6440 8726 6452
rect 8938 6440 8944 6452
rect 8720 6412 8944 6440
rect 8720 6400 8726 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 10045 6443 10103 6449
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10091 6412 10517 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10505 6409 10517 6412
rect 10551 6440 10563 6443
rect 11054 6440 11060 6452
rect 10551 6412 11060 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 11054 6400 11060 6412
rect 11112 6440 11118 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11112 6412 11897 6440
rect 11112 6400 11118 6412
rect 11885 6409 11897 6412
rect 11931 6440 11943 6443
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 11931 6412 12357 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 5629 6375 5687 6381
rect 5629 6372 5641 6375
rect 3108 6344 5641 6372
rect 3108 6332 3114 6344
rect 5629 6341 5641 6344
rect 5675 6341 5687 6375
rect 6850 6375 6908 6381
rect 6850 6372 6862 6375
rect 5629 6335 5687 6341
rect 6012 6344 6862 6372
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 3694 6304 3700 6316
rect 3375 6276 3700 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 3234 6196 3240 6248
rect 3292 6196 3298 6248
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6205 3479 6239
rect 5644 6236 5672 6335
rect 6012 6316 6040 6344
rect 6850 6341 6862 6344
rect 6896 6341 6908 6375
rect 6850 6335 6908 6341
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6227 6276 7205 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10100 6276 10517 6304
rect 10100 6264 10106 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11606 6304 11612 6316
rect 11563 6276 11612 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 11606 6264 11612 6276
rect 11664 6304 11670 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11664 6276 11989 6304
rect 11664 6264 11670 6276
rect 11977 6273 11989 6276
rect 12023 6304 12035 6307
rect 12066 6304 12072 6316
rect 12023 6276 12072 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12360 6313 12388 6403
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5644 6208 6377 6236
rect 3421 6199 3479 6205
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 6641 6199 6699 6205
rect 7024 6208 7757 6236
rect 2884 6168 2912 6196
rect 3436 6168 3464 6199
rect 2884 6140 3464 6168
rect 5810 6128 5816 6180
rect 5868 6168 5874 6180
rect 6270 6168 6276 6180
rect 5868 6140 6276 6168
rect 5868 6128 5874 6140
rect 6270 6128 6276 6140
rect 6328 6168 6334 6180
rect 6656 6168 6684 6199
rect 7024 6177 7052 6208
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8570 6236 8576 6248
rect 8067 6208 8576 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 8570 6196 8576 6208
rect 8628 6236 8634 6248
rect 9122 6236 9128 6248
rect 8628 6208 9128 6236
rect 8628 6196 8634 6208
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 10376 6208 10425 6236
rect 10376 6196 10382 6208
rect 10413 6205 10425 6208
rect 10459 6236 10471 6239
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10459 6208 10885 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12360 6236 12388 6267
rect 11940 6208 12388 6236
rect 11940 6196 11946 6208
rect 6328 6140 6684 6168
rect 7009 6171 7067 6177
rect 6328 6128 6334 6140
rect 7009 6137 7021 6171
rect 7055 6137 7067 6171
rect 7009 6131 7067 6137
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3970 6100 3976 6112
rect 3384 6072 3976 6100
rect 3384 6060 3390 6072
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9306 6100 9312 6112
rect 8904 6072 9312 6100
rect 8904 6060 8910 6072
rect 9306 6060 9312 6072
rect 9364 6100 9370 6112
rect 9950 6100 9956 6112
rect 9364 6072 9956 6100
rect 9364 6060 9370 6072
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 1104 6010 12788 6032
rect 1104 5958 2410 6010
rect 2462 5958 2474 6010
rect 2526 5958 2538 6010
rect 2590 5958 2602 6010
rect 2654 5958 2666 6010
rect 2718 5958 5331 6010
rect 5383 5958 5395 6010
rect 5447 5958 5459 6010
rect 5511 5958 5523 6010
rect 5575 5958 5587 6010
rect 5639 5958 8252 6010
rect 8304 5958 8316 6010
rect 8368 5958 8380 6010
rect 8432 5958 8444 6010
rect 8496 5958 8508 6010
rect 8560 5958 11173 6010
rect 11225 5958 11237 6010
rect 11289 5958 11301 6010
rect 11353 5958 11365 6010
rect 11417 5958 11429 6010
rect 11481 5958 12788 6010
rect 1104 5936 12788 5958
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 5810 5896 5816 5908
rect 3712 5868 5816 5896
rect 3712 5828 3740 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 5902 5856 5908 5908
rect 5960 5856 5966 5908
rect 6362 5856 6368 5908
rect 6420 5856 6426 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 7576 5868 9076 5896
rect 3160 5800 3740 5828
rect 3789 5831 3847 5837
rect 3160 5704 3188 5800
rect 3789 5797 3801 5831
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 5629 5831 5687 5837
rect 5629 5797 5641 5831
rect 5675 5828 5687 5831
rect 5675 5800 7328 5828
rect 5675 5797 5687 5800
rect 5629 5791 5687 5797
rect 3804 5760 3832 5791
rect 4430 5760 4436 5772
rect 3436 5732 3832 5760
rect 3988 5732 4436 5760
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1489 5695 1547 5701
rect 1489 5692 1501 5695
rect 1452 5664 1501 5692
rect 1452 5652 1458 5664
rect 1489 5661 1501 5664
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 3142 5652 3148 5704
rect 3200 5652 3206 5704
rect 3436 5701 3464 5732
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3988 5692 4016 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 7300 5769 7328 5800
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 4540 5732 6561 5760
rect 4540 5701 4568 5732
rect 6549 5729 6561 5732
rect 6595 5760 6607 5763
rect 7285 5763 7343 5769
rect 6595 5732 6776 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 3651 5664 4016 5692
rect 4065 5695 4123 5701
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4525 5655 4583 5661
rect 4632 5664 5457 5692
rect 1756 5627 1814 5633
rect 1756 5593 1768 5627
rect 1802 5624 1814 5627
rect 1946 5624 1952 5636
rect 1802 5596 1952 5624
rect 1802 5593 1814 5596
rect 1756 5587 1814 5593
rect 1946 5584 1952 5596
rect 2004 5584 2010 5636
rect 3694 5584 3700 5636
rect 3752 5624 3758 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3752 5596 3801 5624
rect 3752 5584 3758 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 4080 5624 4108 5655
rect 3789 5587 3847 5593
rect 3896 5596 4108 5624
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 3234 5556 3240 5568
rect 2915 5528 3240 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3602 5516 3608 5568
rect 3660 5556 3666 5568
rect 3896 5556 3924 5596
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 4632 5624 4660 5664
rect 5445 5661 5457 5664
rect 5491 5692 5503 5695
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5491 5664 5733 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 4396 5596 4660 5624
rect 4396 5584 4402 5596
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 5261 5627 5319 5633
rect 5261 5624 5273 5627
rect 4764 5596 5273 5624
rect 4764 5584 4770 5596
rect 5261 5593 5273 5596
rect 5307 5624 5319 5627
rect 5920 5624 5948 5655
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 6052 5664 6193 5692
rect 6052 5652 6058 5664
rect 6181 5661 6193 5664
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6748 5692 6776 5732
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 7374 5760 7380 5772
rect 7331 5732 7380 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 6748 5664 7481 5692
rect 6641 5655 6699 5661
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 5307 5596 5948 5624
rect 6656 5624 6684 5655
rect 6656 5596 6776 5624
rect 5307 5593 5319 5596
rect 5261 5587 5319 5593
rect 3660 5528 3924 5556
rect 3660 5516 3666 5528
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 4246 5556 4252 5568
rect 4203 5528 4252 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 6748 5556 6776 5596
rect 7190 5584 7196 5636
rect 7248 5584 7254 5636
rect 7576 5556 7604 5868
rect 7653 5831 7711 5837
rect 7653 5797 7665 5831
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 7668 5760 7696 5791
rect 8846 5760 8852 5772
rect 7668 5732 8852 5760
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9048 5760 9076 5868
rect 9122 5856 9128 5908
rect 9180 5856 9186 5908
rect 9398 5856 9404 5908
rect 9456 5856 9462 5908
rect 9585 5899 9643 5905
rect 9585 5865 9597 5899
rect 9631 5896 9643 5899
rect 9631 5868 10272 5896
rect 9631 5865 9643 5868
rect 9585 5859 9643 5865
rect 9140 5760 9168 5856
rect 8956 5732 9076 5760
rect 9114 5732 9168 5760
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8662 5692 8668 5704
rect 8527 5664 8668 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8956 5701 8984 5732
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 8179 5627 8237 5633
rect 8179 5593 8191 5627
rect 8225 5624 8237 5627
rect 8225 5593 8248 5624
rect 8179 5587 8248 5593
rect 5224 5528 7604 5556
rect 8220 5556 8248 5587
rect 8386 5584 8392 5636
rect 8444 5584 8450 5636
rect 9114 5633 9142 5732
rect 9416 5701 9444 5856
rect 10244 5760 10272 5868
rect 11514 5856 11520 5908
rect 11572 5856 11578 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 11940 5868 11989 5896
rect 11940 5856 11946 5868
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 11532 5760 11560 5856
rect 10244 5732 11560 5760
rect 9400 5695 9458 5701
rect 9400 5661 9412 5695
rect 9446 5661 9458 5695
rect 9400 5655 9458 5661
rect 9674 5652 9680 5704
rect 9732 5652 9738 5704
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 9079 5627 9142 5633
rect 9079 5593 9091 5627
rect 9125 5596 9142 5627
rect 9125 5593 9137 5596
rect 9079 5587 9137 5593
rect 9214 5584 9220 5636
rect 9272 5584 9278 5636
rect 9306 5584 9312 5636
rect 9364 5584 9370 5636
rect 9876 5624 9904 5655
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 10244 5701 10272 5732
rect 11606 5720 11612 5772
rect 11664 5720 11670 5772
rect 11992 5769 12020 5859
rect 11977 5763 12035 5769
rect 11977 5729 11989 5763
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10376 5664 10609 5692
rect 10376 5652 10382 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10827 5664 11161 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 10152 5624 10180 5652
rect 10796 5624 10824 5655
rect 9876 5596 10180 5624
rect 10428 5596 10824 5624
rect 11164 5624 11192 5655
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11624 5624 11652 5720
rect 11164 5596 11652 5624
rect 8570 5556 8576 5568
rect 8220 5528 8576 5556
rect 5224 5516 5230 5528
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 9861 5559 9919 5565
rect 9861 5525 9873 5559
rect 9907 5556 9919 5559
rect 10042 5556 10048 5568
rect 9907 5528 10048 5556
rect 9907 5525 9919 5528
rect 9861 5519 9919 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 10134 5516 10140 5568
rect 10192 5516 10198 5568
rect 10428 5565 10456 5596
rect 10413 5559 10471 5565
rect 10413 5525 10425 5559
rect 10459 5525 10471 5559
rect 10413 5519 10471 5525
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5556 10747 5559
rect 10962 5556 10968 5568
rect 10735 5528 10968 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 11992 5556 12020 5723
rect 12066 5652 12072 5704
rect 12124 5652 12130 5704
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 12437 5695 12495 5701
rect 12437 5692 12449 5695
rect 12216 5664 12449 5692
rect 12216 5652 12222 5664
rect 12437 5661 12449 5664
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 11572 5528 12449 5556
rect 11572 5516 11578 5528
rect 12437 5525 12449 5528
rect 12483 5525 12495 5559
rect 12437 5519 12495 5525
rect 1104 5466 12947 5488
rect 1104 5414 3870 5466
rect 3922 5414 3934 5466
rect 3986 5414 3998 5466
rect 4050 5414 4062 5466
rect 4114 5414 4126 5466
rect 4178 5414 6791 5466
rect 6843 5414 6855 5466
rect 6907 5414 6919 5466
rect 6971 5414 6983 5466
rect 7035 5414 7047 5466
rect 7099 5414 9712 5466
rect 9764 5414 9776 5466
rect 9828 5414 9840 5466
rect 9892 5414 9904 5466
rect 9956 5414 9968 5466
rect 10020 5414 12633 5466
rect 12685 5414 12697 5466
rect 12749 5414 12761 5466
rect 12813 5414 12825 5466
rect 12877 5414 12889 5466
rect 12941 5414 12947 5466
rect 1104 5392 12947 5414
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4488 5324 4997 5352
rect 4488 5312 4494 5324
rect 4985 5321 4997 5324
rect 5031 5321 5043 5355
rect 4985 5315 5043 5321
rect 5994 5312 6000 5364
rect 6052 5352 6058 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6052 5324 6561 5352
rect 6052 5312 6058 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 8294 5352 8300 5364
rect 7791 5324 8300 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 8266 5312 8300 5324
rect 8352 5312 8358 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 8478 5352 8484 5364
rect 8435 5324 8484 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 8478 5312 8484 5324
rect 8536 5352 8542 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 8536 5324 9689 5352
rect 8536 5312 8542 5324
rect 9677 5321 9689 5324
rect 9723 5352 9735 5355
rect 9766 5352 9772 5364
rect 9723 5324 9772 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 9766 5312 9772 5324
rect 9824 5352 9830 5364
rect 11514 5352 11520 5364
rect 9824 5324 11520 5352
rect 9824 5312 9830 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 12158 5352 12164 5364
rect 11747 5324 12164 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 4246 5284 4252 5296
rect 2639 5256 4252 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 6178 5284 6184 5296
rect 5092 5256 6184 5284
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 2179 5188 2237 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2372 5188 2421 5216
rect 2372 5176 2378 5188
rect 2409 5185 2421 5188
rect 2455 5216 2467 5219
rect 3510 5216 3516 5228
rect 2455 5188 3516 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 5092 5225 5120 5256
rect 6178 5244 6184 5256
rect 6236 5284 6242 5296
rect 6638 5284 6644 5296
rect 6236 5256 6644 5284
rect 6236 5244 6242 5256
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 7101 5287 7159 5293
rect 7101 5284 7113 5287
rect 6840 5256 7113 5284
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 4908 5148 4936 5179
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6656 5215 6684 5244
rect 6840 5225 6868 5256
rect 7101 5253 7113 5256
rect 7147 5284 7159 5287
rect 8266 5284 8294 5312
rect 9582 5284 9588 5296
rect 7147 5256 7604 5284
rect 8266 5256 9588 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 6825 5219 6883 5225
rect 6641 5209 6699 5215
rect 6641 5175 6653 5209
rect 6687 5175 6699 5209
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6825 5179 6883 5185
rect 6932 5188 7205 5216
rect 6641 5169 6699 5175
rect 4908 5120 5120 5148
rect 5092 5024 5120 5120
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 5736 5080 5764 5108
rect 6932 5080 6960 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7300 5148 7328 5179
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7576 5225 7604 5256
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 10152 5256 11621 5284
rect 10152 5228 10180 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7432 5188 7481 5216
rect 7432 5176 7438 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8662 5216 8668 5228
rect 8067 5188 8668 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 10042 5216 10048 5228
rect 9723 5188 10048 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10134 5176 10140 5228
rect 10192 5176 10198 5228
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10962 5216 10968 5228
rect 10735 5188 10968 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 7208 5120 7328 5148
rect 8389 5151 8447 5157
rect 7208 5092 7236 5120
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 8478 5148 8484 5160
rect 8435 5120 8484 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9398 5148 9404 5160
rect 9355 5120 9404 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 7006 5080 7012 5092
rect 5736 5052 7012 5080
rect 7006 5040 7012 5052
rect 7064 5040 7070 5092
rect 7190 5040 7196 5092
rect 7248 5040 7254 5092
rect 5074 4972 5080 5024
rect 5132 4972 5138 5024
rect 6730 4972 6736 5024
rect 6788 4972 6794 5024
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 10318 5012 10324 5024
rect 8628 4984 10324 5012
rect 8628 4972 8634 4984
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 10560 4984 10609 5012
rect 10560 4972 10566 4984
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 1104 4922 12788 4944
rect 1104 4870 2410 4922
rect 2462 4870 2474 4922
rect 2526 4870 2538 4922
rect 2590 4870 2602 4922
rect 2654 4870 2666 4922
rect 2718 4870 5331 4922
rect 5383 4870 5395 4922
rect 5447 4870 5459 4922
rect 5511 4870 5523 4922
rect 5575 4870 5587 4922
rect 5639 4870 8252 4922
rect 8304 4870 8316 4922
rect 8368 4870 8380 4922
rect 8432 4870 8444 4922
rect 8496 4870 8508 4922
rect 8560 4870 11173 4922
rect 11225 4870 11237 4922
rect 11289 4870 11301 4922
rect 11353 4870 11365 4922
rect 11417 4870 11429 4922
rect 11481 4870 12788 4922
rect 1104 4848 12788 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 3050 4808 3056 4820
rect 2823 4780 3056 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 3050 4768 3056 4780
rect 3108 4808 3114 4820
rect 3418 4808 3424 4820
rect 3108 4780 3424 4808
rect 3108 4768 3114 4780
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4706 4808 4712 4820
rect 4212 4780 4712 4808
rect 4212 4768 4218 4780
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5810 4768 5816 4820
rect 5868 4768 5874 4820
rect 6730 4808 6736 4820
rect 6012 4780 6736 4808
rect 3602 4740 3608 4752
rect 3252 4712 3608 4740
rect 3252 4681 3280 4712
rect 3602 4700 3608 4712
rect 3660 4740 3666 4752
rect 4433 4743 4491 4749
rect 4433 4740 4445 4743
rect 3660 4712 4445 4740
rect 3660 4700 3666 4712
rect 4433 4709 4445 4712
rect 4479 4740 4491 4743
rect 5534 4740 5540 4752
rect 4479 4712 5540 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 5828 4740 5856 4768
rect 5828 4712 5948 4740
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 3160 4604 3188 4635
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 3384 4644 3556 4672
rect 3384 4632 3390 4644
rect 3528 4616 3556 4644
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3752 4644 3985 4672
rect 3752 4632 3758 4644
rect 3973 4641 3985 4644
rect 4019 4672 4031 4675
rect 4019 4644 4752 4672
rect 4019 4641 4031 4644
rect 3973 4635 4031 4641
rect 3160 4576 3280 4604
rect 1664 4539 1722 4545
rect 1664 4505 1676 4539
rect 1710 4536 1722 4539
rect 2222 4536 2228 4548
rect 1710 4508 2228 4536
rect 1710 4505 1722 4508
rect 1664 4499 1722 4505
rect 2222 4496 2228 4508
rect 2280 4496 2286 4548
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 3252 4536 3280 4576
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3510 4564 3516 4616
rect 3568 4564 3574 4616
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 3786 4604 3792 4616
rect 3660 4576 3792 4604
rect 3660 4564 3666 4576
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4080 4536 4108 4567
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4724 4613 4752 4644
rect 4890 4632 4896 4684
rect 4948 4632 4954 4684
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5810 4672 5816 4684
rect 5031 4644 5816 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4908 4604 4936 4632
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4908 4576 5089 4604
rect 4709 4567 4767 4573
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 5920 4604 5948 4712
rect 6012 4613 6040 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7064 4780 7481 4808
rect 7064 4768 7070 4780
rect 7469 4777 7481 4780
rect 7515 4808 7527 4811
rect 8018 4808 8024 4820
rect 7515 4780 8024 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 8662 4808 8668 4820
rect 8312 4780 8668 4808
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8312 4672 8340 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9766 4768 9772 4820
rect 9824 4768 9830 4820
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 9784 4740 9812 4768
rect 8435 4712 9812 4740
rect 9861 4743 9919 4749
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 8067 4644 8340 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 5767 4576 5948 4604
rect 5997 4607 6055 4613
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 4356 4536 4384 4564
rect 3200 4508 3924 4536
rect 4080 4508 4384 4536
rect 3200 4496 3206 4508
rect 2958 4428 2964 4480
rect 3016 4428 3022 4480
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 3896 4468 3924 4508
rect 4617 4471 4675 4477
rect 4617 4468 4629 4471
rect 3896 4440 4629 4468
rect 4617 4437 4629 4440
rect 4663 4437 4675 4471
rect 4617 4431 4675 4437
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5169 4471 5227 4477
rect 5169 4468 5181 4471
rect 5132 4440 5181 4468
rect 5132 4428 5138 4440
rect 5169 4437 5181 4440
rect 5215 4437 5227 4471
rect 5276 4468 5304 4567
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 5537 4539 5595 4545
rect 5537 4505 5549 4539
rect 5583 4536 5595 4539
rect 6334 4539 6392 4545
rect 6334 4536 6346 4539
rect 5583 4508 6346 4536
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 6334 4505 6346 4508
rect 6380 4505 6392 4539
rect 6334 4499 6392 4505
rect 5626 4468 5632 4480
rect 5276 4440 5632 4468
rect 5169 4431 5227 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5902 4428 5908 4480
rect 5960 4428 5966 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8404 4477 8432 4703
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9324 4681 9352 4712
rect 9861 4709 9873 4743
rect 9907 4740 9919 4743
rect 10042 4740 10048 4752
rect 9907 4712 10048 4740
rect 9907 4709 9919 4712
rect 9861 4703 9919 4709
rect 9309 4675 9367 4681
rect 8720 4644 8800 4672
rect 8720 4632 8726 4644
rect 8570 4564 8576 4616
rect 8628 4564 8634 4616
rect 8772 4613 8800 4644
rect 9309 4641 9321 4675
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 9876 4672 9904 4703
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 10870 4700 10876 4752
rect 10928 4740 10934 4752
rect 11333 4743 11391 4749
rect 11333 4740 11345 4743
rect 10928 4712 11345 4740
rect 10928 4700 10934 4712
rect 11333 4709 11345 4712
rect 11379 4740 11391 4743
rect 12158 4740 12164 4752
rect 11379 4712 12164 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 9815 4644 9904 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 10502 4632 10508 4684
rect 10560 4672 10566 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10560 4644 10977 4672
rect 10560 4632 10566 4644
rect 10965 4641 10977 4644
rect 11011 4672 11023 4675
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11011 4644 11805 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11793 4641 11805 4644
rect 11839 4672 11851 4675
rect 12066 4672 12072 4684
rect 11839 4644 12072 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8803 4576 8953 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9456 4576 10241 4604
rect 9456 4564 9462 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 8665 4539 8723 4545
rect 8665 4505 8677 4539
rect 8711 4536 8723 4539
rect 9416 4536 9444 4564
rect 8711 4508 9444 4536
rect 8711 4505 8723 4508
rect 8665 4499 8723 4505
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 8352 4440 8401 4468
rect 8352 4428 8358 4440
rect 8389 4437 8401 4440
rect 8435 4437 8447 4471
rect 8389 4431 8447 4437
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 9582 4468 9588 4480
rect 9355 4440 9588 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 9582 4428 9588 4440
rect 9640 4468 9646 4480
rect 9766 4477 9772 4480
rect 9723 4471 9772 4477
rect 9723 4468 9735 4471
rect 9640 4440 9735 4468
rect 9640 4428 9646 4440
rect 9723 4437 9735 4440
rect 9769 4437 9772 4471
rect 9723 4431 9772 4437
rect 9766 4428 9772 4431
rect 9824 4468 9830 4480
rect 9861 4471 9919 4477
rect 9861 4468 9873 4471
rect 9824 4440 9873 4468
rect 9824 4428 9830 4440
rect 9861 4437 9873 4440
rect 9907 4468 9919 4471
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 9907 4440 10885 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 10873 4437 10885 4440
rect 10919 4468 10931 4471
rect 11333 4471 11391 4477
rect 11333 4468 11345 4471
rect 10919 4440 11345 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 11333 4437 11345 4440
rect 11379 4468 11391 4471
rect 11974 4468 11980 4480
rect 11379 4440 11980 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 11974 4428 11980 4440
rect 12032 4468 12038 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 12032 4440 12173 4468
rect 12032 4428 12038 4440
rect 12161 4437 12173 4440
rect 12207 4437 12219 4471
rect 12161 4431 12219 4437
rect 1104 4378 12947 4400
rect 1104 4326 3870 4378
rect 3922 4326 3934 4378
rect 3986 4326 3998 4378
rect 4050 4326 4062 4378
rect 4114 4326 4126 4378
rect 4178 4326 6791 4378
rect 6843 4326 6855 4378
rect 6907 4326 6919 4378
rect 6971 4326 6983 4378
rect 7035 4326 7047 4378
rect 7099 4326 9712 4378
rect 9764 4326 9776 4378
rect 9828 4326 9840 4378
rect 9892 4326 9904 4378
rect 9956 4326 9968 4378
rect 10020 4326 12633 4378
rect 12685 4326 12697 4378
rect 12749 4326 12761 4378
rect 12813 4326 12825 4378
rect 12877 4326 12889 4378
rect 12941 4326 12947 4378
rect 1104 4304 12947 4326
rect 2222 4224 2228 4276
rect 2280 4224 2286 4276
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 3200 4236 3249 4264
rect 3200 4224 3206 4236
rect 3237 4233 3249 4236
rect 3283 4233 3295 4267
rect 3237 4227 3295 4233
rect 3418 4224 3424 4276
rect 3476 4224 3482 4276
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 3752 4236 4077 4264
rect 3752 4224 3758 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 4065 4227 4123 4233
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 5902 4224 5908 4276
rect 5960 4224 5966 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 9677 4267 9735 4273
rect 9677 4264 9689 4267
rect 9640 4236 9689 4264
rect 9640 4224 9646 4236
rect 9677 4233 9689 4236
rect 9723 4264 9735 4267
rect 10226 4264 10232 4276
rect 9723 4236 10232 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 10226 4224 10232 4236
rect 10284 4264 10290 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10284 4236 10885 4264
rect 10284 4224 10290 4236
rect 10873 4233 10885 4236
rect 10919 4264 10931 4267
rect 11609 4267 11667 4273
rect 11609 4264 11621 4267
rect 10919 4236 11621 4264
rect 10919 4233 10931 4236
rect 10873 4227 10931 4233
rect 11609 4233 11621 4236
rect 11655 4233 11667 4267
rect 11609 4227 11667 4233
rect 12066 4224 12072 4276
rect 12124 4224 12130 4276
rect 3436 4196 3464 4224
rect 2516 4168 3096 4196
rect 3436 4168 3927 4196
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2516 4128 2544 4168
rect 2455 4100 2544 4128
rect 2593 4131 2651 4137
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2608 4060 2636 4091
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3068 4128 3096 4168
rect 3326 4128 3332 4140
rect 3068 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3436 4060 3464 4091
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3694 4128 3700 4140
rect 3568 4100 3700 4128
rect 3568 4088 3574 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3899 4137 3927 4168
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4126 3939 4131
rect 5077 4131 5135 4137
rect 3927 4098 4016 4126
rect 3927 4097 3939 4098
rect 3881 4091 3939 4097
rect 2608 4032 2774 4060
rect 3436 4032 3556 4060
rect 2746 3924 2774 4032
rect 3528 4004 3556 4032
rect 3602 4020 3608 4072
rect 3660 4020 3666 4072
rect 3988 4060 4016 4098
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5184 4128 5212 4224
rect 5123 4100 5212 4128
rect 5261 4131 5319 4137
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5552 4128 5580 4224
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5552 4100 5825 4128
rect 5261 4091 5319 4097
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8294 4128 8300 4140
rect 8067 4100 8300 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 5276 4060 5304 4091
rect 3988 4032 5304 4060
rect 3510 3952 3516 4004
rect 3568 3952 3574 4004
rect 3620 3992 3648 4020
rect 5626 3992 5632 4004
rect 3620 3964 5632 3992
rect 5626 3952 5632 3964
rect 5684 3992 5690 4004
rect 6012 3992 6040 4091
rect 5684 3964 6040 3992
rect 5684 3952 5690 3964
rect 3694 3924 3700 3936
rect 2746 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 5040 3896 5181 3924
rect 5040 3884 5046 3896
rect 5169 3893 5181 3896
rect 5215 3924 5227 3927
rect 5994 3924 6000 3936
rect 5215 3896 6000 3924
rect 5215 3893 5227 3896
rect 5169 3887 5227 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 8036 3933 8064 4091
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8662 4128 8668 4140
rect 8435 4100 8668 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 9398 4128 9404 4140
rect 9355 4100 9404 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 9677 4131 9735 4137
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 10042 4128 10048 4140
rect 9723 4100 10048 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 10962 4088 10968 4140
rect 11020 4088 11026 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12084 4128 12112 4224
rect 12023 4100 12112 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 10888 4060 10916 4088
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 10888 4032 11621 4060
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12216 4032 12449 4060
rect 12216 4020 12222 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 12176 3992 12204 4020
rect 11195 3964 12204 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 10318 3884 10324 3936
rect 10376 3884 10382 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 12032 3896 12081 3924
rect 12032 3884 12038 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 1104 3834 12788 3856
rect 1104 3782 2410 3834
rect 2462 3782 2474 3834
rect 2526 3782 2538 3834
rect 2590 3782 2602 3834
rect 2654 3782 2666 3834
rect 2718 3782 5331 3834
rect 5383 3782 5395 3834
rect 5447 3782 5459 3834
rect 5511 3782 5523 3834
rect 5575 3782 5587 3834
rect 5639 3782 8252 3834
rect 8304 3782 8316 3834
rect 8368 3782 8380 3834
rect 8432 3782 8444 3834
rect 8496 3782 8508 3834
rect 8560 3782 11173 3834
rect 11225 3782 11237 3834
rect 11289 3782 11301 3834
rect 11353 3782 11365 3834
rect 11417 3782 11429 3834
rect 11481 3782 12788 3834
rect 1104 3760 12788 3782
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 4890 3720 4896 3732
rect 3568 3692 4896 3720
rect 3568 3680 3574 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 4982 3680 4988 3732
rect 5040 3680 5046 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5132 3692 5641 3720
rect 5132 3680 5138 3692
rect 5629 3689 5641 3692
rect 5675 3720 5687 3723
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5675 3692 6009 3720
rect 5675 3689 5687 3692
rect 5629 3683 5687 3689
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 10318 3680 10324 3732
rect 10376 3680 10382 3732
rect 5000 3593 5028 3680
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 5224 3624 5764 3652
rect 5224 3612 5230 3624
rect 4985 3587 5043 3593
rect 4985 3553 4997 3587
rect 5031 3584 5043 3587
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5031 3556 5457 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5736 3584 5764 3624
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 6638 3652 6644 3664
rect 5868 3624 6644 3652
rect 5868 3612 5874 3624
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 10229 3655 10287 3661
rect 10229 3621 10241 3655
rect 10275 3652 10287 3655
rect 10336 3652 10364 3680
rect 10689 3655 10747 3661
rect 10689 3652 10701 3655
rect 10275 3624 10701 3652
rect 10275 3621 10287 3624
rect 10229 3615 10287 3621
rect 10689 3621 10701 3624
rect 10735 3652 10747 3655
rect 11054 3652 11060 3664
rect 10735 3624 11060 3652
rect 10735 3621 10747 3624
rect 10689 3615 10747 3621
rect 11054 3612 11060 3624
rect 11112 3652 11118 3664
rect 11149 3655 11207 3661
rect 11149 3652 11161 3655
rect 11112 3624 11161 3652
rect 11112 3612 11118 3624
rect 11149 3621 11161 3624
rect 11195 3652 11207 3655
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11195 3624 11621 3652
rect 11195 3621 11207 3624
rect 11149 3615 11207 3621
rect 11609 3621 11621 3624
rect 11655 3652 11667 3655
rect 12066 3652 12072 3664
rect 11655 3624 12072 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5736 3556 6101 3584
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4798 3516 4804 3528
rect 4663 3488 4804 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5629 3519 5687 3525
rect 5184 3488 5488 3516
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 5184 3448 5212 3488
rect 3752 3420 5212 3448
rect 3752 3408 3758 3420
rect 5350 3408 5356 3460
rect 5408 3408 5414 3460
rect 5460 3448 5488 3488
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 5736 3516 5764 3556
rect 6089 3553 6101 3556
rect 6135 3584 6147 3587
rect 6178 3584 6184 3596
rect 6135 3556 6184 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 9907 3556 10333 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 10321 3553 10333 3556
rect 10367 3584 10379 3587
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 10367 3556 10793 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10781 3553 10793 3556
rect 10827 3584 10839 3587
rect 11238 3584 11244 3596
rect 10827 3556 11244 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 11238 3544 11244 3556
rect 11296 3584 11302 3596
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11296 3556 11713 3584
rect 11296 3544 11302 3556
rect 11701 3553 11713 3556
rect 11747 3584 11759 3587
rect 12158 3584 12164 3596
rect 11747 3556 12164 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 5675 3488 5764 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 5994 3476 6000 3528
rect 6052 3476 6058 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 5460 3420 6408 3448
rect 5258 3340 5264 3392
rect 5316 3340 5322 3392
rect 5810 3340 5816 3392
rect 5868 3340 5874 3392
rect 6380 3389 6408 3420
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3349 6423 3383
rect 6365 3343 6423 3349
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 7374 3380 7380 3392
rect 6604 3352 7380 3380
rect 6604 3340 6610 3352
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 10244 3389 10272 3476
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3380 10287 3383
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 10275 3352 10701 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 10689 3349 10701 3352
rect 10735 3380 10747 3383
rect 10778 3380 10784 3392
rect 10735 3352 10784 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 10778 3340 10784 3352
rect 10836 3380 10842 3392
rect 11149 3383 11207 3389
rect 11149 3380 11161 3383
rect 10836 3352 11161 3380
rect 10836 3340 10842 3352
rect 11149 3349 11161 3352
rect 11195 3380 11207 3383
rect 11609 3383 11667 3389
rect 11609 3380 11621 3383
rect 11195 3352 11621 3380
rect 11195 3349 11207 3352
rect 11149 3343 11207 3349
rect 11609 3349 11621 3352
rect 11655 3380 11667 3383
rect 12069 3383 12127 3389
rect 12069 3380 12081 3383
rect 11655 3352 12081 3380
rect 11655 3349 11667 3352
rect 11609 3343 11667 3349
rect 12069 3349 12081 3352
rect 12115 3349 12127 3383
rect 12069 3343 12127 3349
rect 1104 3290 12947 3312
rect 1104 3238 3870 3290
rect 3922 3238 3934 3290
rect 3986 3238 3998 3290
rect 4050 3238 4062 3290
rect 4114 3238 4126 3290
rect 4178 3238 6791 3290
rect 6843 3238 6855 3290
rect 6907 3238 6919 3290
rect 6971 3238 6983 3290
rect 7035 3238 7047 3290
rect 7099 3238 9712 3290
rect 9764 3238 9776 3290
rect 9828 3238 9840 3290
rect 9892 3238 9904 3290
rect 9956 3238 9968 3290
rect 10020 3238 12633 3290
rect 12685 3238 12697 3290
rect 12749 3238 12761 3290
rect 12813 3238 12825 3290
rect 12877 3238 12889 3290
rect 12941 3238 12947 3290
rect 1104 3216 12947 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3145 2007 3179
rect 3694 3176 3700 3188
rect 1949 3139 2007 3145
rect 2746 3148 3700 3176
rect 1964 3108 1992 3139
rect 2041 3111 2099 3117
rect 2041 3108 2053 3111
rect 1964 3080 2053 3108
rect 2041 3077 2053 3080
rect 2087 3077 2099 3111
rect 2746 3108 2774 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 4338 3176 4344 3188
rect 3927 3148 4344 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 3988 3117 4016 3148
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4798 3176 4804 3188
rect 4571 3148 4804 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5350 3176 5356 3188
rect 5031 3148 5356 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 6089 3179 6147 3185
rect 6089 3145 6101 3179
rect 6135 3176 6147 3179
rect 6362 3176 6368 3188
rect 6135 3148 6368 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 9049 3179 9107 3185
rect 9049 3176 9061 3179
rect 6696 3148 9061 3176
rect 6696 3136 6702 3148
rect 2041 3071 2099 3077
rect 2148 3080 2774 3108
rect 3973 3111 4031 3117
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1596 2904 1624 3003
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2148 2972 2176 3080
rect 3973 3077 3985 3111
rect 4019 3077 4031 3111
rect 3973 3071 4031 3077
rect 4246 3068 4252 3120
rect 4304 3108 4310 3120
rect 5813 3111 5871 3117
rect 5813 3108 5825 3111
rect 4304 3080 5825 3108
rect 4304 3068 4310 3080
rect 5813 3077 5825 3080
rect 5859 3108 5871 3111
rect 5859 3080 6684 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2768 3043 2826 3049
rect 2768 3009 2780 3043
rect 2814 3040 2826 3043
rect 3142 3040 3148 3052
rect 2814 3012 3148 3040
rect 2814 3009 2826 3012
rect 2768 3003 2826 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 1719 2944 2176 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2501 2975 2559 2981
rect 2501 2972 2513 2975
rect 2372 2944 2513 2972
rect 2372 2932 2378 2944
rect 2501 2941 2513 2944
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 1596 2876 2544 2904
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 2409 2839 2467 2845
rect 2409 2836 2421 2839
rect 2188 2808 2421 2836
rect 2188 2796 2194 2808
rect 2409 2805 2421 2808
rect 2455 2805 2467 2839
rect 2516 2836 2544 2876
rect 2774 2836 2780 2848
rect 2516 2808 2780 2836
rect 2409 2799 2467 2805
rect 2774 2796 2780 2808
rect 2832 2836 2838 2848
rect 4172 2836 4200 3003
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 4706 3000 4712 3052
rect 4764 3040 4770 3052
rect 6656 3049 6684 3080
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4764 3012 4813 3040
rect 4764 3000 4770 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6227 3012 6377 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6365 3009 6377 3012
rect 6411 3040 6423 3043
rect 6641 3043 6699 3049
rect 6411 3012 6592 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 4356 2904 4384 3000
rect 4448 2972 4476 3000
rect 5000 2972 5028 3003
rect 4448 2944 5028 2972
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2972 6055 2975
rect 6457 2975 6515 2981
rect 6457 2972 6469 2975
rect 6043 2944 6469 2972
rect 6043 2941 6055 2944
rect 5997 2935 6055 2941
rect 6457 2941 6469 2944
rect 6503 2941 6515 2975
rect 6564 2972 6592 3012
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6748 3040 6776 3148
rect 9049 3145 9061 3148
rect 9095 3145 9107 3179
rect 9049 3139 9107 3145
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3145 9275 3179
rect 9217 3139 9275 3145
rect 6822 3068 6828 3120
rect 6880 3108 6886 3120
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 6880 3080 7113 3108
rect 6880 3068 6886 3080
rect 7101 3077 7113 3080
rect 7147 3108 7159 3111
rect 8846 3108 8852 3120
rect 7147 3080 8852 3108
rect 7147 3077 7159 3080
rect 7101 3071 7159 3077
rect 8846 3068 8852 3080
rect 8904 3068 8910 3120
rect 9232 3108 9260 3139
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 10836 3148 11345 3176
rect 10836 3136 10842 3148
rect 11333 3145 11345 3148
rect 11379 3176 11391 3179
rect 11698 3176 11704 3188
rect 11379 3148 11704 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11698 3136 11704 3148
rect 11756 3176 11762 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11756 3148 12081 3176
rect 11756 3136 11762 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 12069 3139 12127 3145
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 9232 3080 9413 3108
rect 9401 3077 9413 3080
rect 9447 3077 9459 3111
rect 9401 3071 9459 3077
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6748 3012 7021 3040
rect 6641 3003 6699 3009
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7300 2972 7328 3003
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 7633 3043 7691 3049
rect 7633 3040 7645 3043
rect 7524 3012 7645 3040
rect 7524 3000 7530 3012
rect 7633 3009 7645 3012
rect 7679 3009 7691 3043
rect 7633 3003 7691 3009
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11054 3040 11060 3052
rect 10827 3012 11060 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 11112 3012 11345 3040
rect 11112 3000 11118 3012
rect 11333 3009 11345 3012
rect 11379 3040 11391 3043
rect 11606 3040 11612 3052
rect 11379 3012 11612 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11606 3000 11612 3012
rect 11664 3040 11670 3052
rect 12069 3043 12127 3049
rect 12069 3040 12081 3043
rect 11664 3012 12081 3040
rect 11664 3000 11670 3012
rect 12069 3009 12081 3012
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 6564 2944 7328 2972
rect 6457 2935 6515 2941
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 4356 2876 5917 2904
rect 5905 2873 5917 2876
rect 5951 2904 5963 2907
rect 6178 2904 6184 2916
rect 5951 2876 6184 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 6178 2864 6184 2876
rect 6236 2904 6242 2916
rect 6472 2904 6500 2935
rect 6638 2904 6644 2916
rect 6236 2876 6408 2904
rect 6472 2876 6644 2904
rect 6236 2864 6242 2876
rect 4706 2836 4712 2848
rect 2832 2808 4712 2836
rect 2832 2796 2838 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6380 2845 6408 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7190 2904 7196 2916
rect 6871 2876 7196 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7300 2904 7328 2944
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 10459 2944 10977 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 10965 2941 10977 2944
rect 11011 2972 11023 2975
rect 11238 2972 11244 2984
rect 11011 2944 11244 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11238 2932 11244 2944
rect 11296 2972 11302 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11296 2944 11713 2972
rect 11296 2932 11302 2944
rect 11701 2941 11713 2944
rect 11747 2972 11759 2975
rect 11790 2972 11796 2984
rect 11747 2944 11796 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 7300 2876 7420 2904
rect 6365 2839 6423 2845
rect 6365 2805 6377 2839
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 7282 2796 7288 2848
rect 7340 2796 7346 2848
rect 7392 2836 7420 2876
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 7392 2808 8769 2836
rect 8757 2805 8769 2808
rect 8803 2836 8815 2839
rect 9033 2839 9091 2845
rect 9033 2836 9045 2839
rect 8803 2808 9045 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 9033 2805 9045 2808
rect 9079 2805 9091 2839
rect 9033 2799 9091 2805
rect 9490 2796 9496 2848
rect 9548 2796 9554 2848
rect 1104 2746 12788 2768
rect 1104 2694 2410 2746
rect 2462 2694 2474 2746
rect 2526 2694 2538 2746
rect 2590 2694 2602 2746
rect 2654 2694 2666 2746
rect 2718 2694 5331 2746
rect 5383 2694 5395 2746
rect 5447 2694 5459 2746
rect 5511 2694 5523 2746
rect 5575 2694 5587 2746
rect 5639 2694 8252 2746
rect 8304 2694 8316 2746
rect 8368 2694 8380 2746
rect 8432 2694 8444 2746
rect 8496 2694 8508 2746
rect 8560 2694 11173 2746
rect 11225 2694 11237 2746
rect 11289 2694 11301 2746
rect 11353 2694 11365 2746
rect 11417 2694 11429 2746
rect 11481 2694 12788 2746
rect 1104 2672 12788 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2866 2632 2872 2644
rect 1627 2604 2872 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3142 2592 3148 2644
rect 3200 2592 3206 2644
rect 7466 2592 7472 2644
rect 7524 2592 7530 2644
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 3344 2536 7205 2564
rect 3344 2440 3372 2536
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 7193 2527 7251 2533
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 11664 2536 11713 2564
rect 11664 2524 11670 2536
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 4338 2456 4344 2508
rect 4396 2456 4402 2508
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 4488 2468 5120 2496
rect 4488 2456 4494 2468
rect 750 2388 756 2440
rect 808 2428 814 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 808 2400 1409 2428
rect 808 2388 814 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2130 2428 2136 2440
rect 1903 2400 2136 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3786 2428 3792 2440
rect 3651 2400 3792 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4356 2428 4384 2456
rect 5092 2437 5120 2468
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11848 2468 12081 2496
rect 11848 2456 11854 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4356 2400 4813 2428
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5828 2428 5856 2456
rect 5123 2400 5856 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 2464 2332 4660 2360
rect 2464 2320 2470 2332
rect 4632 2304 4660 2332
rect 4706 2320 4712 2372
rect 4764 2360 4770 2372
rect 4908 2360 4936 2391
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7340 2400 7481 2428
rect 7340 2388 7346 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 8570 2428 8576 2440
rect 7699 2400 8576 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8570 2388 8576 2400
rect 8628 2428 8634 2440
rect 9490 2428 9496 2440
rect 8628 2400 9496 2428
rect 8628 2388 8634 2400
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 4764 2332 4936 2360
rect 4764 2320 4770 2332
rect 1670 2252 1676 2304
rect 1728 2252 1734 2304
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 4430 2292 4436 2304
rect 3559 2264 4436 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 4614 2252 4620 2304
rect 4672 2252 4678 2304
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 11716 2301 11744 2388
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4856 2264 4905 2292
rect 4856 2252 4862 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 1104 2202 12947 2224
rect 1104 2150 3870 2202
rect 3922 2150 3934 2202
rect 3986 2150 3998 2202
rect 4050 2150 4062 2202
rect 4114 2150 4126 2202
rect 4178 2150 6791 2202
rect 6843 2150 6855 2202
rect 6907 2150 6919 2202
rect 6971 2150 6983 2202
rect 7035 2150 7047 2202
rect 7099 2150 9712 2202
rect 9764 2150 9776 2202
rect 9828 2150 9840 2202
rect 9892 2150 9904 2202
rect 9956 2150 9968 2202
rect 10020 2150 12633 2202
rect 12685 2150 12697 2202
rect 12749 2150 12761 2202
rect 12813 2150 12825 2202
rect 12877 2150 12889 2202
rect 12941 2150 12947 2202
rect 1104 2128 12947 2150
rect 2038 2088 2044 2100
rect 1688 2060 2044 2088
rect 1688 1961 1716 2060
rect 2038 2048 2044 2060
rect 2096 2048 2102 2100
rect 2866 2048 2872 2100
rect 2924 2048 2930 2100
rect 3697 2091 3755 2097
rect 3697 2057 3709 2091
rect 3743 2088 3755 2091
rect 4246 2088 4252 2100
rect 3743 2060 4252 2088
rect 3743 2057 3755 2060
rect 3697 2051 3755 2057
rect 2884 2020 2912 2048
rect 1964 1992 2912 2020
rect 1964 1961 1992 1992
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 1949 1955 2007 1961
rect 1949 1921 1961 1955
rect 1995 1921 2007 1955
rect 1949 1915 2007 1921
rect 2317 1955 2375 1961
rect 2317 1921 2329 1955
rect 2363 1952 2375 1955
rect 2406 1952 2412 1964
rect 2363 1924 2412 1952
rect 2363 1921 2375 1924
rect 2317 1915 2375 1921
rect 1394 1776 1400 1828
rect 1452 1816 1458 1828
rect 1489 1819 1547 1825
rect 1489 1816 1501 1819
rect 1452 1788 1501 1816
rect 1452 1776 1458 1788
rect 1489 1785 1501 1788
rect 1535 1816 1547 1819
rect 2332 1816 2360 1915
rect 2406 1912 2412 1924
rect 2464 1912 2470 1964
rect 2584 1955 2642 1961
rect 2584 1921 2596 1955
rect 2630 1952 2642 1955
rect 3142 1952 3148 1964
rect 2630 1924 3148 1952
rect 2630 1921 2642 1924
rect 2584 1915 2642 1921
rect 3142 1912 3148 1924
rect 3200 1912 3206 1964
rect 3804 1893 3832 2060
rect 4246 2048 4252 2060
rect 4304 2048 4310 2100
rect 4706 2088 4712 2100
rect 4540 2060 4712 2088
rect 4540 2029 4568 2060
rect 4706 2048 4712 2060
rect 4764 2048 4770 2100
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 4948 2060 5120 2088
rect 4948 2048 4954 2060
rect 5092 2029 5120 2060
rect 6178 2048 6184 2100
rect 6236 2048 6242 2100
rect 7193 2091 7251 2097
rect 7193 2057 7205 2091
rect 7239 2088 7251 2091
rect 7239 2060 7420 2088
rect 7239 2057 7251 2060
rect 7193 2051 7251 2057
rect 4525 2023 4583 2029
rect 4525 2020 4537 2023
rect 4264 1992 4537 2020
rect 4264 1961 4292 1992
rect 4525 1989 4537 1992
rect 4571 1989 4583 2023
rect 4525 1983 4583 1989
rect 5068 2023 5126 2029
rect 5068 1989 5080 2023
rect 5114 1989 5126 2023
rect 5994 2020 6000 2032
rect 5068 1983 5126 1989
rect 5920 1992 6000 2020
rect 4065 1955 4123 1961
rect 4065 1921 4077 1955
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 4341 1955 4399 1961
rect 4341 1921 4353 1955
rect 4387 1952 4399 1955
rect 4430 1952 4436 1964
rect 4387 1924 4436 1952
rect 4387 1921 4399 1924
rect 4341 1915 4399 1921
rect 3789 1887 3847 1893
rect 3789 1853 3801 1887
rect 3835 1853 3847 1887
rect 4080 1884 4108 1915
rect 4356 1884 4384 1915
rect 4430 1912 4436 1924
rect 4488 1912 4494 1964
rect 4706 1912 4712 1964
rect 4764 1952 4770 1964
rect 4801 1955 4859 1961
rect 4801 1952 4813 1955
rect 4764 1924 4813 1952
rect 4764 1912 4770 1924
rect 4801 1921 4813 1924
rect 4847 1952 4859 1955
rect 5920 1952 5948 1992
rect 5994 1980 6000 1992
rect 6052 2020 6058 2032
rect 7392 2020 7420 2060
rect 8662 2048 8668 2100
rect 8720 2048 8726 2100
rect 7530 2023 7588 2029
rect 7530 2020 7542 2023
rect 6052 1992 7328 2020
rect 7392 1992 7542 2020
rect 6052 1980 6058 1992
rect 4847 1924 5948 1952
rect 6549 1955 6607 1961
rect 4847 1921 4859 1924
rect 4801 1915 4859 1921
rect 6549 1921 6561 1955
rect 6595 1952 6607 1955
rect 6638 1952 6644 1964
rect 6595 1924 6644 1952
rect 6595 1921 6607 1924
rect 6549 1915 6607 1921
rect 6638 1912 6644 1924
rect 6696 1912 6702 1964
rect 7006 1912 7012 1964
rect 7064 1912 7070 1964
rect 7300 1961 7328 1992
rect 7530 1989 7542 1992
rect 7576 1989 7588 2023
rect 7530 1983 7588 1989
rect 7285 1955 7343 1961
rect 7285 1921 7297 1955
rect 7331 1921 7343 1955
rect 7285 1915 7343 1921
rect 6457 1887 6515 1893
rect 6457 1884 6469 1887
rect 4080 1856 4384 1884
rect 5828 1856 6469 1884
rect 3789 1847 3847 1853
rect 1535 1788 2360 1816
rect 3344 1788 4844 1816
rect 1535 1785 1547 1788
rect 1489 1779 1547 1785
rect 2133 1751 2191 1757
rect 2133 1717 2145 1751
rect 2179 1748 2191 1751
rect 2222 1748 2228 1760
rect 2179 1720 2228 1748
rect 2179 1717 2191 1720
rect 2133 1711 2191 1717
rect 2222 1708 2228 1720
rect 2280 1748 2286 1760
rect 3344 1748 3372 1788
rect 2280 1720 3372 1748
rect 2280 1708 2286 1720
rect 3878 1708 3884 1760
rect 3936 1748 3942 1760
rect 4065 1751 4123 1757
rect 4065 1748 4077 1751
rect 3936 1720 4077 1748
rect 3936 1708 3942 1720
rect 4065 1717 4077 1720
rect 4111 1717 4123 1751
rect 4065 1711 4123 1717
rect 4706 1708 4712 1760
rect 4764 1708 4770 1760
rect 4816 1748 4844 1788
rect 4982 1748 4988 1760
rect 4816 1720 4988 1748
rect 4982 1708 4988 1720
rect 5040 1708 5046 1760
rect 5166 1708 5172 1760
rect 5224 1748 5230 1760
rect 5828 1748 5856 1856
rect 6457 1853 6469 1856
rect 6503 1853 6515 1887
rect 6457 1847 6515 1853
rect 6914 1776 6920 1828
rect 6972 1776 6978 1828
rect 5224 1720 5856 1748
rect 5224 1708 5230 1720
rect 1104 1658 12788 1680
rect 1104 1606 2410 1658
rect 2462 1606 2474 1658
rect 2526 1606 2538 1658
rect 2590 1606 2602 1658
rect 2654 1606 2666 1658
rect 2718 1606 5331 1658
rect 5383 1606 5395 1658
rect 5447 1606 5459 1658
rect 5511 1606 5523 1658
rect 5575 1606 5587 1658
rect 5639 1606 8252 1658
rect 8304 1606 8316 1658
rect 8368 1606 8380 1658
rect 8432 1606 8444 1658
rect 8496 1606 8508 1658
rect 8560 1606 11173 1658
rect 11225 1606 11237 1658
rect 11289 1606 11301 1658
rect 11353 1606 11365 1658
rect 11417 1606 11429 1658
rect 11481 1606 12788 1658
rect 1104 1584 12788 1606
rect 2038 1504 2044 1556
rect 2096 1544 2102 1556
rect 2096 1516 2636 1544
rect 2096 1504 2102 1516
rect 1394 1368 1400 1420
rect 1452 1368 1458 1420
rect 2608 1408 2636 1516
rect 2774 1504 2780 1556
rect 2832 1504 2838 1556
rect 3142 1504 3148 1556
rect 3200 1504 3206 1556
rect 4890 1504 4896 1556
rect 4948 1544 4954 1556
rect 5261 1547 5319 1553
rect 5261 1544 5273 1547
rect 4948 1516 5273 1544
rect 4948 1504 4954 1516
rect 5261 1513 5273 1516
rect 5307 1513 5319 1547
rect 5261 1507 5319 1513
rect 7006 1504 7012 1556
rect 7064 1544 7070 1556
rect 7377 1547 7435 1553
rect 7377 1544 7389 1547
rect 7064 1516 7389 1544
rect 7064 1504 7070 1516
rect 7377 1513 7389 1516
rect 7423 1513 7435 1547
rect 7377 1507 7435 1513
rect 3344 1448 5120 1476
rect 2608 1380 2820 1408
rect 1670 1349 1676 1352
rect 1664 1340 1676 1349
rect 1631 1312 1676 1340
rect 1664 1303 1676 1312
rect 1670 1300 1676 1303
rect 1728 1300 1734 1352
rect 2792 1272 2820 1380
rect 3344 1352 3372 1448
rect 3878 1408 3884 1420
rect 3620 1380 3884 1408
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 3620 1349 3648 1380
rect 3878 1368 3884 1380
rect 3936 1368 3942 1420
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1309 3663 1343
rect 3605 1303 3663 1309
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 4080 1272 4108 1303
rect 4706 1300 4712 1352
rect 4764 1300 4770 1352
rect 4798 1300 4804 1352
rect 4856 1300 4862 1352
rect 5092 1349 5120 1448
rect 5184 1448 7236 1476
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1309 5135 1343
rect 5077 1303 5135 1309
rect 2792 1244 4108 1272
rect 4724 1272 4752 1300
rect 4893 1275 4951 1281
rect 4893 1272 4905 1275
rect 4724 1244 4905 1272
rect 4893 1241 4905 1244
rect 4939 1241 4951 1275
rect 4893 1235 4951 1241
rect 4982 1232 4988 1284
rect 5040 1272 5046 1284
rect 5184 1272 5212 1448
rect 6914 1300 6920 1352
rect 6972 1340 6978 1352
rect 7208 1349 7236 1448
rect 7009 1343 7067 1349
rect 7009 1340 7021 1343
rect 6972 1312 7021 1340
rect 6972 1300 6978 1312
rect 7009 1309 7021 1312
rect 7055 1309 7067 1343
rect 7009 1303 7067 1309
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 5040 1244 5212 1272
rect 5040 1232 5046 1244
rect 3513 1207 3571 1213
rect 3513 1173 3525 1207
rect 3559 1204 3571 1207
rect 5166 1204 5172 1216
rect 3559 1176 5172 1204
rect 3559 1173 3571 1176
rect 3513 1167 3571 1173
rect 5166 1164 5172 1176
rect 5224 1164 5230 1216
rect 1104 1114 12947 1136
rect 1104 1062 3870 1114
rect 3922 1062 3934 1114
rect 3986 1062 3998 1114
rect 4050 1062 4062 1114
rect 4114 1062 4126 1114
rect 4178 1062 6791 1114
rect 6843 1062 6855 1114
rect 6907 1062 6919 1114
rect 6971 1062 6983 1114
rect 7035 1062 7047 1114
rect 7099 1062 9712 1114
rect 9764 1062 9776 1114
rect 9828 1062 9840 1114
rect 9892 1062 9904 1114
rect 9956 1062 9968 1114
rect 10020 1062 12633 1114
rect 12685 1062 12697 1114
rect 12749 1062 12761 1114
rect 12813 1062 12825 1114
rect 12877 1062 12889 1114
rect 12941 1062 12947 1114
rect 1104 1040 12947 1062
<< via1 >>
rect 2410 12486 2462 12538
rect 2474 12486 2526 12538
rect 2538 12486 2590 12538
rect 2602 12486 2654 12538
rect 2666 12486 2718 12538
rect 5331 12486 5383 12538
rect 5395 12486 5447 12538
rect 5459 12486 5511 12538
rect 5523 12486 5575 12538
rect 5587 12486 5639 12538
rect 8252 12486 8304 12538
rect 8316 12486 8368 12538
rect 8380 12486 8432 12538
rect 8444 12486 8496 12538
rect 8508 12486 8560 12538
rect 11173 12486 11225 12538
rect 11237 12486 11289 12538
rect 11301 12486 11353 12538
rect 11365 12486 11417 12538
rect 11429 12486 11481 12538
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 5816 12248 5868 12300
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 1308 12112 1360 12164
rect 3516 12155 3568 12164
rect 3516 12121 3525 12155
rect 3525 12121 3559 12155
rect 3559 12121 3568 12155
rect 3516 12112 3568 12121
rect 5540 12112 5592 12164
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6460 12223 6512 12232
rect 6460 12189 6475 12223
rect 6475 12189 6509 12223
rect 6509 12189 6512 12223
rect 6460 12180 6512 12189
rect 6092 12112 6144 12164
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 10048 12180 10100 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 8944 12044 8996 12096
rect 3870 11942 3922 11994
rect 3934 11942 3986 11994
rect 3998 11942 4050 11994
rect 4062 11942 4114 11994
rect 4126 11942 4178 11994
rect 6791 11942 6843 11994
rect 6855 11942 6907 11994
rect 6919 11942 6971 11994
rect 6983 11942 7035 11994
rect 7047 11942 7099 11994
rect 9712 11942 9764 11994
rect 9776 11942 9828 11994
rect 9840 11942 9892 11994
rect 9904 11942 9956 11994
rect 9968 11942 10020 11994
rect 12633 11942 12685 11994
rect 12697 11942 12749 11994
rect 12761 11942 12813 11994
rect 12825 11942 12877 11994
rect 12889 11942 12941 11994
rect 3516 11840 3568 11892
rect 5540 11840 5592 11892
rect 5632 11840 5684 11892
rect 5816 11840 5868 11892
rect 6184 11840 6236 11892
rect 8392 11840 8444 11892
rect 10048 11840 10100 11892
rect 10324 11840 10376 11892
rect 10600 11840 10652 11892
rect 10876 11840 10928 11892
rect 11152 11840 11204 11892
rect 3792 11704 3844 11756
rect 1308 11500 1360 11552
rect 3516 11500 3568 11552
rect 4344 11636 4396 11688
rect 6460 11636 6512 11688
rect 6736 11704 6788 11756
rect 8852 11745 8904 11756
rect 8852 11711 8861 11745
rect 8861 11711 8895 11745
rect 8895 11711 8904 11745
rect 8852 11704 8904 11711
rect 8944 11747 8996 11756
rect 8944 11713 8976 11747
rect 8976 11713 8996 11747
rect 8944 11704 8996 11713
rect 4436 11611 4488 11620
rect 4436 11577 4445 11611
rect 4445 11577 4479 11611
rect 4479 11577 4488 11611
rect 4436 11568 4488 11577
rect 8944 11568 8996 11620
rect 6092 11500 6144 11552
rect 8852 11500 8904 11552
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 11888 11500 11940 11552
rect 2410 11398 2462 11450
rect 2474 11398 2526 11450
rect 2538 11398 2590 11450
rect 2602 11398 2654 11450
rect 2666 11398 2718 11450
rect 5331 11398 5383 11450
rect 5395 11398 5447 11450
rect 5459 11398 5511 11450
rect 5523 11398 5575 11450
rect 5587 11398 5639 11450
rect 8252 11398 8304 11450
rect 8316 11398 8368 11450
rect 8380 11398 8432 11450
rect 8444 11398 8496 11450
rect 8508 11398 8560 11450
rect 11173 11398 11225 11450
rect 11237 11398 11289 11450
rect 11301 11398 11353 11450
rect 11365 11398 11417 11450
rect 11429 11398 11481 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4436 11296 4488 11348
rect 6736 11296 6788 11348
rect 1308 11092 1360 11144
rect 1492 11092 1544 11144
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 3792 11092 3844 11144
rect 2596 11024 2648 11076
rect 4344 11092 4396 11144
rect 11520 11160 11572 11212
rect 11980 11160 12032 11212
rect 5816 11092 5868 11144
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 5172 11024 5224 11076
rect 2320 10956 2372 11008
rect 4528 10999 4580 11008
rect 4528 10965 4537 10999
rect 4537 10965 4571 10999
rect 4571 10965 4580 10999
rect 4528 10956 4580 10965
rect 7288 10956 7340 11008
rect 10232 10956 10284 11008
rect 11888 10956 11940 11008
rect 3870 10854 3922 10906
rect 3934 10854 3986 10906
rect 3998 10854 4050 10906
rect 4062 10854 4114 10906
rect 4126 10854 4178 10906
rect 6791 10854 6843 10906
rect 6855 10854 6907 10906
rect 6919 10854 6971 10906
rect 6983 10854 7035 10906
rect 7047 10854 7099 10906
rect 9712 10854 9764 10906
rect 9776 10854 9828 10906
rect 9840 10854 9892 10906
rect 9904 10854 9956 10906
rect 9968 10854 10020 10906
rect 12633 10854 12685 10906
rect 12697 10854 12749 10906
rect 12761 10854 12813 10906
rect 12825 10854 12877 10906
rect 12889 10854 12941 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2228 10752 2280 10804
rect 2596 10795 2648 10804
rect 2596 10761 2605 10795
rect 2605 10761 2639 10795
rect 2639 10761 2648 10795
rect 2596 10752 2648 10761
rect 6368 10752 6420 10804
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 1768 10616 1820 10668
rect 2964 10684 3016 10736
rect 6092 10727 6144 10736
rect 6092 10693 6101 10727
rect 6101 10693 6135 10727
rect 6135 10693 6144 10727
rect 6092 10684 6144 10693
rect 6920 10684 6972 10736
rect 2228 10616 2280 10668
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 3148 10616 3200 10668
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 4344 10616 4396 10668
rect 3516 10412 3568 10464
rect 4620 10412 4672 10464
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 5816 10548 5868 10600
rect 4988 10412 5040 10464
rect 7564 10659 7616 10668
rect 7564 10625 7598 10659
rect 7598 10625 7616 10659
rect 7564 10616 7616 10625
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 10048 10684 10100 10736
rect 10232 10684 10284 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 10048 10548 10100 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 9772 10523 9824 10532
rect 9772 10489 9781 10523
rect 9781 10489 9815 10523
rect 9815 10489 9824 10523
rect 9772 10480 9824 10489
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 10232 10412 10284 10464
rect 2410 10310 2462 10362
rect 2474 10310 2526 10362
rect 2538 10310 2590 10362
rect 2602 10310 2654 10362
rect 2666 10310 2718 10362
rect 5331 10310 5383 10362
rect 5395 10310 5447 10362
rect 5459 10310 5511 10362
rect 5523 10310 5575 10362
rect 5587 10310 5639 10362
rect 8252 10310 8304 10362
rect 8316 10310 8368 10362
rect 8380 10310 8432 10362
rect 8444 10310 8496 10362
rect 8508 10310 8560 10362
rect 11173 10310 11225 10362
rect 11237 10310 11289 10362
rect 11301 10310 11353 10362
rect 11365 10310 11417 10362
rect 11429 10310 11481 10362
rect 4344 10251 4396 10260
rect 4344 10217 4353 10251
rect 4353 10217 4387 10251
rect 4387 10217 4396 10251
rect 4344 10208 4396 10217
rect 4988 10208 5040 10260
rect 5724 10208 5776 10260
rect 7564 10208 7616 10260
rect 8668 10208 8720 10260
rect 3148 10072 3200 10124
rect 1492 10004 1544 10056
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 3608 9936 3660 9988
rect 1768 9868 1820 9920
rect 2320 9868 2372 9920
rect 4988 10004 5040 10056
rect 5172 10072 5224 10124
rect 6828 10072 6880 10124
rect 5540 9868 5592 9920
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 8116 10004 8168 10056
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 11520 10208 11572 10260
rect 11888 10208 11940 10260
rect 10048 10004 10100 10056
rect 10140 10004 10192 10056
rect 7104 9868 7156 9920
rect 7380 9868 7432 9920
rect 7656 9868 7708 9920
rect 8576 9868 8628 9920
rect 10232 9868 10284 9920
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11520 9936 11572 9988
rect 3870 9766 3922 9818
rect 3934 9766 3986 9818
rect 3998 9766 4050 9818
rect 4062 9766 4114 9818
rect 4126 9766 4178 9818
rect 6791 9766 6843 9818
rect 6855 9766 6907 9818
rect 6919 9766 6971 9818
rect 6983 9766 7035 9818
rect 7047 9766 7099 9818
rect 9712 9766 9764 9818
rect 9776 9766 9828 9818
rect 9840 9766 9892 9818
rect 9904 9766 9956 9818
rect 9968 9766 10020 9818
rect 12633 9766 12685 9818
rect 12697 9766 12749 9818
rect 12761 9766 12813 9818
rect 12825 9766 12877 9818
rect 12889 9766 12941 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 2228 9528 2280 9580
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3148 9596 3200 9648
rect 5540 9596 5592 9648
rect 10232 9664 10284 9716
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6184 9528 6236 9580
rect 3608 9460 3660 9512
rect 4436 9460 4488 9512
rect 4988 9460 5040 9512
rect 5172 9460 5224 9512
rect 9496 9528 9548 9580
rect 6552 9460 6604 9512
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 10048 9528 10100 9580
rect 5724 9324 5776 9376
rect 10140 9392 10192 9444
rect 11060 9528 11112 9580
rect 11704 9528 11756 9580
rect 10968 9392 11020 9444
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 2410 9222 2462 9274
rect 2474 9222 2526 9274
rect 2538 9222 2590 9274
rect 2602 9222 2654 9274
rect 2666 9222 2718 9274
rect 5331 9222 5383 9274
rect 5395 9222 5447 9274
rect 5459 9222 5511 9274
rect 5523 9222 5575 9274
rect 5587 9222 5639 9274
rect 8252 9222 8304 9274
rect 8316 9222 8368 9274
rect 8380 9222 8432 9274
rect 8444 9222 8496 9274
rect 8508 9222 8560 9274
rect 11173 9222 11225 9274
rect 11237 9222 11289 9274
rect 11301 9222 11353 9274
rect 11365 9222 11417 9274
rect 11429 9222 11481 9274
rect 4436 9163 4488 9172
rect 4436 9129 4445 9163
rect 4445 9129 4479 9163
rect 4479 9129 4488 9163
rect 4436 9120 4488 9129
rect 7564 9120 7616 9172
rect 8576 9120 8628 9172
rect 8668 9120 8720 9172
rect 10968 9120 11020 9172
rect 1308 8916 1360 8968
rect 2044 8916 2096 8968
rect 2228 8916 2280 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 7196 8984 7248 9036
rect 5724 8916 5776 8968
rect 7288 8916 7340 8968
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 7840 8984 7892 9036
rect 5540 8848 5592 8900
rect 7472 8848 7524 8900
rect 8300 8891 8352 8900
rect 8300 8857 8309 8891
rect 8309 8857 8343 8891
rect 8343 8857 8352 8891
rect 8300 8848 8352 8857
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 10048 9052 10100 9104
rect 9128 8916 9180 8968
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 11060 8984 11112 9036
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2688 8780 2740 8832
rect 3332 8780 3384 8832
rect 3608 8780 3660 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 6644 8780 6696 8832
rect 8852 8780 8904 8832
rect 9036 8780 9088 8832
rect 10140 8891 10192 8900
rect 10140 8857 10149 8891
rect 10149 8857 10183 8891
rect 10183 8857 10192 8891
rect 10140 8848 10192 8857
rect 10968 8916 11020 8968
rect 10232 8780 10284 8832
rect 3870 8678 3922 8730
rect 3934 8678 3986 8730
rect 3998 8678 4050 8730
rect 4062 8678 4114 8730
rect 4126 8678 4178 8730
rect 6791 8678 6843 8730
rect 6855 8678 6907 8730
rect 6919 8678 6971 8730
rect 6983 8678 7035 8730
rect 7047 8678 7099 8730
rect 9712 8678 9764 8730
rect 9776 8678 9828 8730
rect 9840 8678 9892 8730
rect 9904 8678 9956 8730
rect 9968 8678 10020 8730
rect 12633 8678 12685 8730
rect 12697 8678 12749 8730
rect 12761 8678 12813 8730
rect 12825 8678 12877 8730
rect 12889 8678 12941 8730
rect 2688 8576 2740 8628
rect 1768 8440 1820 8492
rect 2228 8440 2280 8492
rect 3332 8508 3384 8560
rect 3608 8576 3660 8628
rect 4804 8576 4856 8628
rect 5080 8576 5132 8628
rect 5816 8551 5868 8560
rect 5816 8517 5825 8551
rect 5825 8517 5859 8551
rect 5859 8517 5868 8551
rect 5816 8508 5868 8517
rect 6092 8576 6144 8628
rect 7196 8619 7248 8628
rect 7196 8585 7205 8619
rect 7205 8585 7239 8619
rect 7239 8585 7248 8619
rect 7196 8576 7248 8585
rect 6644 8508 6696 8560
rect 7656 8551 7708 8560
rect 7656 8517 7665 8551
rect 7665 8517 7699 8551
rect 7699 8517 7708 8551
rect 7656 8508 7708 8517
rect 3516 8440 3568 8492
rect 5540 8440 5592 8492
rect 1676 8279 1728 8288
rect 1676 8245 1685 8279
rect 1685 8245 1719 8279
rect 1719 8245 1728 8279
rect 1676 8236 1728 8245
rect 6000 8304 6052 8356
rect 6460 8347 6512 8356
rect 6460 8313 6469 8347
rect 6469 8313 6503 8347
rect 6503 8313 6512 8347
rect 6460 8304 6512 8313
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 9036 8576 9088 8628
rect 9220 8576 9272 8628
rect 9956 8576 10008 8628
rect 10048 8440 10100 8492
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10968 8576 11020 8628
rect 11060 8440 11112 8492
rect 8300 8372 8352 8424
rect 8024 8304 8076 8356
rect 3976 8236 4028 8288
rect 5724 8236 5776 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 2410 8134 2462 8186
rect 2474 8134 2526 8186
rect 2538 8134 2590 8186
rect 2602 8134 2654 8186
rect 2666 8134 2718 8186
rect 5331 8134 5383 8186
rect 5395 8134 5447 8186
rect 5459 8134 5511 8186
rect 5523 8134 5575 8186
rect 5587 8134 5639 8186
rect 8252 8134 8304 8186
rect 8316 8134 8368 8186
rect 8380 8134 8432 8186
rect 8444 8134 8496 8186
rect 8508 8134 8560 8186
rect 11173 8134 11225 8186
rect 11237 8134 11289 8186
rect 11301 8134 11353 8186
rect 11365 8134 11417 8186
rect 11429 8134 11481 8186
rect 1768 8032 1820 8084
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 3240 8032 3292 8084
rect 3976 8075 4028 8084
rect 3976 8041 3985 8075
rect 3985 8041 4019 8075
rect 4019 8041 4028 8075
rect 3976 8032 4028 8041
rect 4252 8032 4304 8084
rect 4804 8032 4856 8084
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 3148 7896 3200 7948
rect 8944 7964 8996 8016
rect 3700 7896 3752 7948
rect 1492 7828 1544 7880
rect 1676 7871 1728 7880
rect 1676 7837 1710 7871
rect 1710 7837 1728 7871
rect 1676 7828 1728 7837
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 5080 7828 5132 7880
rect 5724 7828 5776 7880
rect 6460 7828 6512 7880
rect 7840 7828 7892 7880
rect 8852 7828 8904 7880
rect 9128 7871 9180 7880
rect 9128 7837 9145 7871
rect 9145 7837 9180 7871
rect 9128 7828 9180 7837
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 5448 7760 5500 7812
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10048 7828 10100 7880
rect 3608 7692 3660 7744
rect 6276 7692 6328 7744
rect 6644 7692 6696 7744
rect 8760 7692 8812 7744
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 11060 7692 11112 7744
rect 12440 7735 12492 7744
rect 12440 7701 12449 7735
rect 12449 7701 12483 7735
rect 12483 7701 12492 7735
rect 12440 7692 12492 7701
rect 3870 7590 3922 7642
rect 3934 7590 3986 7642
rect 3998 7590 4050 7642
rect 4062 7590 4114 7642
rect 4126 7590 4178 7642
rect 6791 7590 6843 7642
rect 6855 7590 6907 7642
rect 6919 7590 6971 7642
rect 6983 7590 7035 7642
rect 7047 7590 7099 7642
rect 9712 7590 9764 7642
rect 9776 7590 9828 7642
rect 9840 7590 9892 7642
rect 9904 7590 9956 7642
rect 9968 7590 10020 7642
rect 12633 7590 12685 7642
rect 12697 7590 12749 7642
rect 12761 7590 12813 7642
rect 12825 7590 12877 7642
rect 12889 7590 12941 7642
rect 5448 7488 5500 7540
rect 8576 7488 8628 7540
rect 8760 7531 8812 7540
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 10048 7488 10100 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 2872 7420 2924 7472
rect 3148 7420 3200 7472
rect 2228 7352 2280 7404
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 3700 7352 3752 7404
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 3792 7284 3844 7336
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 6276 7420 6328 7472
rect 8116 7420 8168 7472
rect 6460 7352 6512 7404
rect 8024 7352 8076 7404
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 3516 7148 3568 7200
rect 5540 7216 5592 7268
rect 7748 7284 7800 7336
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9220 7284 9272 7336
rect 9864 7284 9916 7336
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 6552 7148 6604 7200
rect 7472 7148 7524 7200
rect 2410 7046 2462 7098
rect 2474 7046 2526 7098
rect 2538 7046 2590 7098
rect 2602 7046 2654 7098
rect 2666 7046 2718 7098
rect 5331 7046 5383 7098
rect 5395 7046 5447 7098
rect 5459 7046 5511 7098
rect 5523 7046 5575 7098
rect 5587 7046 5639 7098
rect 8252 7046 8304 7098
rect 8316 7046 8368 7098
rect 8380 7046 8432 7098
rect 8444 7046 8496 7098
rect 8508 7046 8560 7098
rect 11173 7046 11225 7098
rect 11237 7046 11289 7098
rect 11301 7046 11353 7098
rect 11365 7046 11417 7098
rect 11429 7046 11481 7098
rect 1768 6944 1820 6996
rect 2320 6944 2372 6996
rect 6460 6944 6512 6996
rect 7472 6944 7524 6996
rect 11060 6944 11112 6996
rect 2688 6876 2740 6928
rect 3148 6876 3200 6928
rect 8944 6876 8996 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 6184 6808 6236 6860
rect 7748 6851 7800 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 5724 6740 5776 6792
rect 6000 6740 6052 6792
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 6644 6740 6696 6792
rect 7380 6740 7432 6792
rect 7840 6740 7892 6792
rect 8576 6740 8628 6792
rect 9128 6783 9180 6792
rect 9128 6749 9145 6783
rect 9145 6749 9180 6783
rect 9128 6740 9180 6749
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 3424 6672 3476 6724
rect 7196 6672 7248 6724
rect 8024 6672 8076 6724
rect 3792 6604 3844 6656
rect 4896 6604 4948 6656
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 6644 6604 6696 6656
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 12072 6808 12124 6860
rect 10232 6740 10284 6792
rect 11060 6740 11112 6792
rect 9956 6604 10008 6656
rect 10324 6604 10376 6656
rect 3870 6502 3922 6554
rect 3934 6502 3986 6554
rect 3998 6502 4050 6554
rect 4062 6502 4114 6554
rect 4126 6502 4178 6554
rect 6791 6502 6843 6554
rect 6855 6502 6907 6554
rect 6919 6502 6971 6554
rect 6983 6502 7035 6554
rect 7047 6502 7099 6554
rect 9712 6502 9764 6554
rect 9776 6502 9828 6554
rect 9840 6502 9892 6554
rect 9904 6502 9956 6554
rect 9968 6502 10020 6554
rect 12633 6502 12685 6554
rect 12697 6502 12749 6554
rect 12761 6502 12813 6554
rect 12825 6502 12877 6554
rect 12889 6502 12941 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 8668 6400 8720 6452
rect 8944 6400 8996 6452
rect 11060 6400 11112 6452
rect 3056 6332 3108 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 3700 6264 3752 6316
rect 2872 6196 2924 6248
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 11612 6264 11664 6316
rect 12072 6264 12124 6316
rect 5816 6128 5868 6180
rect 6276 6128 6328 6180
rect 8576 6196 8628 6248
rect 9128 6196 9180 6248
rect 10324 6196 10376 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 3332 6060 3384 6112
rect 3976 6060 4028 6112
rect 8852 6060 8904 6112
rect 9312 6060 9364 6112
rect 9956 6060 10008 6112
rect 2410 5958 2462 6010
rect 2474 5958 2526 6010
rect 2538 5958 2590 6010
rect 2602 5958 2654 6010
rect 2666 5958 2718 6010
rect 5331 5958 5383 6010
rect 5395 5958 5447 6010
rect 5459 5958 5511 6010
rect 5523 5958 5575 6010
rect 5587 5958 5639 6010
rect 8252 5958 8304 6010
rect 8316 5958 8368 6010
rect 8380 5958 8432 6010
rect 8444 5958 8496 6010
rect 8508 5958 8560 6010
rect 11173 5958 11225 6010
rect 11237 5958 11289 6010
rect 11301 5958 11353 6010
rect 11365 5958 11417 6010
rect 11429 5958 11481 6010
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 5816 5856 5868 5908
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 4436 5763 4488 5772
rect 1400 5652 1452 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 1952 5584 2004 5636
rect 3700 5584 3752 5636
rect 3240 5516 3292 5568
rect 3608 5516 3660 5568
rect 4344 5584 4396 5636
rect 4712 5584 4764 5636
rect 6000 5652 6052 5704
rect 7380 5720 7432 5772
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 4252 5516 4304 5568
rect 5172 5516 5224 5568
rect 7196 5627 7248 5636
rect 7196 5593 7205 5627
rect 7205 5593 7239 5627
rect 7239 5593 7248 5627
rect 7196 5584 7248 5593
rect 8852 5720 8904 5772
rect 9128 5856 9180 5908
rect 9404 5856 9456 5908
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8668 5652 8720 5704
rect 8392 5627 8444 5636
rect 8392 5593 8401 5627
rect 8401 5593 8435 5627
rect 8435 5593 8444 5627
rect 8392 5584 8444 5593
rect 11520 5856 11572 5908
rect 11888 5856 11940 5908
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 9220 5627 9272 5636
rect 9220 5593 9229 5627
rect 9229 5593 9263 5627
rect 9263 5593 9272 5627
rect 9220 5584 9272 5593
rect 9312 5627 9364 5636
rect 9312 5593 9321 5627
rect 9321 5593 9355 5627
rect 9355 5593 9364 5627
rect 9312 5584 9364 5593
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 10324 5652 10376 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 8576 5516 8628 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 10048 5516 10100 5568
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 10968 5516 11020 5568
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12164 5652 12216 5704
rect 11520 5516 11572 5525
rect 3870 5414 3922 5466
rect 3934 5414 3986 5466
rect 3998 5414 4050 5466
rect 4062 5414 4114 5466
rect 4126 5414 4178 5466
rect 6791 5414 6843 5466
rect 6855 5414 6907 5466
rect 6919 5414 6971 5466
rect 6983 5414 7035 5466
rect 7047 5414 7099 5466
rect 9712 5414 9764 5466
rect 9776 5414 9828 5466
rect 9840 5414 9892 5466
rect 9904 5414 9956 5466
rect 9968 5414 10020 5466
rect 12633 5414 12685 5466
rect 12697 5414 12749 5466
rect 12761 5414 12813 5466
rect 12825 5414 12877 5466
rect 12889 5414 12941 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 4436 5312 4488 5364
rect 6000 5312 6052 5364
rect 8300 5312 8352 5364
rect 8484 5312 8536 5364
rect 9772 5312 9824 5364
rect 11520 5312 11572 5364
rect 12164 5312 12216 5364
rect 4252 5244 4304 5296
rect 2320 5176 2372 5228
rect 3516 5176 3568 5228
rect 6184 5244 6236 5296
rect 6644 5244 6696 5296
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 5724 5108 5776 5160
rect 7380 5176 7432 5228
rect 9588 5244 9640 5296
rect 8668 5176 8720 5228
rect 10048 5176 10100 5228
rect 10140 5176 10192 5228
rect 10968 5176 11020 5228
rect 8484 5108 8536 5160
rect 9404 5108 9456 5160
rect 7012 5040 7064 5092
rect 7196 5040 7248 5092
rect 5080 4972 5132 5024
rect 6736 5015 6788 5024
rect 6736 4981 6745 5015
rect 6745 4981 6779 5015
rect 6779 4981 6788 5015
rect 6736 4972 6788 4981
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 8576 4972 8628 5024
rect 10324 4972 10376 5024
rect 10508 4972 10560 5024
rect 2410 4870 2462 4922
rect 2474 4870 2526 4922
rect 2538 4870 2590 4922
rect 2602 4870 2654 4922
rect 2666 4870 2718 4922
rect 5331 4870 5383 4922
rect 5395 4870 5447 4922
rect 5459 4870 5511 4922
rect 5523 4870 5575 4922
rect 5587 4870 5639 4922
rect 8252 4870 8304 4922
rect 8316 4870 8368 4922
rect 8380 4870 8432 4922
rect 8444 4870 8496 4922
rect 8508 4870 8560 4922
rect 11173 4870 11225 4922
rect 11237 4870 11289 4922
rect 11301 4870 11353 4922
rect 11365 4870 11417 4922
rect 11429 4870 11481 4922
rect 3056 4768 3108 4820
rect 3424 4768 3476 4820
rect 4160 4768 4212 4820
rect 4712 4768 4764 4820
rect 5816 4768 5868 4820
rect 3608 4700 3660 4752
rect 5540 4700 5592 4752
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 3700 4632 3752 4684
rect 2228 4496 2280 4548
rect 3148 4496 3200 4548
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3516 4564 3568 4616
rect 3608 4564 3660 4616
rect 3792 4564 3844 4616
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4344 4564 4396 4616
rect 4896 4632 4948 4684
rect 5816 4632 5868 4684
rect 6736 4768 6788 4820
rect 7012 4768 7064 4820
rect 8024 4768 8076 4820
rect 8668 4768 8720 4820
rect 9772 4768 9824 4820
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 5080 4428 5132 4480
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 5632 4428 5684 4480
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 8300 4428 8352 4480
rect 8668 4632 8720 4684
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 10048 4700 10100 4752
rect 10876 4743 10928 4752
rect 10876 4709 10885 4743
rect 10885 4709 10919 4743
rect 10919 4709 10928 4743
rect 10876 4700 10928 4709
rect 12164 4743 12216 4752
rect 12164 4709 12173 4743
rect 12173 4709 12207 4743
rect 12207 4709 12216 4743
rect 12164 4700 12216 4709
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 12072 4632 12124 4684
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9588 4428 9640 4480
rect 9772 4428 9824 4480
rect 11980 4428 12032 4480
rect 3870 4326 3922 4378
rect 3934 4326 3986 4378
rect 3998 4326 4050 4378
rect 4062 4326 4114 4378
rect 4126 4326 4178 4378
rect 6791 4326 6843 4378
rect 6855 4326 6907 4378
rect 6919 4326 6971 4378
rect 6983 4326 7035 4378
rect 7047 4326 7099 4378
rect 9712 4326 9764 4378
rect 9776 4326 9828 4378
rect 9840 4326 9892 4378
rect 9904 4326 9956 4378
rect 9968 4326 10020 4378
rect 12633 4326 12685 4378
rect 12697 4326 12749 4378
rect 12761 4326 12813 4378
rect 12825 4326 12877 4378
rect 12889 4326 12941 4378
rect 2228 4267 2280 4276
rect 2228 4233 2237 4267
rect 2237 4233 2271 4267
rect 2271 4233 2280 4267
rect 2228 4224 2280 4233
rect 3148 4224 3200 4276
rect 3424 4224 3476 4276
rect 3700 4224 3752 4276
rect 5172 4224 5224 4276
rect 5540 4224 5592 4276
rect 5908 4267 5960 4276
rect 5908 4233 5917 4267
rect 5917 4233 5951 4267
rect 5951 4233 5960 4267
rect 5908 4224 5960 4233
rect 9588 4224 9640 4276
rect 10232 4224 10284 4276
rect 12072 4224 12124 4276
rect 2964 4088 3016 4140
rect 3332 4088 3384 4140
rect 3516 4088 3568 4140
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 3516 3952 3568 4004
rect 5632 3952 5684 4004
rect 3700 3884 3752 3936
rect 4988 3884 5040 3936
rect 6000 3884 6052 3936
rect 8300 4088 8352 4140
rect 8668 4088 8720 4140
rect 9404 4088 9456 4140
rect 10048 4088 10100 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 12164 4020 12216 4072
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11980 3884 12032 3936
rect 2410 3782 2462 3834
rect 2474 3782 2526 3834
rect 2538 3782 2590 3834
rect 2602 3782 2654 3834
rect 2666 3782 2718 3834
rect 5331 3782 5383 3834
rect 5395 3782 5447 3834
rect 5459 3782 5511 3834
rect 5523 3782 5575 3834
rect 5587 3782 5639 3834
rect 8252 3782 8304 3834
rect 8316 3782 8368 3834
rect 8380 3782 8432 3834
rect 8444 3782 8496 3834
rect 8508 3782 8560 3834
rect 11173 3782 11225 3834
rect 11237 3782 11289 3834
rect 11301 3782 11353 3834
rect 11365 3782 11417 3834
rect 11429 3782 11481 3834
rect 3516 3680 3568 3732
rect 4896 3680 4948 3732
rect 4988 3680 5040 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 10324 3680 10376 3732
rect 5172 3612 5224 3664
rect 5816 3612 5868 3664
rect 6644 3612 6696 3664
rect 11060 3612 11112 3664
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 4804 3476 4856 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 3700 3408 3752 3460
rect 5356 3451 5408 3460
rect 5356 3417 5365 3451
rect 5365 3417 5399 3451
rect 5399 3417 5408 3451
rect 5356 3408 5408 3417
rect 6184 3544 6236 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 12164 3544 12216 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 10232 3476 10284 3528
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5816 3383 5868 3392
rect 5816 3349 5825 3383
rect 5825 3349 5859 3383
rect 5859 3349 5868 3383
rect 5816 3340 5868 3349
rect 6552 3340 6604 3392
rect 7380 3340 7432 3392
rect 10784 3340 10836 3392
rect 3870 3238 3922 3290
rect 3934 3238 3986 3290
rect 3998 3238 4050 3290
rect 4062 3238 4114 3290
rect 4126 3238 4178 3290
rect 6791 3238 6843 3290
rect 6855 3238 6907 3290
rect 6919 3238 6971 3290
rect 6983 3238 7035 3290
rect 7047 3238 7099 3290
rect 9712 3238 9764 3290
rect 9776 3238 9828 3290
rect 9840 3238 9892 3290
rect 9904 3238 9956 3290
rect 9968 3238 10020 3290
rect 12633 3238 12685 3290
rect 12697 3238 12749 3290
rect 12761 3238 12813 3290
rect 12825 3238 12877 3290
rect 12889 3238 12941 3290
rect 3700 3136 3752 3188
rect 4344 3136 4396 3188
rect 4804 3136 4856 3188
rect 5356 3136 5408 3188
rect 6368 3136 6420 3188
rect 6644 3136 6696 3188
rect 4252 3111 4304 3120
rect 4252 3077 4261 3111
rect 4261 3077 4295 3111
rect 4295 3077 4304 3111
rect 4252 3068 4304 3077
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 3148 3000 3200 3052
rect 2320 2932 2372 2984
rect 2136 2796 2188 2848
rect 2780 2796 2832 2848
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4436 3000 4488 3052
rect 4712 3000 4764 3052
rect 6828 3068 6880 3120
rect 8852 3111 8904 3120
rect 8852 3077 8861 3111
rect 8861 3077 8895 3111
rect 8895 3077 8904 3111
rect 8852 3068 8904 3077
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11704 3136 11756 3188
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7472 3000 7524 3052
rect 11060 3000 11112 3052
rect 11612 3000 11664 3052
rect 6184 2864 6236 2916
rect 4712 2796 4764 2848
rect 6644 2864 6696 2916
rect 7196 2864 7248 2916
rect 11244 2932 11296 2984
rect 11796 2932 11848 2984
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 9496 2839 9548 2848
rect 9496 2805 9505 2839
rect 9505 2805 9539 2839
rect 9539 2805 9548 2839
rect 9496 2796 9548 2805
rect 2410 2694 2462 2746
rect 2474 2694 2526 2746
rect 2538 2694 2590 2746
rect 2602 2694 2654 2746
rect 2666 2694 2718 2746
rect 5331 2694 5383 2746
rect 5395 2694 5447 2746
rect 5459 2694 5511 2746
rect 5523 2694 5575 2746
rect 5587 2694 5639 2746
rect 8252 2694 8304 2746
rect 8316 2694 8368 2746
rect 8380 2694 8432 2746
rect 8444 2694 8496 2746
rect 8508 2694 8560 2746
rect 11173 2694 11225 2746
rect 11237 2694 11289 2746
rect 11301 2694 11353 2746
rect 11365 2694 11417 2746
rect 11429 2694 11481 2746
rect 2872 2592 2924 2644
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 11612 2524 11664 2576
rect 4344 2456 4396 2508
rect 4436 2456 4488 2508
rect 756 2388 808 2440
rect 2136 2388 2188 2440
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 3792 2388 3844 2440
rect 5816 2456 5868 2508
rect 11796 2456 11848 2508
rect 2412 2320 2464 2372
rect 4712 2363 4764 2372
rect 4712 2329 4721 2363
rect 4721 2329 4755 2363
rect 4755 2329 4764 2363
rect 7288 2388 7340 2440
rect 8576 2388 8628 2440
rect 9496 2388 9548 2440
rect 11704 2388 11756 2440
rect 4712 2320 4764 2329
rect 1676 2295 1728 2304
rect 1676 2261 1685 2295
rect 1685 2261 1719 2295
rect 1719 2261 1728 2295
rect 1676 2252 1728 2261
rect 4436 2252 4488 2304
rect 4620 2252 4672 2304
rect 4804 2252 4856 2304
rect 3870 2150 3922 2202
rect 3934 2150 3986 2202
rect 3998 2150 4050 2202
rect 4062 2150 4114 2202
rect 4126 2150 4178 2202
rect 6791 2150 6843 2202
rect 6855 2150 6907 2202
rect 6919 2150 6971 2202
rect 6983 2150 7035 2202
rect 7047 2150 7099 2202
rect 9712 2150 9764 2202
rect 9776 2150 9828 2202
rect 9840 2150 9892 2202
rect 9904 2150 9956 2202
rect 9968 2150 10020 2202
rect 12633 2150 12685 2202
rect 12697 2150 12749 2202
rect 12761 2150 12813 2202
rect 12825 2150 12877 2202
rect 12889 2150 12941 2202
rect 2044 2048 2096 2100
rect 2872 2048 2924 2100
rect 1400 1776 1452 1828
rect 2412 1912 2464 1964
rect 3148 1912 3200 1964
rect 4252 2048 4304 2100
rect 4712 2048 4764 2100
rect 4896 2048 4948 2100
rect 6184 2091 6236 2100
rect 6184 2057 6193 2091
rect 6193 2057 6227 2091
rect 6227 2057 6236 2091
rect 6184 2048 6236 2057
rect 4436 1912 4488 1964
rect 4712 1912 4764 1964
rect 6000 1980 6052 2032
rect 8668 2091 8720 2100
rect 8668 2057 8677 2091
rect 8677 2057 8711 2091
rect 8711 2057 8720 2091
rect 8668 2048 8720 2057
rect 6644 1912 6696 1964
rect 7012 1955 7064 1964
rect 7012 1921 7021 1955
rect 7021 1921 7055 1955
rect 7055 1921 7064 1955
rect 7012 1912 7064 1921
rect 2228 1708 2280 1760
rect 3884 1708 3936 1760
rect 4712 1751 4764 1760
rect 4712 1717 4721 1751
rect 4721 1717 4755 1751
rect 4755 1717 4764 1751
rect 4712 1708 4764 1717
rect 4988 1708 5040 1760
rect 5172 1708 5224 1760
rect 6920 1819 6972 1828
rect 6920 1785 6929 1819
rect 6929 1785 6963 1819
rect 6963 1785 6972 1819
rect 6920 1776 6972 1785
rect 2410 1606 2462 1658
rect 2474 1606 2526 1658
rect 2538 1606 2590 1658
rect 2602 1606 2654 1658
rect 2666 1606 2718 1658
rect 5331 1606 5383 1658
rect 5395 1606 5447 1658
rect 5459 1606 5511 1658
rect 5523 1606 5575 1658
rect 5587 1606 5639 1658
rect 8252 1606 8304 1658
rect 8316 1606 8368 1658
rect 8380 1606 8432 1658
rect 8444 1606 8496 1658
rect 8508 1606 8560 1658
rect 11173 1606 11225 1658
rect 11237 1606 11289 1658
rect 11301 1606 11353 1658
rect 11365 1606 11417 1658
rect 11429 1606 11481 1658
rect 2044 1504 2096 1556
rect 1400 1411 1452 1420
rect 1400 1377 1409 1411
rect 1409 1377 1443 1411
rect 1443 1377 1452 1411
rect 1400 1368 1452 1377
rect 2780 1547 2832 1556
rect 2780 1513 2789 1547
rect 2789 1513 2823 1547
rect 2823 1513 2832 1547
rect 2780 1504 2832 1513
rect 3148 1547 3200 1556
rect 3148 1513 3157 1547
rect 3157 1513 3191 1547
rect 3191 1513 3200 1547
rect 3148 1504 3200 1513
rect 4896 1504 4948 1556
rect 7012 1504 7064 1556
rect 1676 1343 1728 1352
rect 1676 1309 1710 1343
rect 1710 1309 1728 1343
rect 1676 1300 1728 1309
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 3884 1368 3936 1420
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4712 1300 4764 1352
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4804 1300 4856 1309
rect 4988 1232 5040 1284
rect 6920 1300 6972 1352
rect 5172 1164 5224 1216
rect 3870 1062 3922 1114
rect 3934 1062 3986 1114
rect 3998 1062 4050 1114
rect 4062 1062 4114 1114
rect 4126 1062 4178 1114
rect 6791 1062 6843 1114
rect 6855 1062 6907 1114
rect 6919 1062 6971 1114
rect 6983 1062 7035 1114
rect 7047 1062 7099 1114
rect 9712 1062 9764 1114
rect 9776 1062 9828 1114
rect 9840 1062 9892 1114
rect 9904 1062 9956 1114
rect 9968 1062 10020 1114
rect 12633 1062 12685 1114
rect 12697 1062 12749 1114
rect 12761 1062 12813 1114
rect 12825 1062 12877 1114
rect 12889 1062 12941 1114
<< metal2 >>
rect 4342 12880 4398 12889
rect 4342 12815 4398 12824
rect 2410 12540 2718 12549
rect 2410 12538 2416 12540
rect 2472 12538 2496 12540
rect 2552 12538 2576 12540
rect 2632 12538 2656 12540
rect 2712 12538 2718 12540
rect 2472 12486 2474 12538
rect 2654 12486 2656 12538
rect 2410 12484 2416 12486
rect 2472 12484 2496 12486
rect 2552 12484 2576 12486
rect 2632 12484 2656 12486
rect 2712 12484 2718 12486
rect 2410 12475 2718 12484
rect 4356 12442 4384 12815
rect 5331 12540 5639 12549
rect 5331 12538 5337 12540
rect 5393 12538 5417 12540
rect 5473 12538 5497 12540
rect 5553 12538 5577 12540
rect 5633 12538 5639 12540
rect 5393 12486 5395 12538
rect 5575 12486 5577 12538
rect 5331 12484 5337 12486
rect 5393 12484 5417 12486
rect 5473 12484 5497 12486
rect 5553 12484 5577 12486
rect 5633 12484 5639 12486
rect 5331 12475 5639 12484
rect 8252 12540 8560 12549
rect 8252 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8498 12540
rect 8554 12538 8560 12540
rect 8314 12486 8316 12538
rect 8496 12486 8498 12538
rect 8252 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8498 12486
rect 8554 12484 8560 12486
rect 8252 12475 8560 12484
rect 11173 12540 11481 12549
rect 11173 12538 11179 12540
rect 11235 12538 11259 12540
rect 11315 12538 11339 12540
rect 11395 12538 11419 12540
rect 11475 12538 11481 12540
rect 11235 12486 11237 12538
rect 11417 12486 11419 12538
rect 11173 12484 11179 12486
rect 11235 12484 11259 12486
rect 11315 12484 11339 12486
rect 11395 12484 11419 12486
rect 11475 12484 11481 12486
rect 11173 12475 11481 12484
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 1308 12164 1360 12170
rect 1308 12106 1360 12112
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 1320 12073 1348 12106
rect 1306 12064 1362 12073
rect 1306 11999 1362 12008
rect 3528 11898 3556 12106
rect 3870 11996 4178 12005
rect 3870 11994 3876 11996
rect 3932 11994 3956 11996
rect 4012 11994 4036 11996
rect 4092 11994 4116 11996
rect 4172 11994 4178 11996
rect 3932 11942 3934 11994
rect 4114 11942 4116 11994
rect 3870 11940 3876 11942
rect 3932 11940 3956 11942
rect 4012 11940 4036 11942
rect 4092 11940 4116 11942
rect 4172 11940 4178 11942
rect 3870 11931 4178 11940
rect 5552 11898 5580 12106
rect 5644 11898 5672 12174
rect 5828 11898 5856 12242
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 1320 11257 1348 11494
rect 2410 11452 2718 11461
rect 2410 11450 2416 11452
rect 2472 11450 2496 11452
rect 2552 11450 2576 11452
rect 2632 11450 2656 11452
rect 2712 11450 2718 11452
rect 2472 11398 2474 11450
rect 2654 11398 2656 11450
rect 2410 11396 2416 11398
rect 2472 11396 2496 11398
rect 2552 11396 2576 11398
rect 2632 11396 2656 11398
rect 2712 11396 2718 11398
rect 2410 11387 2718 11396
rect 1306 11248 1362 11257
rect 1306 11183 1362 11192
rect 1320 11150 1348 11183
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1504 10062 1532 11086
rect 1688 10810 1716 11086
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2240 10674 2268 10746
rect 2332 10674 2360 10950
rect 2608 10810 2636 11018
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 1780 10441 1808 10610
rect 1766 10432 1822 10441
rect 1766 10367 1822 10376
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1320 8809 1348 8910
rect 1504 8838 1532 9998
rect 1688 9722 1716 9998
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1780 9625 1808 9862
rect 1766 9616 1822 9625
rect 2240 9586 2268 10610
rect 2410 10364 2718 10373
rect 2410 10362 2416 10364
rect 2472 10362 2496 10364
rect 2552 10362 2576 10364
rect 2632 10362 2656 10364
rect 2712 10362 2718 10364
rect 2472 10310 2474 10362
rect 2654 10310 2656 10362
rect 2410 10308 2416 10310
rect 2472 10308 2496 10310
rect 2552 10308 2576 10310
rect 2632 10308 2656 10310
rect 2712 10308 2718 10310
rect 2410 10299 2718 10308
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2332 9586 2360 9862
rect 1766 9551 1822 9560
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2240 8974 2268 9522
rect 2410 9276 2718 9285
rect 2410 9274 2416 9276
rect 2472 9274 2496 9276
rect 2552 9274 2576 9276
rect 2632 9274 2656 9276
rect 2712 9274 2718 9276
rect 2472 9222 2474 9274
rect 2654 9222 2656 9274
rect 2410 9220 2416 9222
rect 2472 9220 2496 9222
rect 2552 9220 2576 9222
rect 2632 9220 2656 9222
rect 2712 9220 2718 9222
rect 2410 9211 2718 9220
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 1492 8832 1544 8838
rect 1306 8800 1362 8809
rect 1492 8774 1544 8780
rect 1306 8735 1362 8744
rect 1504 7886 1532 8774
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1676 8288 1728 8294
rect 1676 8230 1728 8236
rect 1688 7886 1716 8230
rect 1780 8090 1808 8434
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1780 7993 1808 8026
rect 1766 7984 1822 7993
rect 1766 7919 1822 7928
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2056 7313 2084 8910
rect 2240 8498 2268 8910
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8634 2728 8774
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2240 7410 2268 8434
rect 2410 8188 2718 8197
rect 2410 8186 2416 8188
rect 2472 8186 2496 8188
rect 2552 8186 2576 8188
rect 2632 8186 2656 8188
rect 2712 8186 2718 8188
rect 2472 8134 2474 8186
rect 2654 8134 2656 8186
rect 2410 8132 2416 8134
rect 2472 8132 2496 8134
rect 2552 8132 2576 8134
rect 2632 8132 2656 8134
rect 2712 8132 2718 8134
rect 2410 8123 2718 8132
rect 2872 7472 2924 7478
rect 2792 7420 2872 7426
rect 2792 7414 2924 7420
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2792 7398 2912 7414
rect 2042 7304 2098 7313
rect 2042 7239 2098 7248
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1766 7168 1822 7177
rect 1688 6866 1716 7142
rect 1766 7103 1822 7112
rect 1780 7002 1808 7103
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5710 1440 6734
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 4622 1440 5646
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1964 5370 1992 5578
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 756 2440 808 2446
rect 756 2382 808 2388
rect 768 1465 796 2382
rect 1412 1834 1440 4558
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1400 1828 1452 1834
rect 1400 1770 1452 1776
rect 754 1456 810 1465
rect 1412 1426 1440 1770
rect 754 1391 810 1400
rect 1400 1420 1452 1426
rect 1400 1362 1452 1368
rect 1688 1358 1716 2246
rect 2056 2106 2084 7239
rect 2332 7002 2360 7346
rect 2410 7100 2718 7109
rect 2410 7098 2416 7100
rect 2472 7098 2496 7100
rect 2552 7098 2576 7100
rect 2632 7098 2656 7100
rect 2712 7098 2718 7100
rect 2472 7046 2474 7098
rect 2654 7046 2656 7098
rect 2410 7044 2416 7046
rect 2472 7044 2496 7046
rect 2552 7044 2576 7046
rect 2632 7044 2656 7046
rect 2712 7044 2718 7046
rect 2410 7035 2718 7044
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2688 6928 2740 6934
rect 2792 6914 2820 7398
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2740 6886 2820 6914
rect 2688 6870 2740 6876
rect 2884 6254 2912 7278
rect 2976 6458 3004 10678
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3160 10130 3188 10610
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3160 9654 3188 10066
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8090 3096 8910
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3160 7954 3188 9590
rect 3252 9586 3280 10610
rect 3528 10470 3556 11494
rect 3804 11354 3832 11698
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 4356 11150 4384 11630
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4448 11354 4476 11562
rect 6104 11558 6132 12106
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6472 11694 6500 12174
rect 6791 11996 7099 12005
rect 6791 11994 6797 11996
rect 6853 11994 6877 11996
rect 6933 11994 6957 11996
rect 7013 11994 7037 11996
rect 7093 11994 7099 11996
rect 6853 11942 6855 11994
rect 7035 11942 7037 11994
rect 6791 11940 6797 11942
rect 6853 11940 6877 11942
rect 6933 11940 6957 11942
rect 7013 11940 7037 11942
rect 7093 11940 7099 11942
rect 6791 11931 7099 11940
rect 8404 11898 8432 12174
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8956 11762 8984 12038
rect 9712 11996 10020 12005
rect 9712 11994 9718 11996
rect 9774 11994 9798 11996
rect 9854 11994 9878 11996
rect 9934 11994 9958 11996
rect 10014 11994 10020 11996
rect 9774 11942 9776 11994
rect 9956 11942 9958 11994
rect 9712 11940 9718 11942
rect 9774 11940 9798 11942
rect 9854 11940 9878 11942
rect 9934 11940 9958 11942
rect 10014 11940 10020 11942
rect 9712 11931 10020 11940
rect 10060 11898 10088 12174
rect 10336 11898 10364 12174
rect 10612 11898 10640 12174
rect 10888 11898 10916 12174
rect 11164 11898 11192 12174
rect 12633 11996 12941 12005
rect 12633 11994 12639 11996
rect 12695 11994 12719 11996
rect 12775 11994 12799 11996
rect 12855 11994 12879 11996
rect 12935 11994 12941 11996
rect 12695 11942 12697 11994
rect 12877 11942 12879 11994
rect 12633 11940 12639 11942
rect 12695 11940 12719 11942
rect 12775 11940 12799 11942
rect 12855 11940 12879 11942
rect 12935 11940 12941 11942
rect 12633 11931 12941 11940
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5331 11452 5639 11461
rect 5331 11450 5337 11452
rect 5393 11450 5417 11452
rect 5473 11450 5497 11452
rect 5553 11450 5577 11452
rect 5633 11450 5639 11452
rect 5393 11398 5395 11450
rect 5575 11398 5577 11450
rect 5331 11396 5337 11398
rect 5393 11396 5417 11398
rect 5473 11396 5497 11398
rect 5553 11396 5577 11398
rect 5633 11396 5639 11398
rect 5331 11387 5639 11396
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 8090 3280 9522
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8566 3372 8774
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3528 8498 3556 10406
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3620 9518 3648 9930
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8634 3648 8774
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3160 7478 3188 7890
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3160 7342 3188 7414
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3068 6390 3096 7278
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2410 6012 2718 6021
rect 2410 6010 2416 6012
rect 2472 6010 2496 6012
rect 2552 6010 2576 6012
rect 2632 6010 2656 6012
rect 2712 6010 2718 6012
rect 2472 5958 2474 6010
rect 2654 5958 2656 6010
rect 2410 5956 2416 5958
rect 2472 5956 2496 5958
rect 2552 5956 2576 5958
rect 2632 5956 2656 5958
rect 2712 5956 2718 5958
rect 2410 5947 2718 5956
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2240 4282 2268 4490
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2332 4162 2360 5170
rect 2410 4924 2718 4933
rect 2410 4922 2416 4924
rect 2472 4922 2496 4924
rect 2552 4922 2576 4924
rect 2632 4922 2656 4924
rect 2712 4922 2718 4924
rect 2472 4870 2474 4922
rect 2654 4870 2656 4922
rect 2410 4868 2416 4870
rect 2472 4868 2496 4870
rect 2552 4868 2576 4870
rect 2632 4868 2656 4870
rect 2712 4868 2718 4870
rect 2410 4859 2718 4868
rect 2240 4134 2360 4162
rect 2240 3058 2268 4134
rect 2410 3836 2718 3845
rect 2410 3834 2416 3836
rect 2472 3834 2496 3836
rect 2552 3834 2576 3836
rect 2632 3834 2656 3836
rect 2712 3834 2718 3836
rect 2472 3782 2474 3834
rect 2654 3782 2656 3834
rect 2410 3780 2416 3782
rect 2472 3780 2496 3782
rect 2552 3780 2576 3782
rect 2632 3780 2656 3782
rect 2712 3780 2718 3782
rect 2410 3771 2718 3780
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2446 2176 2790
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2056 1562 2084 2042
rect 2240 1766 2268 2994
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 2530 2360 2926
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2410 2748 2718 2757
rect 2410 2746 2416 2748
rect 2472 2746 2496 2748
rect 2552 2746 2576 2748
rect 2632 2746 2656 2748
rect 2712 2746 2718 2748
rect 2472 2694 2474 2746
rect 2654 2694 2656 2746
rect 2410 2692 2416 2694
rect 2472 2692 2496 2694
rect 2552 2692 2576 2694
rect 2632 2692 2656 2694
rect 2712 2692 2718 2694
rect 2410 2683 2718 2692
rect 2332 2502 2452 2530
rect 2424 2378 2452 2502
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2424 1970 2452 2314
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2228 1760 2280 1766
rect 2228 1702 2280 1708
rect 2410 1660 2718 1669
rect 2410 1658 2416 1660
rect 2472 1658 2496 1660
rect 2552 1658 2576 1660
rect 2632 1658 2656 1660
rect 2712 1658 2718 1660
rect 2472 1606 2474 1658
rect 2654 1606 2656 1658
rect 2410 1604 2416 1606
rect 2472 1604 2496 1606
rect 2552 1604 2576 1606
rect 2632 1604 2656 1606
rect 2712 1604 2718 1606
rect 2410 1595 2718 1604
rect 2792 1562 2820 2790
rect 2884 2650 2912 6190
rect 3068 4826 3096 6326
rect 3160 6322 3188 6870
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 4978 3188 5646
rect 3252 5574 3280 6190
rect 3344 6118 3372 7822
rect 3528 7206 3556 7822
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3436 5914 3464 6666
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5148 3280 5510
rect 3528 5234 3556 7142
rect 3620 5574 3648 7686
rect 3712 7410 3740 7890
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3712 6322 3740 7346
rect 3804 7342 3832 11086
rect 3870 10908 4178 10917
rect 3870 10906 3876 10908
rect 3932 10906 3956 10908
rect 4012 10906 4036 10908
rect 4092 10906 4116 10908
rect 4172 10906 4178 10908
rect 3932 10854 3934 10906
rect 4114 10854 4116 10906
rect 3870 10852 3876 10854
rect 3932 10852 3956 10854
rect 4012 10852 4036 10854
rect 4092 10852 4116 10854
rect 4172 10852 4178 10854
rect 3870 10843 4178 10852
rect 4356 10792 4384 11086
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4264 10764 4384 10792
rect 3870 9820 4178 9829
rect 3870 9818 3876 9820
rect 3932 9818 3956 9820
rect 4012 9818 4036 9820
rect 4092 9818 4116 9820
rect 4172 9818 4178 9820
rect 3932 9766 3934 9818
rect 4114 9766 4116 9818
rect 3870 9764 3876 9766
rect 3932 9764 3956 9766
rect 4012 9764 4036 9766
rect 4092 9764 4116 9766
rect 4172 9764 4178 9766
rect 3870 9755 4178 9764
rect 4264 8974 4292 10764
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4356 10266 4384 10610
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4540 10062 4568 10950
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4632 10062 4660 10406
rect 5000 10266 5028 10406
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5184 10130 5212 11018
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5331 10364 5639 10373
rect 5331 10362 5337 10364
rect 5393 10362 5417 10364
rect 5473 10362 5497 10364
rect 5553 10362 5577 10364
rect 5633 10362 5639 10364
rect 5393 10310 5395 10362
rect 5575 10310 5577 10362
rect 5331 10308 5337 10310
rect 5393 10308 5417 10310
rect 5473 10308 5497 10310
rect 5553 10308 5577 10310
rect 5633 10308 5639 10310
rect 5331 10299 5639 10308
rect 5736 10266 5764 10610
rect 5828 10606 5856 11086
rect 6104 10742 6132 11494
rect 6748 11354 6776 11698
rect 8864 11558 8892 11698
rect 8956 11626 8984 11698
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 8252 11452 8560 11461
rect 8252 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8498 11452
rect 8554 11450 8560 11452
rect 8314 11398 8316 11450
rect 8496 11398 8498 11450
rect 8252 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8498 11398
rect 8554 11396 8560 11398
rect 8252 11387 8560 11396
rect 11173 11452 11481 11461
rect 11173 11450 11179 11452
rect 11235 11450 11259 11452
rect 11315 11450 11339 11452
rect 11395 11450 11419 11452
rect 11475 11450 11481 11452
rect 11235 11398 11237 11450
rect 11417 11398 11419 11450
rect 11173 11396 11179 11398
rect 11235 11396 11259 11398
rect 11315 11396 11339 11398
rect 11395 11396 11419 11398
rect 11475 11396 11481 11398
rect 11173 11387 11481 11396
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9518 5028 9998
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9654 5580 9862
rect 5736 9674 5764 10202
rect 5540 9648 5592 9654
rect 5736 9646 5856 9674
rect 5540 9590 5592 9596
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4448 9178 4476 9454
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 3870 8732 4178 8741
rect 3870 8730 3876 8732
rect 3932 8730 3956 8732
rect 4012 8730 4036 8732
rect 4092 8730 4116 8732
rect 4172 8730 4178 8732
rect 3932 8678 3934 8730
rect 4114 8678 4116 8730
rect 3870 8676 3876 8678
rect 3932 8676 3956 8678
rect 4012 8676 4036 8678
rect 4092 8676 4116 8678
rect 4172 8676 4178 8678
rect 3870 8667 4178 8676
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 8090 4016 8230
rect 4264 8090 4292 8910
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4448 7886 4476 9114
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8634 4844 8774
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 3870 7644 4178 7653
rect 3870 7642 3876 7644
rect 3932 7642 3956 7644
rect 4012 7642 4036 7644
rect 4092 7642 4116 7644
rect 4172 7642 4178 7644
rect 3932 7590 3934 7642
rect 4114 7590 4116 7642
rect 3870 7588 3876 7590
rect 3932 7588 3956 7590
rect 4012 7588 4036 7590
rect 4092 7588 4116 7590
rect 4172 7588 4178 7590
rect 3870 7579 4178 7588
rect 4448 7342 4476 7822
rect 4816 7410 4844 8026
rect 5092 7886 5120 8570
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5092 7410 5120 7822
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 5184 6662 5212 9454
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5331 9276 5639 9285
rect 5331 9274 5337 9276
rect 5393 9274 5417 9276
rect 5473 9274 5497 9276
rect 5553 9274 5577 9276
rect 5633 9274 5639 9276
rect 5393 9222 5395 9274
rect 5575 9222 5577 9274
rect 5331 9220 5337 9222
rect 5393 9220 5417 9222
rect 5473 9220 5497 9222
rect 5553 9220 5577 9222
rect 5633 9220 5639 9222
rect 5331 9211 5639 9220
rect 5736 8974 5764 9318
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8498 5580 8842
rect 5828 8566 5856 9646
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5331 8188 5639 8197
rect 5331 8186 5337 8188
rect 5393 8186 5417 8188
rect 5473 8186 5497 8188
rect 5553 8186 5577 8188
rect 5633 8186 5639 8188
rect 5393 8134 5395 8186
rect 5575 8134 5577 8186
rect 5331 8132 5337 8134
rect 5393 8132 5417 8134
rect 5473 8132 5497 8134
rect 5553 8132 5577 8134
rect 5633 8132 5639 8134
rect 5331 8123 5639 8132
rect 5736 7886 5764 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5460 7546 5488 7754
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5538 7304 5594 7313
rect 5538 7239 5540 7248
rect 5592 7239 5594 7248
rect 5540 7210 5592 7216
rect 5331 7100 5639 7109
rect 5331 7098 5337 7100
rect 5393 7098 5417 7100
rect 5473 7098 5497 7100
rect 5553 7098 5577 7100
rect 5633 7098 5639 7100
rect 5393 7046 5395 7098
rect 5575 7046 5577 7098
rect 5331 7044 5337 7046
rect 5393 7044 5417 7046
rect 5473 7044 5497 7046
rect 5553 7044 5577 7046
rect 5633 7044 5639 7046
rect 5331 7035 5639 7044
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3804 5794 3832 6598
rect 3870 6556 4178 6565
rect 3870 6554 3876 6556
rect 3932 6554 3956 6556
rect 4012 6554 4036 6556
rect 4092 6554 4116 6556
rect 4172 6554 4178 6556
rect 3932 6502 3934 6554
rect 4114 6502 4116 6554
rect 3870 6500 3876 6502
rect 3932 6500 3956 6502
rect 4012 6500 4036 6502
rect 4092 6500 4116 6502
rect 4172 6500 4178 6502
rect 3870 6491 4178 6500
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3712 5766 3832 5794
rect 3712 5642 3740 5766
rect 3988 5658 4016 6054
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3804 5630 4016 5658
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3252 5120 3372 5148
rect 3160 4950 3280 4978
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3252 4570 3280 4950
rect 3344 4690 3372 5120
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 4622 3464 4762
rect 3620 4758 3648 5510
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3424 4616 3476 4622
rect 3148 4548 3200 4554
rect 3252 4542 3372 4570
rect 3424 4558 3476 4564
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3148 4490 3200 4496
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 4146 3004 4422
rect 3160 4282 3188 4490
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3344 4146 3372 4542
rect 3436 4282 3464 4558
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3528 4146 3556 4558
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3160 2650 3188 2994
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 2884 2106 2912 2586
rect 3344 2446 3372 4082
rect 3620 4078 3648 4558
rect 3712 4282 3740 4626
rect 3804 4622 3832 5630
rect 3988 5574 4016 5630
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3870 5468 4178 5477
rect 3870 5466 3876 5468
rect 3932 5466 3956 5468
rect 4012 5466 4036 5468
rect 4092 5466 4116 5468
rect 4172 5466 4178 5468
rect 3932 5414 3934 5466
rect 4114 5414 4116 5466
rect 3870 5412 3876 5414
rect 3932 5412 3956 5414
rect 4012 5412 4036 5414
rect 4092 5412 4116 5414
rect 4172 5412 4178 5414
rect 3870 5403 4178 5412
rect 4264 5302 4292 5510
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4356 4842 4384 5578
rect 4448 5370 4476 5714
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4264 4814 4384 4842
rect 4172 4622 4200 4762
rect 4264 4622 4292 4814
rect 4448 4706 4476 5306
rect 4724 4826 4752 5578
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4356 4678 4476 4706
rect 4356 4622 4384 4678
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3698 4176 3754 4185
rect 3698 4111 3700 4120
rect 3752 4111 3754 4120
rect 3700 4082 3752 4088
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3528 3738 3556 3946
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3712 3466 3740 3878
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3712 3194 3740 3402
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3804 2446 3832 4422
rect 3870 4380 4178 4389
rect 3870 4378 3876 4380
rect 3932 4378 3956 4380
rect 4012 4378 4036 4380
rect 4092 4378 4116 4380
rect 4172 4378 4178 4380
rect 3932 4326 3934 4378
rect 4114 4326 4116 4378
rect 3870 4324 3876 4326
rect 3932 4324 3956 4326
rect 4012 4324 4036 4326
rect 4092 4324 4116 4326
rect 4172 4324 4178 4326
rect 3870 4315 4178 4324
rect 3870 3292 4178 3301
rect 3870 3290 3876 3292
rect 3932 3290 3956 3292
rect 4012 3290 4036 3292
rect 4092 3290 4116 3292
rect 4172 3290 4178 3292
rect 3932 3238 3934 3290
rect 4114 3238 4116 3290
rect 3870 3236 3876 3238
rect 3932 3236 3956 3238
rect 4012 3236 4036 3238
rect 4092 3236 4116 3238
rect 4172 3236 4178 3238
rect 3870 3227 4178 3236
rect 4264 3210 4292 4558
rect 4264 3188 4476 3210
rect 4264 3182 4344 3188
rect 4396 3182 4476 3188
rect 4344 3130 4396 3136
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 3160 1562 3188 1906
rect 2044 1556 2096 1562
rect 2044 1498 2096 1504
rect 2780 1556 2832 1562
rect 2780 1498 2832 1504
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3344 1358 3372 2382
rect 3870 2204 4178 2213
rect 3870 2202 3876 2204
rect 3932 2202 3956 2204
rect 4012 2202 4036 2204
rect 4092 2202 4116 2204
rect 4172 2202 4178 2204
rect 3932 2150 3934 2202
rect 4114 2150 4116 2202
rect 3870 2148 3876 2150
rect 3932 2148 3956 2150
rect 4012 2148 4036 2150
rect 4092 2148 4116 2150
rect 4172 2148 4178 2150
rect 3870 2139 4178 2148
rect 4264 2106 4292 3062
rect 4448 3058 4476 3182
rect 4724 3058 4752 4762
rect 4908 4690 4936 6598
rect 5736 6066 5764 6734
rect 5920 6458 5948 10610
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6012 8362 6040 9522
rect 6104 8634 6132 9522
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6798 6040 7142
rect 6196 6866 6224 9522
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7478 6316 7686
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5828 6186 5856 6258
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5736 6038 5856 6066
rect 5331 6012 5639 6021
rect 5331 6010 5337 6012
rect 5393 6010 5417 6012
rect 5473 6010 5497 6012
rect 5553 6010 5577 6012
rect 5633 6010 5639 6012
rect 5393 5958 5395 6010
rect 5575 5958 5577 6010
rect 5331 5956 5337 5958
rect 5393 5956 5417 5958
rect 5473 5956 5497 5958
rect 5553 5956 5577 5958
rect 5633 5956 5639 5958
rect 5331 5947 5639 5956
rect 5828 5914 5856 6038
rect 5920 5914 5948 6394
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 3534 4844 4422
rect 4908 3738 4936 4626
rect 5092 4486 5120 4966
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 5092 3738 5120 4422
rect 5184 4282 5212 5510
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5331 4924 5639 4933
rect 5331 4922 5337 4924
rect 5393 4922 5417 4924
rect 5473 4922 5497 4924
rect 5553 4922 5577 4924
rect 5633 4922 5639 4924
rect 5393 4870 5395 4922
rect 5575 4870 5577 4922
rect 5331 4868 5337 4870
rect 5393 4868 5417 4870
rect 5473 4868 5497 4870
rect 5553 4868 5577 4870
rect 5633 4868 5639 4870
rect 5331 4859 5639 4868
rect 5540 4752 5592 4758
rect 5736 4706 5764 5102
rect 5828 4826 5856 5850
rect 6012 5710 6040 6258
rect 6288 6186 6316 7414
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6380 5914 6408 10746
rect 6564 9518 6592 11086
rect 6791 10908 7099 10917
rect 6791 10906 6797 10908
rect 6853 10906 6877 10908
rect 6933 10906 6957 10908
rect 7013 10906 7037 10908
rect 7093 10906 7099 10908
rect 6853 10854 6855 10906
rect 7035 10854 7037 10906
rect 6791 10852 6797 10854
rect 6853 10852 6877 10854
rect 6933 10852 6957 10854
rect 7013 10852 7037 10854
rect 7093 10852 7099 10854
rect 6791 10843 7099 10852
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6932 10146 6960 10678
rect 6840 10130 6960 10146
rect 6828 10124 6960 10130
rect 6880 10118 6960 10124
rect 6828 10066 6880 10072
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9926 7144 9998
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6791 9820 7099 9829
rect 6791 9818 6797 9820
rect 6853 9818 6877 9820
rect 6933 9818 6957 9820
rect 7013 9818 7037 9820
rect 7093 9818 7099 9820
rect 6853 9766 6855 9818
rect 7035 9766 7037 9818
rect 6791 9764 6797 9766
rect 6853 9764 6877 9766
rect 6933 9764 6957 9766
rect 7013 9764 7037 9766
rect 7093 9764 7099 9766
rect 6791 9755 7099 9764
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 7208 9042 7236 11086
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10606 7328 10950
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8566 6684 8774
rect 6791 8732 7099 8741
rect 6791 8730 6797 8732
rect 6853 8730 6877 8732
rect 6933 8730 6957 8732
rect 7013 8730 7037 8732
rect 7093 8730 7099 8732
rect 6853 8678 6855 8730
rect 7035 8678 7037 8730
rect 6791 8676 6797 8678
rect 6853 8676 6877 8678
rect 6933 8676 6957 8678
rect 7013 8676 7037 8678
rect 7093 8676 7099 8678
rect 6791 8667 7099 8676
rect 7208 8634 7236 8978
rect 7300 8974 7328 10542
rect 7392 9926 7420 11086
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9712 10908 10020 10917
rect 9712 10906 9718 10908
rect 9774 10906 9798 10908
rect 9854 10906 9878 10908
rect 9934 10906 9958 10908
rect 10014 10906 10020 10908
rect 9774 10854 9776 10906
rect 9956 10854 9958 10906
rect 9712 10852 9718 10854
rect 9774 10852 9798 10854
rect 9854 10852 9878 10854
rect 9934 10852 9958 10854
rect 10014 10852 10020 10854
rect 9712 10843 10020 10852
rect 10244 10742 10272 10950
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10266 7604 10610
rect 10060 10606 10088 10678
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8252 10364 8560 10373
rect 8252 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8498 10364
rect 8554 10362 8560 10364
rect 8314 10310 8316 10362
rect 8496 10310 8498 10362
rect 8252 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8498 10310
rect 8554 10308 8560 10310
rect 8252 10299 8560 10308
rect 8680 10266 8708 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 9784 10130 9812 10474
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10060 10062 10088 10542
rect 10244 10470 10272 10678
rect 11532 10674 11560 11154
rect 11900 11014 11928 11494
rect 11992 11218 12020 11630
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10810 11928 10950
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9178 7604 9454
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7668 9042 7696 9862
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6472 7886 6500 8298
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 7002 6500 7346
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5370 6040 5646
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5540 4694 5592 4700
rect 5552 4282 5580 4694
rect 5644 4678 5764 4706
rect 5816 4684 5868 4690
rect 5644 4486 5672 4678
rect 5816 4626 5868 4632
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5184 4185 5212 4218
rect 5170 4176 5226 4185
rect 5170 4111 5226 4120
rect 5644 4010 5672 4422
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5331 3836 5639 3845
rect 5331 3834 5337 3836
rect 5393 3834 5417 3836
rect 5473 3834 5497 3836
rect 5553 3834 5577 3836
rect 5633 3834 5639 3836
rect 5393 3782 5395 3834
rect 5575 3782 5577 3834
rect 5331 3780 5337 3782
rect 5393 3780 5417 3782
rect 5473 3780 5497 3782
rect 5553 3780 5577 3782
rect 5633 3780 5639 3782
rect 5331 3771 5639 3780
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5828 3670 5856 4626
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 4282 5948 4422
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5172 3664 5224 3670
rect 5092 3612 5172 3618
rect 5092 3606 5224 3612
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5092 3590 5212 3606
rect 5092 3534 5120 3590
rect 6012 3534 6040 3878
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 4816 3194 4844 3470
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4356 2514 4384 2994
rect 4724 2854 4752 2994
rect 5276 2972 5304 3334
rect 5368 3194 5396 3402
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5184 2944 5304 2972
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4448 2310 4476 2450
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 4448 1970 4476 2246
rect 4632 1986 4660 2246
rect 4724 2106 4752 2314
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 4632 1970 4752 1986
rect 4436 1964 4488 1970
rect 4632 1964 4764 1970
rect 4632 1958 4712 1964
rect 4436 1906 4488 1912
rect 4712 1906 4764 1912
rect 3884 1760 3936 1766
rect 3884 1702 3936 1708
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 3896 1426 3924 1702
rect 3884 1420 3936 1426
rect 3884 1362 3936 1368
rect 4724 1358 4752 1702
rect 4816 1358 4844 2246
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 4908 1562 4936 2042
rect 5184 1766 5212 2944
rect 5331 2748 5639 2757
rect 5331 2746 5337 2748
rect 5393 2746 5417 2748
rect 5473 2746 5497 2748
rect 5553 2746 5577 2748
rect 5633 2746 5639 2748
rect 5393 2694 5395 2746
rect 5575 2694 5577 2746
rect 5331 2692 5337 2694
rect 5393 2692 5417 2694
rect 5473 2692 5497 2694
rect 5553 2692 5577 2694
rect 5633 2692 5639 2694
rect 5331 2683 5639 2692
rect 5828 2514 5856 3334
rect 6104 2774 6132 4558
rect 6196 3602 6224 5238
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6380 3194 6408 5170
rect 6564 3398 6592 7142
rect 6656 6798 6684 7686
rect 6791 7644 7099 7653
rect 6791 7642 6797 7644
rect 6853 7642 6877 7644
rect 6933 7642 6957 7644
rect 7013 7642 7037 7644
rect 7093 7642 7099 7644
rect 6853 7590 6855 7642
rect 7035 7590 7037 7642
rect 6791 7588 6797 7590
rect 6853 7588 6877 7590
rect 6933 7588 6957 7590
rect 7013 7588 7037 7590
rect 7093 7588 7099 7590
rect 6791 7579 7099 7588
rect 7484 7206 7512 8842
rect 7668 8566 7696 8978
rect 7852 8922 7880 8978
rect 7760 8894 7880 8922
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7760 8294 7788 8894
rect 8128 8498 8156 9998
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8252 9276 8560 9285
rect 8252 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8498 9276
rect 8554 9274 8560 9276
rect 8314 9222 8316 9274
rect 8496 9222 8498 9274
rect 8252 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8498 9222
rect 8554 9220 8560 9222
rect 8252 9211 8560 9220
rect 8588 9178 8616 9862
rect 9712 9820 10020 9829
rect 9712 9818 9718 9820
rect 9774 9818 9798 9820
rect 9854 9818 9878 9820
rect 9934 9818 9958 9820
rect 10014 9818 10020 9820
rect 9774 9766 9776 9818
rect 9956 9766 9958 9818
rect 9712 9764 9718 9766
rect 9774 9764 9798 9766
rect 9854 9764 9878 9766
rect 9934 9764 9958 9766
rect 10014 9764 10020 9766
rect 9712 9755 10020 9764
rect 10060 9586 10088 9998
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 9178 8708 9318
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7342 7788 8230
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 7002 7512 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 5302 6684 6598
rect 6791 6556 7099 6565
rect 6791 6554 6797 6556
rect 6853 6554 6877 6556
rect 6933 6554 6957 6556
rect 7013 6554 7037 6556
rect 7093 6554 7099 6556
rect 6853 6502 6855 6554
rect 7035 6502 7037 6554
rect 6791 6500 6797 6502
rect 6853 6500 6877 6502
rect 6933 6500 6957 6502
rect 7013 6500 7037 6502
rect 7093 6500 7099 6502
rect 6791 6491 7099 6500
rect 7208 5642 7236 6666
rect 7392 5778 7420 6734
rect 7484 5914 7512 6938
rect 7760 6866 7788 7278
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7852 6798 7880 7822
rect 8036 7410 8064 8298
rect 8128 7478 8156 8434
rect 8312 8430 8340 8842
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8252 8188 8560 8197
rect 8252 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8498 8188
rect 8554 8186 8560 8188
rect 8314 8134 8316 8186
rect 8496 8134 8498 8186
rect 8252 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8498 8134
rect 8554 8132 8560 8134
rect 8252 8123 8560 8132
rect 8864 7886 8892 8774
rect 8956 8022 8984 8978
rect 9508 8974 9536 9522
rect 10060 9110 10088 9522
rect 10152 9450 10180 9998
rect 10244 9926 10272 10406
rect 11173 10364 11481 10373
rect 11173 10362 11179 10364
rect 11235 10362 11259 10364
rect 11315 10362 11339 10364
rect 11395 10362 11419 10364
rect 11475 10362 11481 10364
rect 11235 10310 11237 10362
rect 11417 10310 11419 10362
rect 11173 10308 11179 10310
rect 11235 10308 11259 10310
rect 11315 10308 11339 10310
rect 11395 10308 11419 10310
rect 11475 10308 11481 10310
rect 11173 10299 11481 10308
rect 11532 10266 11560 10610
rect 11900 10606 11928 10746
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 10266 11928 10542
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 9722 10272 9862
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7546 8800 7686
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8036 6730 8064 7346
rect 8252 7100 8560 7109
rect 8252 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8498 7100
rect 8554 7098 8560 7100
rect 8314 7046 8316 7098
rect 8496 7046 8498 7098
rect 8252 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8498 7046
rect 8554 7044 8560 7046
rect 8252 7035 8560 7044
rect 8588 6798 8616 7482
rect 8864 7410 8892 7822
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 6934 8984 7958
rect 9140 7886 9168 8910
rect 9712 8732 10020 8741
rect 9712 8730 9718 8732
rect 9774 8730 9798 8732
rect 9854 8730 9878 8732
rect 9934 8730 9958 8732
rect 10014 8730 10020 8732
rect 9774 8678 9776 8730
rect 9956 8678 9958 8730
rect 9712 8676 9718 8678
rect 9774 8676 9798 8678
rect 9854 8676 9878 8678
rect 9934 8676 9958 8678
rect 10014 8676 10020 8678
rect 9712 8667 10020 8676
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9232 7886 9260 8570
rect 9968 8090 9996 8570
rect 10060 8498 10088 9046
rect 10152 8906 10180 9386
rect 10980 9178 11008 9386
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 8974 11008 9114
rect 11072 9042 11100 9522
rect 11173 9276 11481 9285
rect 11173 9274 11179 9276
rect 11235 9274 11259 9276
rect 11315 9274 11339 9276
rect 11395 9274 11419 9276
rect 11475 9274 11481 9276
rect 11235 9222 11237 9274
rect 11417 9222 11419 9274
rect 11173 9220 11179 9222
rect 11235 9220 11259 9222
rect 11315 9220 11339 9222
rect 11395 9220 11419 9222
rect 11475 9220 11481 9222
rect 11173 9211 11481 9220
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8498 10180 8842
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10244 7970 10272 8774
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 8498 11100 8978
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11173 8188 11481 8197
rect 11173 8186 11179 8188
rect 11235 8186 11259 8188
rect 11315 8186 11339 8188
rect 11395 8186 11419 8188
rect 11475 8186 11481 8188
rect 11235 8134 11237 8186
rect 11417 8134 11419 8186
rect 11173 8132 11179 8134
rect 11235 8132 11259 8134
rect 11315 8132 11339 8134
rect 11395 8132 11419 8134
rect 11475 8132 11481 8134
rect 11173 8123 11481 8132
rect 9876 7942 10272 7970
rect 9876 7886 9904 7942
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8956 6458 8984 6870
rect 9140 6798 9168 7822
rect 9232 7342 9260 7822
rect 9712 7644 10020 7653
rect 9712 7642 9718 7644
rect 9774 7642 9798 7644
rect 9854 7642 9878 7644
rect 9934 7642 9958 7644
rect 10014 7642 10020 7644
rect 9774 7590 9776 7642
rect 9956 7590 9958 7642
rect 9712 7588 9718 7590
rect 9774 7588 9798 7590
rect 9854 7588 9878 7590
rect 9934 7588 9958 7590
rect 10014 7588 10020 7590
rect 9712 7579 10020 7588
rect 10060 7546 10088 7822
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9232 6798 9260 7278
rect 9876 6798 9904 7278
rect 10244 6798 10272 7942
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7002 11100 7686
rect 11173 7100 11481 7109
rect 11173 7098 11179 7100
rect 11235 7098 11259 7100
rect 11315 7098 11339 7100
rect 11395 7098 11419 7100
rect 11475 7098 11481 7100
rect 11235 7046 11237 7098
rect 11417 7046 11419 7098
rect 11173 7044 11179 7046
rect 11235 7044 11259 7046
rect 11315 7044 11339 7046
rect 11395 7044 11419 7046
rect 11475 7044 11481 7046
rect 11173 7035 11481 7044
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11072 6798 11100 6938
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9864 6792 9916 6798
rect 10232 6792 10284 6798
rect 9916 6752 10180 6780
rect 9864 6734 9916 6740
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8252 6012 8560 6021
rect 8252 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8498 6012
rect 8554 6010 8560 6012
rect 8314 5958 8316 6010
rect 8496 5958 8498 6010
rect 8252 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8498 5958
rect 8554 5956 8560 5958
rect 8252 5947 8560 5956
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6791 5468 7099 5477
rect 6791 5466 6797 5468
rect 6853 5466 6877 5468
rect 6933 5466 6957 5468
rect 7013 5466 7037 5468
rect 7093 5466 7099 5468
rect 6853 5414 6855 5466
rect 7035 5414 7037 5466
rect 6791 5412 6797 5414
rect 6853 5412 6877 5414
rect 6933 5412 6957 5414
rect 7013 5412 7037 5414
rect 7093 5412 7099 5414
rect 6791 5403 7099 5412
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 7208 5098 7236 5578
rect 7392 5234 7420 5714
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4826 6776 4966
rect 7024 4826 7052 5034
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6791 4380 7099 4389
rect 6791 4378 6797 4380
rect 6853 4378 6877 4380
rect 6933 4378 6957 4380
rect 7013 4378 7037 4380
rect 7093 4378 7099 4380
rect 6853 4326 6855 4378
rect 7035 4326 7037 4378
rect 6791 4324 6797 4326
rect 6853 4324 6877 4326
rect 6933 4324 6957 4326
rect 7013 4324 7037 4326
rect 7093 4324 7099 4326
rect 6791 4315 7099 4324
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6656 3194 6684 3606
rect 6791 3292 7099 3301
rect 6791 3290 6797 3292
rect 6853 3290 6877 3292
rect 6933 3290 6957 3292
rect 7013 3290 7037 3292
rect 7093 3290 7099 3292
rect 6853 3238 6855 3290
rect 7035 3238 7037 3290
rect 6791 3236 6797 3238
rect 6853 3236 6877 3238
rect 6933 3236 6957 3238
rect 7013 3236 7037 3238
rect 7093 3236 7099 3238
rect 6791 3227 7099 3236
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6012 2746 6132 2774
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6012 2038 6040 2746
rect 6196 2106 6224 2858
rect 6656 2774 6684 2858
rect 6840 2774 6868 3062
rect 7208 2922 7236 5034
rect 7484 5030 7512 5850
rect 8024 5704 8076 5710
rect 8300 5704 8352 5710
rect 8024 5646 8076 5652
rect 8298 5672 8300 5681
rect 8352 5672 8354 5681
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 8036 4826 8064 5646
rect 8298 5607 8354 5616
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8300 5364 8352 5370
rect 8404 5352 8432 5578
rect 8588 5574 8616 6190
rect 8680 5710 8708 6394
rect 9140 6254 9168 6734
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 5778 8892 6054
rect 9140 5914 9168 6190
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8668 5704 8720 5710
rect 9232 5681 9260 6734
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 8668 5646 8720 5652
rect 9218 5672 9274 5681
rect 9324 5642 9352 6054
rect 9416 5914 9444 6734
rect 9956 6656 10008 6662
rect 10008 6616 10088 6644
rect 9956 6598 10008 6604
rect 9712 6556 10020 6565
rect 9712 6554 9718 6556
rect 9774 6554 9798 6556
rect 9854 6554 9878 6556
rect 9934 6554 9958 6556
rect 10014 6554 10020 6556
rect 9774 6502 9776 6554
rect 9956 6502 9958 6554
rect 9712 6500 9718 6502
rect 9774 6500 9798 6502
rect 9854 6500 9878 6502
rect 9934 6500 9958 6502
rect 10014 6500 10020 6502
rect 9712 6491 10020 6500
rect 10060 6322 10088 6616
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9968 5710 9996 6054
rect 10152 5710 10180 6752
rect 10232 6734 10284 6740
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10244 6066 10272 6734
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6254 10364 6598
rect 11072 6458 11100 6734
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10244 6038 10364 6066
rect 10336 5710 10364 6038
rect 11173 6012 11481 6021
rect 11173 6010 11179 6012
rect 11235 6010 11259 6012
rect 11315 6010 11339 6012
rect 11395 6010 11419 6012
rect 11475 6010 11481 6012
rect 11235 5958 11237 6010
rect 11417 5958 11419 6010
rect 11173 5956 11179 5958
rect 11235 5956 11259 5958
rect 11315 5956 11339 5958
rect 11395 5956 11419 5958
rect 11475 5956 11481 5958
rect 11173 5947 11481 5956
rect 11532 5914 11560 9930
rect 11716 9586 11744 9998
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 12084 7954 12112 11630
rect 12633 10908 12941 10917
rect 12633 10906 12639 10908
rect 12695 10906 12719 10908
rect 12775 10906 12799 10908
rect 12855 10906 12879 10908
rect 12935 10906 12941 10908
rect 12695 10854 12697 10906
rect 12877 10854 12879 10906
rect 12633 10852 12639 10854
rect 12695 10852 12719 10854
rect 12775 10852 12799 10854
rect 12855 10852 12879 10854
rect 12935 10852 12941 10854
rect 12633 10843 12941 10852
rect 12633 9820 12941 9829
rect 12633 9818 12639 9820
rect 12695 9818 12719 9820
rect 12775 9818 12799 9820
rect 12855 9818 12879 9820
rect 12935 9818 12941 9820
rect 12695 9766 12697 9818
rect 12877 9766 12879 9818
rect 12633 9764 12639 9766
rect 12695 9764 12719 9766
rect 12775 9764 12799 9766
rect 12855 9764 12879 9766
rect 12935 9764 12941 9766
rect 12633 9755 12941 9764
rect 12633 8732 12941 8741
rect 12633 8730 12639 8732
rect 12695 8730 12719 8732
rect 12775 8730 12799 8732
rect 12855 8730 12879 8732
rect 12935 8730 12941 8732
rect 12695 8678 12697 8730
rect 12877 8678 12879 8730
rect 12633 8676 12639 8678
rect 12695 8676 12719 8678
rect 12775 8676 12799 8678
rect 12855 8676 12879 8678
rect 12935 8676 12941 8678
rect 12633 8667 12941 8676
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 6866 12112 7890
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7546 12480 7686
rect 12633 7644 12941 7653
rect 12633 7642 12639 7644
rect 12695 7642 12719 7644
rect 12775 7642 12799 7644
rect 12855 7642 12879 7644
rect 12935 7642 12941 7644
rect 12695 7590 12697 7642
rect 12877 7590 12879 7642
rect 12633 7588 12639 7590
rect 12695 7588 12719 7590
rect 12775 7588 12799 7590
rect 12855 7588 12879 7590
rect 12935 7588 12941 7590
rect 12633 7579 12941 7588
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6322 12112 6802
rect 12633 6556 12941 6565
rect 12633 6554 12639 6556
rect 12695 6554 12719 6556
rect 12775 6554 12799 6556
rect 12855 6554 12879 6556
rect 12935 6554 12941 6556
rect 12695 6502 12697 6554
rect 12877 6502 12879 6554
rect 12633 6500 12639 6502
rect 12695 6500 12719 6502
rect 12775 6500 12799 6502
rect 12855 6500 12879 6502
rect 12935 6500 12941 6502
rect 12633 6491 12941 6500
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11624 5778 11652 6258
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 5914 11928 6190
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 9680 5704 9732 5710
rect 9600 5664 9680 5692
rect 9218 5607 9220 5616
rect 9272 5607 9274 5616
rect 9312 5636 9364 5642
rect 9220 5578 9272 5584
rect 9312 5578 9364 5584
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8352 5324 8432 5352
rect 8484 5364 8536 5370
rect 8300 5306 8352 5312
rect 8484 5306 8536 5312
rect 8496 5166 8524 5306
rect 8680 5234 8708 5510
rect 9600 5302 9628 5664
rect 9680 5646 9732 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9712 5468 10020 5477
rect 9712 5466 9718 5468
rect 9774 5466 9798 5468
rect 9854 5466 9878 5468
rect 9934 5466 9958 5468
rect 10014 5466 10020 5468
rect 9774 5414 9776 5466
rect 9956 5414 9958 5466
rect 9712 5412 9718 5414
rect 9774 5412 9798 5414
rect 9854 5412 9878 5414
rect 9934 5412 9958 5414
rect 10014 5412 10020 5414
rect 9712 5403 10020 5412
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8252 4924 8560 4933
rect 8252 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8498 4924
rect 8554 4922 8560 4924
rect 8314 4870 8316 4922
rect 8496 4870 8498 4922
rect 8252 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8498 4870
rect 8554 4868 8560 4870
rect 8252 4859 8560 4868
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8588 4622 8616 4966
rect 8680 4826 8708 5170
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8680 4690 8708 4762
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8252 3836 8560 3845
rect 8252 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8498 3836
rect 8554 3834 8560 3836
rect 8314 3782 8316 3834
rect 8496 3782 8498 3834
rect 8252 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8498 3782
rect 8554 3780 8560 3782
rect 8252 3771 8560 3780
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3058 7420 3334
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6656 2746 6868 2774
rect 6184 2100 6236 2106
rect 6184 2042 6236 2048
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6656 1970 6684 2746
rect 7300 2446 7328 2790
rect 7484 2650 7512 2994
rect 8252 2748 8560 2757
rect 8252 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8498 2748
rect 8554 2746 8560 2748
rect 8314 2694 8316 2746
rect 8496 2694 8498 2746
rect 8252 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8498 2694
rect 8554 2692 8560 2694
rect 8252 2683 8560 2692
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 8588 2446 8616 4558
rect 8680 4146 8708 4626
rect 9416 4622 9444 5102
rect 9784 4826 9812 5306
rect 10060 5234 10088 5510
rect 10152 5234 10180 5510
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 4146 9444 4558
rect 9784 4486 9812 4762
rect 10060 4758 10088 5170
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9600 4282 9628 4422
rect 9712 4380 10020 4389
rect 9712 4378 9718 4380
rect 9774 4378 9798 4380
rect 9854 4378 9878 4380
rect 9934 4378 9958 4380
rect 10014 4378 10020 4380
rect 9774 4326 9776 4378
rect 9956 4326 9958 4378
rect 9712 4324 9718 4326
rect 9774 4324 9798 4326
rect 9854 4324 9878 4326
rect 9934 4324 9958 4326
rect 10014 4324 10020 4326
rect 9712 4315 10020 4324
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 10060 4146 10088 4694
rect 10152 4146 10180 5170
rect 10336 5030 10364 5646
rect 11532 5574 11560 5646
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 10980 5234 11008 5510
rect 11532 5370 11560 5510
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4690 10548 4966
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10244 3534 10272 4218
rect 10520 4146 10548 4626
rect 10888 4146 10916 4694
rect 10980 4146 11008 5170
rect 11173 4924 11481 4933
rect 11173 4922 11179 4924
rect 11235 4922 11259 4924
rect 11315 4922 11339 4924
rect 11395 4922 11419 4924
rect 11475 4922 11481 4924
rect 11235 4870 11237 4922
rect 11417 4870 11419 4922
rect 11173 4868 11179 4870
rect 11235 4868 11259 4870
rect 11315 4868 11339 4870
rect 11395 4868 11419 4870
rect 11475 4868 11481 4870
rect 11173 4859 11481 4868
rect 12084 4690 12112 5646
rect 12176 5370 12204 5646
rect 12633 5468 12941 5477
rect 12633 5466 12639 5468
rect 12695 5466 12719 5468
rect 12775 5466 12799 5468
rect 12855 5466 12879 5468
rect 12935 5466 12941 5468
rect 12695 5414 12697 5466
rect 12877 5414 12879 5466
rect 12633 5412 12639 5414
rect 12695 5412 12719 5414
rect 12775 5412 12799 5414
rect 12855 5412 12879 5414
rect 12935 5412 12941 5414
rect 12633 5403 12941 5412
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12176 4758 12204 5306
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11992 3942 12020 4422
rect 12084 4282 12112 4626
rect 12633 4380 12941 4389
rect 12633 4378 12639 4380
rect 12695 4378 12719 4380
rect 12775 4378 12799 4380
rect 12855 4378 12879 4380
rect 12935 4378 12941 4380
rect 12695 4326 12697 4378
rect 12877 4326 12879 4378
rect 12633 4324 12639 4326
rect 12695 4324 12719 4326
rect 12775 4324 12799 4326
rect 12855 4324 12879 4326
rect 12935 4324 12941 4326
rect 12633 4315 12941 4324
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 10336 3738 10364 3878
rect 11173 3836 11481 3845
rect 11173 3834 11179 3836
rect 11235 3834 11259 3836
rect 11315 3834 11339 3836
rect 11395 3834 11419 3836
rect 11475 3834 11481 3836
rect 11235 3782 11237 3834
rect 11417 3782 11419 3834
rect 11173 3780 11179 3782
rect 11235 3780 11259 3782
rect 11315 3780 11339 3782
rect 11395 3780 11419 3782
rect 11475 3780 11481 3782
rect 11173 3771 11481 3780
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 12084 3670 12112 4014
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 9712 3292 10020 3301
rect 9712 3290 9718 3292
rect 9774 3290 9798 3292
rect 9854 3290 9878 3292
rect 9934 3290 9958 3292
rect 10014 3290 10020 3292
rect 9774 3238 9776 3290
rect 9956 3238 9958 3290
rect 9712 3236 9718 3238
rect 9774 3236 9798 3238
rect 9854 3236 9878 3238
rect 9934 3236 9958 3238
rect 10014 3236 10020 3238
rect 9712 3227 10020 3236
rect 10796 3194 10824 3334
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8864 2774 8892 3062
rect 11072 3058 11100 3606
rect 12176 3602 12204 4014
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11256 2990 11284 3538
rect 12633 3292 12941 3301
rect 12633 3290 12639 3292
rect 12695 3290 12719 3292
rect 12775 3290 12799 3292
rect 12855 3290 12879 3292
rect 12935 3290 12941 3292
rect 12695 3238 12697 3290
rect 12877 3238 12879 3290
rect 12633 3236 12639 3238
rect 12695 3236 12719 3238
rect 12775 3236 12799 3238
rect 12855 3236 12879 3238
rect 12935 3236 12941 3238
rect 12633 3227 12941 3236
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 8680 2746 8892 2774
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 6791 2204 7099 2213
rect 6791 2202 6797 2204
rect 6853 2202 6877 2204
rect 6933 2202 6957 2204
rect 7013 2202 7037 2204
rect 7093 2202 7099 2204
rect 6853 2150 6855 2202
rect 7035 2150 7037 2202
rect 6791 2148 6797 2150
rect 6853 2148 6877 2150
rect 6933 2148 6957 2150
rect 7013 2148 7037 2150
rect 7093 2148 7099 2150
rect 6791 2139 7099 2148
rect 8680 2106 8708 2746
rect 9508 2446 9536 2790
rect 11173 2748 11481 2757
rect 11173 2746 11179 2748
rect 11235 2746 11259 2748
rect 11315 2746 11339 2748
rect 11395 2746 11419 2748
rect 11475 2746 11481 2748
rect 11235 2694 11237 2746
rect 11417 2694 11419 2746
rect 11173 2692 11179 2694
rect 11235 2692 11259 2694
rect 11315 2692 11339 2694
rect 11395 2692 11419 2694
rect 11475 2692 11481 2694
rect 11173 2683 11481 2692
rect 11624 2582 11652 2994
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11716 2446 11744 3130
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11808 2514 11836 2926
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 9712 2204 10020 2213
rect 9712 2202 9718 2204
rect 9774 2202 9798 2204
rect 9854 2202 9878 2204
rect 9934 2202 9958 2204
rect 10014 2202 10020 2204
rect 9774 2150 9776 2202
rect 9956 2150 9958 2202
rect 9712 2148 9718 2150
rect 9774 2148 9798 2150
rect 9854 2148 9878 2150
rect 9934 2148 9958 2150
rect 10014 2148 10020 2150
rect 9712 2139 10020 2148
rect 12633 2204 12941 2213
rect 12633 2202 12639 2204
rect 12695 2202 12719 2204
rect 12775 2202 12799 2204
rect 12855 2202 12879 2204
rect 12935 2202 12941 2204
rect 12695 2150 12697 2202
rect 12877 2150 12879 2202
rect 12633 2148 12639 2150
rect 12695 2148 12719 2150
rect 12775 2148 12799 2150
rect 12855 2148 12879 2150
rect 12935 2148 12941 2150
rect 12633 2139 12941 2148
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 6920 1828 6972 1834
rect 6920 1770 6972 1776
rect 4988 1760 5040 1766
rect 4988 1702 5040 1708
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 3804 649 3832 1294
rect 5000 1290 5028 1702
rect 4988 1284 5040 1290
rect 4988 1226 5040 1232
rect 5184 1222 5212 1702
rect 5331 1660 5639 1669
rect 5331 1658 5337 1660
rect 5393 1658 5417 1660
rect 5473 1658 5497 1660
rect 5553 1658 5577 1660
rect 5633 1658 5639 1660
rect 5393 1606 5395 1658
rect 5575 1606 5577 1658
rect 5331 1604 5337 1606
rect 5393 1604 5417 1606
rect 5473 1604 5497 1606
rect 5553 1604 5577 1606
rect 5633 1604 5639 1606
rect 5331 1595 5639 1604
rect 6932 1358 6960 1770
rect 7024 1562 7052 1906
rect 8252 1660 8560 1669
rect 8252 1658 8258 1660
rect 8314 1658 8338 1660
rect 8394 1658 8418 1660
rect 8474 1658 8498 1660
rect 8554 1658 8560 1660
rect 8314 1606 8316 1658
rect 8496 1606 8498 1658
rect 8252 1604 8258 1606
rect 8314 1604 8338 1606
rect 8394 1604 8418 1606
rect 8474 1604 8498 1606
rect 8554 1604 8560 1606
rect 8252 1595 8560 1604
rect 11173 1660 11481 1669
rect 11173 1658 11179 1660
rect 11235 1658 11259 1660
rect 11315 1658 11339 1660
rect 11395 1658 11419 1660
rect 11475 1658 11481 1660
rect 11235 1606 11237 1658
rect 11417 1606 11419 1658
rect 11173 1604 11179 1606
rect 11235 1604 11259 1606
rect 11315 1604 11339 1606
rect 11395 1604 11419 1606
rect 11475 1604 11481 1606
rect 11173 1595 11481 1604
rect 7012 1556 7064 1562
rect 7012 1498 7064 1504
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 3870 1116 4178 1125
rect 3870 1114 3876 1116
rect 3932 1114 3956 1116
rect 4012 1114 4036 1116
rect 4092 1114 4116 1116
rect 4172 1114 4178 1116
rect 3932 1062 3934 1114
rect 4114 1062 4116 1114
rect 3870 1060 3876 1062
rect 3932 1060 3956 1062
rect 4012 1060 4036 1062
rect 4092 1060 4116 1062
rect 4172 1060 4178 1062
rect 3870 1051 4178 1060
rect 6791 1116 7099 1125
rect 6791 1114 6797 1116
rect 6853 1114 6877 1116
rect 6933 1114 6957 1116
rect 7013 1114 7037 1116
rect 7093 1114 7099 1116
rect 6853 1062 6855 1114
rect 7035 1062 7037 1114
rect 6791 1060 6797 1062
rect 6853 1060 6877 1062
rect 6933 1060 6957 1062
rect 7013 1060 7037 1062
rect 7093 1060 7099 1062
rect 6791 1051 7099 1060
rect 9712 1116 10020 1125
rect 9712 1114 9718 1116
rect 9774 1114 9798 1116
rect 9854 1114 9878 1116
rect 9934 1114 9958 1116
rect 10014 1114 10020 1116
rect 9774 1062 9776 1114
rect 9956 1062 9958 1114
rect 9712 1060 9718 1062
rect 9774 1060 9798 1062
rect 9854 1060 9878 1062
rect 9934 1060 9958 1062
rect 10014 1060 10020 1062
rect 9712 1051 10020 1060
rect 12633 1116 12941 1125
rect 12633 1114 12639 1116
rect 12695 1114 12719 1116
rect 12775 1114 12799 1116
rect 12855 1114 12879 1116
rect 12935 1114 12941 1116
rect 12695 1062 12697 1114
rect 12877 1062 12879 1114
rect 12633 1060 12639 1062
rect 12695 1060 12719 1062
rect 12775 1060 12799 1062
rect 12855 1060 12879 1062
rect 12935 1060 12941 1062
rect 12633 1051 12941 1060
rect 3790 640 3846 649
rect 3790 575 3846 584
<< via2 >>
rect 4342 12824 4398 12880
rect 2416 12538 2472 12540
rect 2496 12538 2552 12540
rect 2576 12538 2632 12540
rect 2656 12538 2712 12540
rect 2416 12486 2462 12538
rect 2462 12486 2472 12538
rect 2496 12486 2526 12538
rect 2526 12486 2538 12538
rect 2538 12486 2552 12538
rect 2576 12486 2590 12538
rect 2590 12486 2602 12538
rect 2602 12486 2632 12538
rect 2656 12486 2666 12538
rect 2666 12486 2712 12538
rect 2416 12484 2472 12486
rect 2496 12484 2552 12486
rect 2576 12484 2632 12486
rect 2656 12484 2712 12486
rect 5337 12538 5393 12540
rect 5417 12538 5473 12540
rect 5497 12538 5553 12540
rect 5577 12538 5633 12540
rect 5337 12486 5383 12538
rect 5383 12486 5393 12538
rect 5417 12486 5447 12538
rect 5447 12486 5459 12538
rect 5459 12486 5473 12538
rect 5497 12486 5511 12538
rect 5511 12486 5523 12538
rect 5523 12486 5553 12538
rect 5577 12486 5587 12538
rect 5587 12486 5633 12538
rect 5337 12484 5393 12486
rect 5417 12484 5473 12486
rect 5497 12484 5553 12486
rect 5577 12484 5633 12486
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8498 12538 8554 12540
rect 8258 12486 8304 12538
rect 8304 12486 8314 12538
rect 8338 12486 8368 12538
rect 8368 12486 8380 12538
rect 8380 12486 8394 12538
rect 8418 12486 8432 12538
rect 8432 12486 8444 12538
rect 8444 12486 8474 12538
rect 8498 12486 8508 12538
rect 8508 12486 8554 12538
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8498 12484 8554 12486
rect 11179 12538 11235 12540
rect 11259 12538 11315 12540
rect 11339 12538 11395 12540
rect 11419 12538 11475 12540
rect 11179 12486 11225 12538
rect 11225 12486 11235 12538
rect 11259 12486 11289 12538
rect 11289 12486 11301 12538
rect 11301 12486 11315 12538
rect 11339 12486 11353 12538
rect 11353 12486 11365 12538
rect 11365 12486 11395 12538
rect 11419 12486 11429 12538
rect 11429 12486 11475 12538
rect 11179 12484 11235 12486
rect 11259 12484 11315 12486
rect 11339 12484 11395 12486
rect 11419 12484 11475 12486
rect 1306 12008 1362 12064
rect 3876 11994 3932 11996
rect 3956 11994 4012 11996
rect 4036 11994 4092 11996
rect 4116 11994 4172 11996
rect 3876 11942 3922 11994
rect 3922 11942 3932 11994
rect 3956 11942 3986 11994
rect 3986 11942 3998 11994
rect 3998 11942 4012 11994
rect 4036 11942 4050 11994
rect 4050 11942 4062 11994
rect 4062 11942 4092 11994
rect 4116 11942 4126 11994
rect 4126 11942 4172 11994
rect 3876 11940 3932 11942
rect 3956 11940 4012 11942
rect 4036 11940 4092 11942
rect 4116 11940 4172 11942
rect 2416 11450 2472 11452
rect 2496 11450 2552 11452
rect 2576 11450 2632 11452
rect 2656 11450 2712 11452
rect 2416 11398 2462 11450
rect 2462 11398 2472 11450
rect 2496 11398 2526 11450
rect 2526 11398 2538 11450
rect 2538 11398 2552 11450
rect 2576 11398 2590 11450
rect 2590 11398 2602 11450
rect 2602 11398 2632 11450
rect 2656 11398 2666 11450
rect 2666 11398 2712 11450
rect 2416 11396 2472 11398
rect 2496 11396 2552 11398
rect 2576 11396 2632 11398
rect 2656 11396 2712 11398
rect 1306 11192 1362 11248
rect 1766 10376 1822 10432
rect 1766 9560 1822 9616
rect 2416 10362 2472 10364
rect 2496 10362 2552 10364
rect 2576 10362 2632 10364
rect 2656 10362 2712 10364
rect 2416 10310 2462 10362
rect 2462 10310 2472 10362
rect 2496 10310 2526 10362
rect 2526 10310 2538 10362
rect 2538 10310 2552 10362
rect 2576 10310 2590 10362
rect 2590 10310 2602 10362
rect 2602 10310 2632 10362
rect 2656 10310 2666 10362
rect 2666 10310 2712 10362
rect 2416 10308 2472 10310
rect 2496 10308 2552 10310
rect 2576 10308 2632 10310
rect 2656 10308 2712 10310
rect 2416 9274 2472 9276
rect 2496 9274 2552 9276
rect 2576 9274 2632 9276
rect 2656 9274 2712 9276
rect 2416 9222 2462 9274
rect 2462 9222 2472 9274
rect 2496 9222 2526 9274
rect 2526 9222 2538 9274
rect 2538 9222 2552 9274
rect 2576 9222 2590 9274
rect 2590 9222 2602 9274
rect 2602 9222 2632 9274
rect 2656 9222 2666 9274
rect 2666 9222 2712 9274
rect 2416 9220 2472 9222
rect 2496 9220 2552 9222
rect 2576 9220 2632 9222
rect 2656 9220 2712 9222
rect 1306 8744 1362 8800
rect 1766 7928 1822 7984
rect 2416 8186 2472 8188
rect 2496 8186 2552 8188
rect 2576 8186 2632 8188
rect 2656 8186 2712 8188
rect 2416 8134 2462 8186
rect 2462 8134 2472 8186
rect 2496 8134 2526 8186
rect 2526 8134 2538 8186
rect 2538 8134 2552 8186
rect 2576 8134 2590 8186
rect 2590 8134 2602 8186
rect 2602 8134 2632 8186
rect 2656 8134 2666 8186
rect 2666 8134 2712 8186
rect 2416 8132 2472 8134
rect 2496 8132 2552 8134
rect 2576 8132 2632 8134
rect 2656 8132 2712 8134
rect 2042 7248 2098 7304
rect 1766 7112 1822 7168
rect 754 1400 810 1456
rect 2416 7098 2472 7100
rect 2496 7098 2552 7100
rect 2576 7098 2632 7100
rect 2656 7098 2712 7100
rect 2416 7046 2462 7098
rect 2462 7046 2472 7098
rect 2496 7046 2526 7098
rect 2526 7046 2538 7098
rect 2538 7046 2552 7098
rect 2576 7046 2590 7098
rect 2590 7046 2602 7098
rect 2602 7046 2632 7098
rect 2656 7046 2666 7098
rect 2666 7046 2712 7098
rect 2416 7044 2472 7046
rect 2496 7044 2552 7046
rect 2576 7044 2632 7046
rect 2656 7044 2712 7046
rect 6797 11994 6853 11996
rect 6877 11994 6933 11996
rect 6957 11994 7013 11996
rect 7037 11994 7093 11996
rect 6797 11942 6843 11994
rect 6843 11942 6853 11994
rect 6877 11942 6907 11994
rect 6907 11942 6919 11994
rect 6919 11942 6933 11994
rect 6957 11942 6971 11994
rect 6971 11942 6983 11994
rect 6983 11942 7013 11994
rect 7037 11942 7047 11994
rect 7047 11942 7093 11994
rect 6797 11940 6853 11942
rect 6877 11940 6933 11942
rect 6957 11940 7013 11942
rect 7037 11940 7093 11942
rect 9718 11994 9774 11996
rect 9798 11994 9854 11996
rect 9878 11994 9934 11996
rect 9958 11994 10014 11996
rect 9718 11942 9764 11994
rect 9764 11942 9774 11994
rect 9798 11942 9828 11994
rect 9828 11942 9840 11994
rect 9840 11942 9854 11994
rect 9878 11942 9892 11994
rect 9892 11942 9904 11994
rect 9904 11942 9934 11994
rect 9958 11942 9968 11994
rect 9968 11942 10014 11994
rect 9718 11940 9774 11942
rect 9798 11940 9854 11942
rect 9878 11940 9934 11942
rect 9958 11940 10014 11942
rect 12639 11994 12695 11996
rect 12719 11994 12775 11996
rect 12799 11994 12855 11996
rect 12879 11994 12935 11996
rect 12639 11942 12685 11994
rect 12685 11942 12695 11994
rect 12719 11942 12749 11994
rect 12749 11942 12761 11994
rect 12761 11942 12775 11994
rect 12799 11942 12813 11994
rect 12813 11942 12825 11994
rect 12825 11942 12855 11994
rect 12879 11942 12889 11994
rect 12889 11942 12935 11994
rect 12639 11940 12695 11942
rect 12719 11940 12775 11942
rect 12799 11940 12855 11942
rect 12879 11940 12935 11942
rect 5337 11450 5393 11452
rect 5417 11450 5473 11452
rect 5497 11450 5553 11452
rect 5577 11450 5633 11452
rect 5337 11398 5383 11450
rect 5383 11398 5393 11450
rect 5417 11398 5447 11450
rect 5447 11398 5459 11450
rect 5459 11398 5473 11450
rect 5497 11398 5511 11450
rect 5511 11398 5523 11450
rect 5523 11398 5553 11450
rect 5577 11398 5587 11450
rect 5587 11398 5633 11450
rect 5337 11396 5393 11398
rect 5417 11396 5473 11398
rect 5497 11396 5553 11398
rect 5577 11396 5633 11398
rect 2416 6010 2472 6012
rect 2496 6010 2552 6012
rect 2576 6010 2632 6012
rect 2656 6010 2712 6012
rect 2416 5958 2462 6010
rect 2462 5958 2472 6010
rect 2496 5958 2526 6010
rect 2526 5958 2538 6010
rect 2538 5958 2552 6010
rect 2576 5958 2590 6010
rect 2590 5958 2602 6010
rect 2602 5958 2632 6010
rect 2656 5958 2666 6010
rect 2666 5958 2712 6010
rect 2416 5956 2472 5958
rect 2496 5956 2552 5958
rect 2576 5956 2632 5958
rect 2656 5956 2712 5958
rect 2416 4922 2472 4924
rect 2496 4922 2552 4924
rect 2576 4922 2632 4924
rect 2656 4922 2712 4924
rect 2416 4870 2462 4922
rect 2462 4870 2472 4922
rect 2496 4870 2526 4922
rect 2526 4870 2538 4922
rect 2538 4870 2552 4922
rect 2576 4870 2590 4922
rect 2590 4870 2602 4922
rect 2602 4870 2632 4922
rect 2656 4870 2666 4922
rect 2666 4870 2712 4922
rect 2416 4868 2472 4870
rect 2496 4868 2552 4870
rect 2576 4868 2632 4870
rect 2656 4868 2712 4870
rect 2416 3834 2472 3836
rect 2496 3834 2552 3836
rect 2576 3834 2632 3836
rect 2656 3834 2712 3836
rect 2416 3782 2462 3834
rect 2462 3782 2472 3834
rect 2496 3782 2526 3834
rect 2526 3782 2538 3834
rect 2538 3782 2552 3834
rect 2576 3782 2590 3834
rect 2590 3782 2602 3834
rect 2602 3782 2632 3834
rect 2656 3782 2666 3834
rect 2666 3782 2712 3834
rect 2416 3780 2472 3782
rect 2496 3780 2552 3782
rect 2576 3780 2632 3782
rect 2656 3780 2712 3782
rect 2416 2746 2472 2748
rect 2496 2746 2552 2748
rect 2576 2746 2632 2748
rect 2656 2746 2712 2748
rect 2416 2694 2462 2746
rect 2462 2694 2472 2746
rect 2496 2694 2526 2746
rect 2526 2694 2538 2746
rect 2538 2694 2552 2746
rect 2576 2694 2590 2746
rect 2590 2694 2602 2746
rect 2602 2694 2632 2746
rect 2656 2694 2666 2746
rect 2666 2694 2712 2746
rect 2416 2692 2472 2694
rect 2496 2692 2552 2694
rect 2576 2692 2632 2694
rect 2656 2692 2712 2694
rect 2416 1658 2472 1660
rect 2496 1658 2552 1660
rect 2576 1658 2632 1660
rect 2656 1658 2712 1660
rect 2416 1606 2462 1658
rect 2462 1606 2472 1658
rect 2496 1606 2526 1658
rect 2526 1606 2538 1658
rect 2538 1606 2552 1658
rect 2576 1606 2590 1658
rect 2590 1606 2602 1658
rect 2602 1606 2632 1658
rect 2656 1606 2666 1658
rect 2666 1606 2712 1658
rect 2416 1604 2472 1606
rect 2496 1604 2552 1606
rect 2576 1604 2632 1606
rect 2656 1604 2712 1606
rect 3876 10906 3932 10908
rect 3956 10906 4012 10908
rect 4036 10906 4092 10908
rect 4116 10906 4172 10908
rect 3876 10854 3922 10906
rect 3922 10854 3932 10906
rect 3956 10854 3986 10906
rect 3986 10854 3998 10906
rect 3998 10854 4012 10906
rect 4036 10854 4050 10906
rect 4050 10854 4062 10906
rect 4062 10854 4092 10906
rect 4116 10854 4126 10906
rect 4126 10854 4172 10906
rect 3876 10852 3932 10854
rect 3956 10852 4012 10854
rect 4036 10852 4092 10854
rect 4116 10852 4172 10854
rect 3876 9818 3932 9820
rect 3956 9818 4012 9820
rect 4036 9818 4092 9820
rect 4116 9818 4172 9820
rect 3876 9766 3922 9818
rect 3922 9766 3932 9818
rect 3956 9766 3986 9818
rect 3986 9766 3998 9818
rect 3998 9766 4012 9818
rect 4036 9766 4050 9818
rect 4050 9766 4062 9818
rect 4062 9766 4092 9818
rect 4116 9766 4126 9818
rect 4126 9766 4172 9818
rect 3876 9764 3932 9766
rect 3956 9764 4012 9766
rect 4036 9764 4092 9766
rect 4116 9764 4172 9766
rect 5337 10362 5393 10364
rect 5417 10362 5473 10364
rect 5497 10362 5553 10364
rect 5577 10362 5633 10364
rect 5337 10310 5383 10362
rect 5383 10310 5393 10362
rect 5417 10310 5447 10362
rect 5447 10310 5459 10362
rect 5459 10310 5473 10362
rect 5497 10310 5511 10362
rect 5511 10310 5523 10362
rect 5523 10310 5553 10362
rect 5577 10310 5587 10362
rect 5587 10310 5633 10362
rect 5337 10308 5393 10310
rect 5417 10308 5473 10310
rect 5497 10308 5553 10310
rect 5577 10308 5633 10310
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8498 11450 8554 11452
rect 8258 11398 8304 11450
rect 8304 11398 8314 11450
rect 8338 11398 8368 11450
rect 8368 11398 8380 11450
rect 8380 11398 8394 11450
rect 8418 11398 8432 11450
rect 8432 11398 8444 11450
rect 8444 11398 8474 11450
rect 8498 11398 8508 11450
rect 8508 11398 8554 11450
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8498 11396 8554 11398
rect 11179 11450 11235 11452
rect 11259 11450 11315 11452
rect 11339 11450 11395 11452
rect 11419 11450 11475 11452
rect 11179 11398 11225 11450
rect 11225 11398 11235 11450
rect 11259 11398 11289 11450
rect 11289 11398 11301 11450
rect 11301 11398 11315 11450
rect 11339 11398 11353 11450
rect 11353 11398 11365 11450
rect 11365 11398 11395 11450
rect 11419 11398 11429 11450
rect 11429 11398 11475 11450
rect 11179 11396 11235 11398
rect 11259 11396 11315 11398
rect 11339 11396 11395 11398
rect 11419 11396 11475 11398
rect 3876 8730 3932 8732
rect 3956 8730 4012 8732
rect 4036 8730 4092 8732
rect 4116 8730 4172 8732
rect 3876 8678 3922 8730
rect 3922 8678 3932 8730
rect 3956 8678 3986 8730
rect 3986 8678 3998 8730
rect 3998 8678 4012 8730
rect 4036 8678 4050 8730
rect 4050 8678 4062 8730
rect 4062 8678 4092 8730
rect 4116 8678 4126 8730
rect 4126 8678 4172 8730
rect 3876 8676 3932 8678
rect 3956 8676 4012 8678
rect 4036 8676 4092 8678
rect 4116 8676 4172 8678
rect 3876 7642 3932 7644
rect 3956 7642 4012 7644
rect 4036 7642 4092 7644
rect 4116 7642 4172 7644
rect 3876 7590 3922 7642
rect 3922 7590 3932 7642
rect 3956 7590 3986 7642
rect 3986 7590 3998 7642
rect 3998 7590 4012 7642
rect 4036 7590 4050 7642
rect 4050 7590 4062 7642
rect 4062 7590 4092 7642
rect 4116 7590 4126 7642
rect 4126 7590 4172 7642
rect 3876 7588 3932 7590
rect 3956 7588 4012 7590
rect 4036 7588 4092 7590
rect 4116 7588 4172 7590
rect 5337 9274 5393 9276
rect 5417 9274 5473 9276
rect 5497 9274 5553 9276
rect 5577 9274 5633 9276
rect 5337 9222 5383 9274
rect 5383 9222 5393 9274
rect 5417 9222 5447 9274
rect 5447 9222 5459 9274
rect 5459 9222 5473 9274
rect 5497 9222 5511 9274
rect 5511 9222 5523 9274
rect 5523 9222 5553 9274
rect 5577 9222 5587 9274
rect 5587 9222 5633 9274
rect 5337 9220 5393 9222
rect 5417 9220 5473 9222
rect 5497 9220 5553 9222
rect 5577 9220 5633 9222
rect 5337 8186 5393 8188
rect 5417 8186 5473 8188
rect 5497 8186 5553 8188
rect 5577 8186 5633 8188
rect 5337 8134 5383 8186
rect 5383 8134 5393 8186
rect 5417 8134 5447 8186
rect 5447 8134 5459 8186
rect 5459 8134 5473 8186
rect 5497 8134 5511 8186
rect 5511 8134 5523 8186
rect 5523 8134 5553 8186
rect 5577 8134 5587 8186
rect 5587 8134 5633 8186
rect 5337 8132 5393 8134
rect 5417 8132 5473 8134
rect 5497 8132 5553 8134
rect 5577 8132 5633 8134
rect 5538 7268 5594 7304
rect 5538 7248 5540 7268
rect 5540 7248 5592 7268
rect 5592 7248 5594 7268
rect 5337 7098 5393 7100
rect 5417 7098 5473 7100
rect 5497 7098 5553 7100
rect 5577 7098 5633 7100
rect 5337 7046 5383 7098
rect 5383 7046 5393 7098
rect 5417 7046 5447 7098
rect 5447 7046 5459 7098
rect 5459 7046 5473 7098
rect 5497 7046 5511 7098
rect 5511 7046 5523 7098
rect 5523 7046 5553 7098
rect 5577 7046 5587 7098
rect 5587 7046 5633 7098
rect 5337 7044 5393 7046
rect 5417 7044 5473 7046
rect 5497 7044 5553 7046
rect 5577 7044 5633 7046
rect 3876 6554 3932 6556
rect 3956 6554 4012 6556
rect 4036 6554 4092 6556
rect 4116 6554 4172 6556
rect 3876 6502 3922 6554
rect 3922 6502 3932 6554
rect 3956 6502 3986 6554
rect 3986 6502 3998 6554
rect 3998 6502 4012 6554
rect 4036 6502 4050 6554
rect 4050 6502 4062 6554
rect 4062 6502 4092 6554
rect 4116 6502 4126 6554
rect 4126 6502 4172 6554
rect 3876 6500 3932 6502
rect 3956 6500 4012 6502
rect 4036 6500 4092 6502
rect 4116 6500 4172 6502
rect 3876 5466 3932 5468
rect 3956 5466 4012 5468
rect 4036 5466 4092 5468
rect 4116 5466 4172 5468
rect 3876 5414 3922 5466
rect 3922 5414 3932 5466
rect 3956 5414 3986 5466
rect 3986 5414 3998 5466
rect 3998 5414 4012 5466
rect 4036 5414 4050 5466
rect 4050 5414 4062 5466
rect 4062 5414 4092 5466
rect 4116 5414 4126 5466
rect 4126 5414 4172 5466
rect 3876 5412 3932 5414
rect 3956 5412 4012 5414
rect 4036 5412 4092 5414
rect 4116 5412 4172 5414
rect 3698 4140 3754 4176
rect 3698 4120 3700 4140
rect 3700 4120 3752 4140
rect 3752 4120 3754 4140
rect 3876 4378 3932 4380
rect 3956 4378 4012 4380
rect 4036 4378 4092 4380
rect 4116 4378 4172 4380
rect 3876 4326 3922 4378
rect 3922 4326 3932 4378
rect 3956 4326 3986 4378
rect 3986 4326 3998 4378
rect 3998 4326 4012 4378
rect 4036 4326 4050 4378
rect 4050 4326 4062 4378
rect 4062 4326 4092 4378
rect 4116 4326 4126 4378
rect 4126 4326 4172 4378
rect 3876 4324 3932 4326
rect 3956 4324 4012 4326
rect 4036 4324 4092 4326
rect 4116 4324 4172 4326
rect 3876 3290 3932 3292
rect 3956 3290 4012 3292
rect 4036 3290 4092 3292
rect 4116 3290 4172 3292
rect 3876 3238 3922 3290
rect 3922 3238 3932 3290
rect 3956 3238 3986 3290
rect 3986 3238 3998 3290
rect 3998 3238 4012 3290
rect 4036 3238 4050 3290
rect 4050 3238 4062 3290
rect 4062 3238 4092 3290
rect 4116 3238 4126 3290
rect 4126 3238 4172 3290
rect 3876 3236 3932 3238
rect 3956 3236 4012 3238
rect 4036 3236 4092 3238
rect 4116 3236 4172 3238
rect 3876 2202 3932 2204
rect 3956 2202 4012 2204
rect 4036 2202 4092 2204
rect 4116 2202 4172 2204
rect 3876 2150 3922 2202
rect 3922 2150 3932 2202
rect 3956 2150 3986 2202
rect 3986 2150 3998 2202
rect 3998 2150 4012 2202
rect 4036 2150 4050 2202
rect 4050 2150 4062 2202
rect 4062 2150 4092 2202
rect 4116 2150 4126 2202
rect 4126 2150 4172 2202
rect 3876 2148 3932 2150
rect 3956 2148 4012 2150
rect 4036 2148 4092 2150
rect 4116 2148 4172 2150
rect 5337 6010 5393 6012
rect 5417 6010 5473 6012
rect 5497 6010 5553 6012
rect 5577 6010 5633 6012
rect 5337 5958 5383 6010
rect 5383 5958 5393 6010
rect 5417 5958 5447 6010
rect 5447 5958 5459 6010
rect 5459 5958 5473 6010
rect 5497 5958 5511 6010
rect 5511 5958 5523 6010
rect 5523 5958 5553 6010
rect 5577 5958 5587 6010
rect 5587 5958 5633 6010
rect 5337 5956 5393 5958
rect 5417 5956 5473 5958
rect 5497 5956 5553 5958
rect 5577 5956 5633 5958
rect 5337 4922 5393 4924
rect 5417 4922 5473 4924
rect 5497 4922 5553 4924
rect 5577 4922 5633 4924
rect 5337 4870 5383 4922
rect 5383 4870 5393 4922
rect 5417 4870 5447 4922
rect 5447 4870 5459 4922
rect 5459 4870 5473 4922
rect 5497 4870 5511 4922
rect 5511 4870 5523 4922
rect 5523 4870 5553 4922
rect 5577 4870 5587 4922
rect 5587 4870 5633 4922
rect 5337 4868 5393 4870
rect 5417 4868 5473 4870
rect 5497 4868 5553 4870
rect 5577 4868 5633 4870
rect 6797 10906 6853 10908
rect 6877 10906 6933 10908
rect 6957 10906 7013 10908
rect 7037 10906 7093 10908
rect 6797 10854 6843 10906
rect 6843 10854 6853 10906
rect 6877 10854 6907 10906
rect 6907 10854 6919 10906
rect 6919 10854 6933 10906
rect 6957 10854 6971 10906
rect 6971 10854 6983 10906
rect 6983 10854 7013 10906
rect 7037 10854 7047 10906
rect 7047 10854 7093 10906
rect 6797 10852 6853 10854
rect 6877 10852 6933 10854
rect 6957 10852 7013 10854
rect 7037 10852 7093 10854
rect 6797 9818 6853 9820
rect 6877 9818 6933 9820
rect 6957 9818 7013 9820
rect 7037 9818 7093 9820
rect 6797 9766 6843 9818
rect 6843 9766 6853 9818
rect 6877 9766 6907 9818
rect 6907 9766 6919 9818
rect 6919 9766 6933 9818
rect 6957 9766 6971 9818
rect 6971 9766 6983 9818
rect 6983 9766 7013 9818
rect 7037 9766 7047 9818
rect 7047 9766 7093 9818
rect 6797 9764 6853 9766
rect 6877 9764 6933 9766
rect 6957 9764 7013 9766
rect 7037 9764 7093 9766
rect 6797 8730 6853 8732
rect 6877 8730 6933 8732
rect 6957 8730 7013 8732
rect 7037 8730 7093 8732
rect 6797 8678 6843 8730
rect 6843 8678 6853 8730
rect 6877 8678 6907 8730
rect 6907 8678 6919 8730
rect 6919 8678 6933 8730
rect 6957 8678 6971 8730
rect 6971 8678 6983 8730
rect 6983 8678 7013 8730
rect 7037 8678 7047 8730
rect 7047 8678 7093 8730
rect 6797 8676 6853 8678
rect 6877 8676 6933 8678
rect 6957 8676 7013 8678
rect 7037 8676 7093 8678
rect 9718 10906 9774 10908
rect 9798 10906 9854 10908
rect 9878 10906 9934 10908
rect 9958 10906 10014 10908
rect 9718 10854 9764 10906
rect 9764 10854 9774 10906
rect 9798 10854 9828 10906
rect 9828 10854 9840 10906
rect 9840 10854 9854 10906
rect 9878 10854 9892 10906
rect 9892 10854 9904 10906
rect 9904 10854 9934 10906
rect 9958 10854 9968 10906
rect 9968 10854 10014 10906
rect 9718 10852 9774 10854
rect 9798 10852 9854 10854
rect 9878 10852 9934 10854
rect 9958 10852 10014 10854
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8498 10362 8554 10364
rect 8258 10310 8304 10362
rect 8304 10310 8314 10362
rect 8338 10310 8368 10362
rect 8368 10310 8380 10362
rect 8380 10310 8394 10362
rect 8418 10310 8432 10362
rect 8432 10310 8444 10362
rect 8444 10310 8474 10362
rect 8498 10310 8508 10362
rect 8508 10310 8554 10362
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8498 10308 8554 10310
rect 5170 4120 5226 4176
rect 5337 3834 5393 3836
rect 5417 3834 5473 3836
rect 5497 3834 5553 3836
rect 5577 3834 5633 3836
rect 5337 3782 5383 3834
rect 5383 3782 5393 3834
rect 5417 3782 5447 3834
rect 5447 3782 5459 3834
rect 5459 3782 5473 3834
rect 5497 3782 5511 3834
rect 5511 3782 5523 3834
rect 5523 3782 5553 3834
rect 5577 3782 5587 3834
rect 5587 3782 5633 3834
rect 5337 3780 5393 3782
rect 5417 3780 5473 3782
rect 5497 3780 5553 3782
rect 5577 3780 5633 3782
rect 5337 2746 5393 2748
rect 5417 2746 5473 2748
rect 5497 2746 5553 2748
rect 5577 2746 5633 2748
rect 5337 2694 5383 2746
rect 5383 2694 5393 2746
rect 5417 2694 5447 2746
rect 5447 2694 5459 2746
rect 5459 2694 5473 2746
rect 5497 2694 5511 2746
rect 5511 2694 5523 2746
rect 5523 2694 5553 2746
rect 5577 2694 5587 2746
rect 5587 2694 5633 2746
rect 5337 2692 5393 2694
rect 5417 2692 5473 2694
rect 5497 2692 5553 2694
rect 5577 2692 5633 2694
rect 6797 7642 6853 7644
rect 6877 7642 6933 7644
rect 6957 7642 7013 7644
rect 7037 7642 7093 7644
rect 6797 7590 6843 7642
rect 6843 7590 6853 7642
rect 6877 7590 6907 7642
rect 6907 7590 6919 7642
rect 6919 7590 6933 7642
rect 6957 7590 6971 7642
rect 6971 7590 6983 7642
rect 6983 7590 7013 7642
rect 7037 7590 7047 7642
rect 7047 7590 7093 7642
rect 6797 7588 6853 7590
rect 6877 7588 6933 7590
rect 6957 7588 7013 7590
rect 7037 7588 7093 7590
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8498 9274 8554 9276
rect 8258 9222 8304 9274
rect 8304 9222 8314 9274
rect 8338 9222 8368 9274
rect 8368 9222 8380 9274
rect 8380 9222 8394 9274
rect 8418 9222 8432 9274
rect 8432 9222 8444 9274
rect 8444 9222 8474 9274
rect 8498 9222 8508 9274
rect 8508 9222 8554 9274
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8498 9220 8554 9222
rect 9718 9818 9774 9820
rect 9798 9818 9854 9820
rect 9878 9818 9934 9820
rect 9958 9818 10014 9820
rect 9718 9766 9764 9818
rect 9764 9766 9774 9818
rect 9798 9766 9828 9818
rect 9828 9766 9840 9818
rect 9840 9766 9854 9818
rect 9878 9766 9892 9818
rect 9892 9766 9904 9818
rect 9904 9766 9934 9818
rect 9958 9766 9968 9818
rect 9968 9766 10014 9818
rect 9718 9764 9774 9766
rect 9798 9764 9854 9766
rect 9878 9764 9934 9766
rect 9958 9764 10014 9766
rect 6797 6554 6853 6556
rect 6877 6554 6933 6556
rect 6957 6554 7013 6556
rect 7037 6554 7093 6556
rect 6797 6502 6843 6554
rect 6843 6502 6853 6554
rect 6877 6502 6907 6554
rect 6907 6502 6919 6554
rect 6919 6502 6933 6554
rect 6957 6502 6971 6554
rect 6971 6502 6983 6554
rect 6983 6502 7013 6554
rect 7037 6502 7047 6554
rect 7047 6502 7093 6554
rect 6797 6500 6853 6502
rect 6877 6500 6933 6502
rect 6957 6500 7013 6502
rect 7037 6500 7093 6502
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8498 8186 8554 8188
rect 8258 8134 8304 8186
rect 8304 8134 8314 8186
rect 8338 8134 8368 8186
rect 8368 8134 8380 8186
rect 8380 8134 8394 8186
rect 8418 8134 8432 8186
rect 8432 8134 8444 8186
rect 8444 8134 8474 8186
rect 8498 8134 8508 8186
rect 8508 8134 8554 8186
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 8498 8132 8554 8134
rect 11179 10362 11235 10364
rect 11259 10362 11315 10364
rect 11339 10362 11395 10364
rect 11419 10362 11475 10364
rect 11179 10310 11225 10362
rect 11225 10310 11235 10362
rect 11259 10310 11289 10362
rect 11289 10310 11301 10362
rect 11301 10310 11315 10362
rect 11339 10310 11353 10362
rect 11353 10310 11365 10362
rect 11365 10310 11395 10362
rect 11419 10310 11429 10362
rect 11429 10310 11475 10362
rect 11179 10308 11235 10310
rect 11259 10308 11315 10310
rect 11339 10308 11395 10310
rect 11419 10308 11475 10310
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8498 7098 8554 7100
rect 8258 7046 8304 7098
rect 8304 7046 8314 7098
rect 8338 7046 8368 7098
rect 8368 7046 8380 7098
rect 8380 7046 8394 7098
rect 8418 7046 8432 7098
rect 8432 7046 8444 7098
rect 8444 7046 8474 7098
rect 8498 7046 8508 7098
rect 8508 7046 8554 7098
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 8498 7044 8554 7046
rect 9718 8730 9774 8732
rect 9798 8730 9854 8732
rect 9878 8730 9934 8732
rect 9958 8730 10014 8732
rect 9718 8678 9764 8730
rect 9764 8678 9774 8730
rect 9798 8678 9828 8730
rect 9828 8678 9840 8730
rect 9840 8678 9854 8730
rect 9878 8678 9892 8730
rect 9892 8678 9904 8730
rect 9904 8678 9934 8730
rect 9958 8678 9968 8730
rect 9968 8678 10014 8730
rect 9718 8676 9774 8678
rect 9798 8676 9854 8678
rect 9878 8676 9934 8678
rect 9958 8676 10014 8678
rect 11179 9274 11235 9276
rect 11259 9274 11315 9276
rect 11339 9274 11395 9276
rect 11419 9274 11475 9276
rect 11179 9222 11225 9274
rect 11225 9222 11235 9274
rect 11259 9222 11289 9274
rect 11289 9222 11301 9274
rect 11301 9222 11315 9274
rect 11339 9222 11353 9274
rect 11353 9222 11365 9274
rect 11365 9222 11395 9274
rect 11419 9222 11429 9274
rect 11429 9222 11475 9274
rect 11179 9220 11235 9222
rect 11259 9220 11315 9222
rect 11339 9220 11395 9222
rect 11419 9220 11475 9222
rect 11179 8186 11235 8188
rect 11259 8186 11315 8188
rect 11339 8186 11395 8188
rect 11419 8186 11475 8188
rect 11179 8134 11225 8186
rect 11225 8134 11235 8186
rect 11259 8134 11289 8186
rect 11289 8134 11301 8186
rect 11301 8134 11315 8186
rect 11339 8134 11353 8186
rect 11353 8134 11365 8186
rect 11365 8134 11395 8186
rect 11419 8134 11429 8186
rect 11429 8134 11475 8186
rect 11179 8132 11235 8134
rect 11259 8132 11315 8134
rect 11339 8132 11395 8134
rect 11419 8132 11475 8134
rect 9718 7642 9774 7644
rect 9798 7642 9854 7644
rect 9878 7642 9934 7644
rect 9958 7642 10014 7644
rect 9718 7590 9764 7642
rect 9764 7590 9774 7642
rect 9798 7590 9828 7642
rect 9828 7590 9840 7642
rect 9840 7590 9854 7642
rect 9878 7590 9892 7642
rect 9892 7590 9904 7642
rect 9904 7590 9934 7642
rect 9958 7590 9968 7642
rect 9968 7590 10014 7642
rect 9718 7588 9774 7590
rect 9798 7588 9854 7590
rect 9878 7588 9934 7590
rect 9958 7588 10014 7590
rect 11179 7098 11235 7100
rect 11259 7098 11315 7100
rect 11339 7098 11395 7100
rect 11419 7098 11475 7100
rect 11179 7046 11225 7098
rect 11225 7046 11235 7098
rect 11259 7046 11289 7098
rect 11289 7046 11301 7098
rect 11301 7046 11315 7098
rect 11339 7046 11353 7098
rect 11353 7046 11365 7098
rect 11365 7046 11395 7098
rect 11419 7046 11429 7098
rect 11429 7046 11475 7098
rect 11179 7044 11235 7046
rect 11259 7044 11315 7046
rect 11339 7044 11395 7046
rect 11419 7044 11475 7046
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8498 6010 8554 6012
rect 8258 5958 8304 6010
rect 8304 5958 8314 6010
rect 8338 5958 8368 6010
rect 8368 5958 8380 6010
rect 8380 5958 8394 6010
rect 8418 5958 8432 6010
rect 8432 5958 8444 6010
rect 8444 5958 8474 6010
rect 8498 5958 8508 6010
rect 8508 5958 8554 6010
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8498 5956 8554 5958
rect 6797 5466 6853 5468
rect 6877 5466 6933 5468
rect 6957 5466 7013 5468
rect 7037 5466 7093 5468
rect 6797 5414 6843 5466
rect 6843 5414 6853 5466
rect 6877 5414 6907 5466
rect 6907 5414 6919 5466
rect 6919 5414 6933 5466
rect 6957 5414 6971 5466
rect 6971 5414 6983 5466
rect 6983 5414 7013 5466
rect 7037 5414 7047 5466
rect 7047 5414 7093 5466
rect 6797 5412 6853 5414
rect 6877 5412 6933 5414
rect 6957 5412 7013 5414
rect 7037 5412 7093 5414
rect 6797 4378 6853 4380
rect 6877 4378 6933 4380
rect 6957 4378 7013 4380
rect 7037 4378 7093 4380
rect 6797 4326 6843 4378
rect 6843 4326 6853 4378
rect 6877 4326 6907 4378
rect 6907 4326 6919 4378
rect 6919 4326 6933 4378
rect 6957 4326 6971 4378
rect 6971 4326 6983 4378
rect 6983 4326 7013 4378
rect 7037 4326 7047 4378
rect 7047 4326 7093 4378
rect 6797 4324 6853 4326
rect 6877 4324 6933 4326
rect 6957 4324 7013 4326
rect 7037 4324 7093 4326
rect 6797 3290 6853 3292
rect 6877 3290 6933 3292
rect 6957 3290 7013 3292
rect 7037 3290 7093 3292
rect 6797 3238 6843 3290
rect 6843 3238 6853 3290
rect 6877 3238 6907 3290
rect 6907 3238 6919 3290
rect 6919 3238 6933 3290
rect 6957 3238 6971 3290
rect 6971 3238 6983 3290
rect 6983 3238 7013 3290
rect 7037 3238 7047 3290
rect 7047 3238 7093 3290
rect 6797 3236 6853 3238
rect 6877 3236 6933 3238
rect 6957 3236 7013 3238
rect 7037 3236 7093 3238
rect 8298 5652 8300 5672
rect 8300 5652 8352 5672
rect 8352 5652 8354 5672
rect 8298 5616 8354 5652
rect 9218 5636 9274 5672
rect 9718 6554 9774 6556
rect 9798 6554 9854 6556
rect 9878 6554 9934 6556
rect 9958 6554 10014 6556
rect 9718 6502 9764 6554
rect 9764 6502 9774 6554
rect 9798 6502 9828 6554
rect 9828 6502 9840 6554
rect 9840 6502 9854 6554
rect 9878 6502 9892 6554
rect 9892 6502 9904 6554
rect 9904 6502 9934 6554
rect 9958 6502 9968 6554
rect 9968 6502 10014 6554
rect 9718 6500 9774 6502
rect 9798 6500 9854 6502
rect 9878 6500 9934 6502
rect 9958 6500 10014 6502
rect 11179 6010 11235 6012
rect 11259 6010 11315 6012
rect 11339 6010 11395 6012
rect 11419 6010 11475 6012
rect 11179 5958 11225 6010
rect 11225 5958 11235 6010
rect 11259 5958 11289 6010
rect 11289 5958 11301 6010
rect 11301 5958 11315 6010
rect 11339 5958 11353 6010
rect 11353 5958 11365 6010
rect 11365 5958 11395 6010
rect 11419 5958 11429 6010
rect 11429 5958 11475 6010
rect 11179 5956 11235 5958
rect 11259 5956 11315 5958
rect 11339 5956 11395 5958
rect 11419 5956 11475 5958
rect 12639 10906 12695 10908
rect 12719 10906 12775 10908
rect 12799 10906 12855 10908
rect 12879 10906 12935 10908
rect 12639 10854 12685 10906
rect 12685 10854 12695 10906
rect 12719 10854 12749 10906
rect 12749 10854 12761 10906
rect 12761 10854 12775 10906
rect 12799 10854 12813 10906
rect 12813 10854 12825 10906
rect 12825 10854 12855 10906
rect 12879 10854 12889 10906
rect 12889 10854 12935 10906
rect 12639 10852 12695 10854
rect 12719 10852 12775 10854
rect 12799 10852 12855 10854
rect 12879 10852 12935 10854
rect 12639 9818 12695 9820
rect 12719 9818 12775 9820
rect 12799 9818 12855 9820
rect 12879 9818 12935 9820
rect 12639 9766 12685 9818
rect 12685 9766 12695 9818
rect 12719 9766 12749 9818
rect 12749 9766 12761 9818
rect 12761 9766 12775 9818
rect 12799 9766 12813 9818
rect 12813 9766 12825 9818
rect 12825 9766 12855 9818
rect 12879 9766 12889 9818
rect 12889 9766 12935 9818
rect 12639 9764 12695 9766
rect 12719 9764 12775 9766
rect 12799 9764 12855 9766
rect 12879 9764 12935 9766
rect 12639 8730 12695 8732
rect 12719 8730 12775 8732
rect 12799 8730 12855 8732
rect 12879 8730 12935 8732
rect 12639 8678 12685 8730
rect 12685 8678 12695 8730
rect 12719 8678 12749 8730
rect 12749 8678 12761 8730
rect 12761 8678 12775 8730
rect 12799 8678 12813 8730
rect 12813 8678 12825 8730
rect 12825 8678 12855 8730
rect 12879 8678 12889 8730
rect 12889 8678 12935 8730
rect 12639 8676 12695 8678
rect 12719 8676 12775 8678
rect 12799 8676 12855 8678
rect 12879 8676 12935 8678
rect 12639 7642 12695 7644
rect 12719 7642 12775 7644
rect 12799 7642 12855 7644
rect 12879 7642 12935 7644
rect 12639 7590 12685 7642
rect 12685 7590 12695 7642
rect 12719 7590 12749 7642
rect 12749 7590 12761 7642
rect 12761 7590 12775 7642
rect 12799 7590 12813 7642
rect 12813 7590 12825 7642
rect 12825 7590 12855 7642
rect 12879 7590 12889 7642
rect 12889 7590 12935 7642
rect 12639 7588 12695 7590
rect 12719 7588 12775 7590
rect 12799 7588 12855 7590
rect 12879 7588 12935 7590
rect 12639 6554 12695 6556
rect 12719 6554 12775 6556
rect 12799 6554 12855 6556
rect 12879 6554 12935 6556
rect 12639 6502 12685 6554
rect 12685 6502 12695 6554
rect 12719 6502 12749 6554
rect 12749 6502 12761 6554
rect 12761 6502 12775 6554
rect 12799 6502 12813 6554
rect 12813 6502 12825 6554
rect 12825 6502 12855 6554
rect 12879 6502 12889 6554
rect 12889 6502 12935 6554
rect 12639 6500 12695 6502
rect 12719 6500 12775 6502
rect 12799 6500 12855 6502
rect 12879 6500 12935 6502
rect 9218 5616 9220 5636
rect 9220 5616 9272 5636
rect 9272 5616 9274 5636
rect 9718 5466 9774 5468
rect 9798 5466 9854 5468
rect 9878 5466 9934 5468
rect 9958 5466 10014 5468
rect 9718 5414 9764 5466
rect 9764 5414 9774 5466
rect 9798 5414 9828 5466
rect 9828 5414 9840 5466
rect 9840 5414 9854 5466
rect 9878 5414 9892 5466
rect 9892 5414 9904 5466
rect 9904 5414 9934 5466
rect 9958 5414 9968 5466
rect 9968 5414 10014 5466
rect 9718 5412 9774 5414
rect 9798 5412 9854 5414
rect 9878 5412 9934 5414
rect 9958 5412 10014 5414
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8498 4922 8554 4924
rect 8258 4870 8304 4922
rect 8304 4870 8314 4922
rect 8338 4870 8368 4922
rect 8368 4870 8380 4922
rect 8380 4870 8394 4922
rect 8418 4870 8432 4922
rect 8432 4870 8444 4922
rect 8444 4870 8474 4922
rect 8498 4870 8508 4922
rect 8508 4870 8554 4922
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8498 4868 8554 4870
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8498 3834 8554 3836
rect 8258 3782 8304 3834
rect 8304 3782 8314 3834
rect 8338 3782 8368 3834
rect 8368 3782 8380 3834
rect 8380 3782 8394 3834
rect 8418 3782 8432 3834
rect 8432 3782 8444 3834
rect 8444 3782 8474 3834
rect 8498 3782 8508 3834
rect 8508 3782 8554 3834
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 8498 3780 8554 3782
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8498 2746 8554 2748
rect 8258 2694 8304 2746
rect 8304 2694 8314 2746
rect 8338 2694 8368 2746
rect 8368 2694 8380 2746
rect 8380 2694 8394 2746
rect 8418 2694 8432 2746
rect 8432 2694 8444 2746
rect 8444 2694 8474 2746
rect 8498 2694 8508 2746
rect 8508 2694 8554 2746
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 8498 2692 8554 2694
rect 9718 4378 9774 4380
rect 9798 4378 9854 4380
rect 9878 4378 9934 4380
rect 9958 4378 10014 4380
rect 9718 4326 9764 4378
rect 9764 4326 9774 4378
rect 9798 4326 9828 4378
rect 9828 4326 9840 4378
rect 9840 4326 9854 4378
rect 9878 4326 9892 4378
rect 9892 4326 9904 4378
rect 9904 4326 9934 4378
rect 9958 4326 9968 4378
rect 9968 4326 10014 4378
rect 9718 4324 9774 4326
rect 9798 4324 9854 4326
rect 9878 4324 9934 4326
rect 9958 4324 10014 4326
rect 11179 4922 11235 4924
rect 11259 4922 11315 4924
rect 11339 4922 11395 4924
rect 11419 4922 11475 4924
rect 11179 4870 11225 4922
rect 11225 4870 11235 4922
rect 11259 4870 11289 4922
rect 11289 4870 11301 4922
rect 11301 4870 11315 4922
rect 11339 4870 11353 4922
rect 11353 4870 11365 4922
rect 11365 4870 11395 4922
rect 11419 4870 11429 4922
rect 11429 4870 11475 4922
rect 11179 4868 11235 4870
rect 11259 4868 11315 4870
rect 11339 4868 11395 4870
rect 11419 4868 11475 4870
rect 12639 5466 12695 5468
rect 12719 5466 12775 5468
rect 12799 5466 12855 5468
rect 12879 5466 12935 5468
rect 12639 5414 12685 5466
rect 12685 5414 12695 5466
rect 12719 5414 12749 5466
rect 12749 5414 12761 5466
rect 12761 5414 12775 5466
rect 12799 5414 12813 5466
rect 12813 5414 12825 5466
rect 12825 5414 12855 5466
rect 12879 5414 12889 5466
rect 12889 5414 12935 5466
rect 12639 5412 12695 5414
rect 12719 5412 12775 5414
rect 12799 5412 12855 5414
rect 12879 5412 12935 5414
rect 12639 4378 12695 4380
rect 12719 4378 12775 4380
rect 12799 4378 12855 4380
rect 12879 4378 12935 4380
rect 12639 4326 12685 4378
rect 12685 4326 12695 4378
rect 12719 4326 12749 4378
rect 12749 4326 12761 4378
rect 12761 4326 12775 4378
rect 12799 4326 12813 4378
rect 12813 4326 12825 4378
rect 12825 4326 12855 4378
rect 12879 4326 12889 4378
rect 12889 4326 12935 4378
rect 12639 4324 12695 4326
rect 12719 4324 12775 4326
rect 12799 4324 12855 4326
rect 12879 4324 12935 4326
rect 11179 3834 11235 3836
rect 11259 3834 11315 3836
rect 11339 3834 11395 3836
rect 11419 3834 11475 3836
rect 11179 3782 11225 3834
rect 11225 3782 11235 3834
rect 11259 3782 11289 3834
rect 11289 3782 11301 3834
rect 11301 3782 11315 3834
rect 11339 3782 11353 3834
rect 11353 3782 11365 3834
rect 11365 3782 11395 3834
rect 11419 3782 11429 3834
rect 11429 3782 11475 3834
rect 11179 3780 11235 3782
rect 11259 3780 11315 3782
rect 11339 3780 11395 3782
rect 11419 3780 11475 3782
rect 9718 3290 9774 3292
rect 9798 3290 9854 3292
rect 9878 3290 9934 3292
rect 9958 3290 10014 3292
rect 9718 3238 9764 3290
rect 9764 3238 9774 3290
rect 9798 3238 9828 3290
rect 9828 3238 9840 3290
rect 9840 3238 9854 3290
rect 9878 3238 9892 3290
rect 9892 3238 9904 3290
rect 9904 3238 9934 3290
rect 9958 3238 9968 3290
rect 9968 3238 10014 3290
rect 9718 3236 9774 3238
rect 9798 3236 9854 3238
rect 9878 3236 9934 3238
rect 9958 3236 10014 3238
rect 12639 3290 12695 3292
rect 12719 3290 12775 3292
rect 12799 3290 12855 3292
rect 12879 3290 12935 3292
rect 12639 3238 12685 3290
rect 12685 3238 12695 3290
rect 12719 3238 12749 3290
rect 12749 3238 12761 3290
rect 12761 3238 12775 3290
rect 12799 3238 12813 3290
rect 12813 3238 12825 3290
rect 12825 3238 12855 3290
rect 12879 3238 12889 3290
rect 12889 3238 12935 3290
rect 12639 3236 12695 3238
rect 12719 3236 12775 3238
rect 12799 3236 12855 3238
rect 12879 3236 12935 3238
rect 6797 2202 6853 2204
rect 6877 2202 6933 2204
rect 6957 2202 7013 2204
rect 7037 2202 7093 2204
rect 6797 2150 6843 2202
rect 6843 2150 6853 2202
rect 6877 2150 6907 2202
rect 6907 2150 6919 2202
rect 6919 2150 6933 2202
rect 6957 2150 6971 2202
rect 6971 2150 6983 2202
rect 6983 2150 7013 2202
rect 7037 2150 7047 2202
rect 7047 2150 7093 2202
rect 6797 2148 6853 2150
rect 6877 2148 6933 2150
rect 6957 2148 7013 2150
rect 7037 2148 7093 2150
rect 11179 2746 11235 2748
rect 11259 2746 11315 2748
rect 11339 2746 11395 2748
rect 11419 2746 11475 2748
rect 11179 2694 11225 2746
rect 11225 2694 11235 2746
rect 11259 2694 11289 2746
rect 11289 2694 11301 2746
rect 11301 2694 11315 2746
rect 11339 2694 11353 2746
rect 11353 2694 11365 2746
rect 11365 2694 11395 2746
rect 11419 2694 11429 2746
rect 11429 2694 11475 2746
rect 11179 2692 11235 2694
rect 11259 2692 11315 2694
rect 11339 2692 11395 2694
rect 11419 2692 11475 2694
rect 9718 2202 9774 2204
rect 9798 2202 9854 2204
rect 9878 2202 9934 2204
rect 9958 2202 10014 2204
rect 9718 2150 9764 2202
rect 9764 2150 9774 2202
rect 9798 2150 9828 2202
rect 9828 2150 9840 2202
rect 9840 2150 9854 2202
rect 9878 2150 9892 2202
rect 9892 2150 9904 2202
rect 9904 2150 9934 2202
rect 9958 2150 9968 2202
rect 9968 2150 10014 2202
rect 9718 2148 9774 2150
rect 9798 2148 9854 2150
rect 9878 2148 9934 2150
rect 9958 2148 10014 2150
rect 12639 2202 12695 2204
rect 12719 2202 12775 2204
rect 12799 2202 12855 2204
rect 12879 2202 12935 2204
rect 12639 2150 12685 2202
rect 12685 2150 12695 2202
rect 12719 2150 12749 2202
rect 12749 2150 12761 2202
rect 12761 2150 12775 2202
rect 12799 2150 12813 2202
rect 12813 2150 12825 2202
rect 12825 2150 12855 2202
rect 12879 2150 12889 2202
rect 12889 2150 12935 2202
rect 12639 2148 12695 2150
rect 12719 2148 12775 2150
rect 12799 2148 12855 2150
rect 12879 2148 12935 2150
rect 5337 1658 5393 1660
rect 5417 1658 5473 1660
rect 5497 1658 5553 1660
rect 5577 1658 5633 1660
rect 5337 1606 5383 1658
rect 5383 1606 5393 1658
rect 5417 1606 5447 1658
rect 5447 1606 5459 1658
rect 5459 1606 5473 1658
rect 5497 1606 5511 1658
rect 5511 1606 5523 1658
rect 5523 1606 5553 1658
rect 5577 1606 5587 1658
rect 5587 1606 5633 1658
rect 5337 1604 5393 1606
rect 5417 1604 5473 1606
rect 5497 1604 5553 1606
rect 5577 1604 5633 1606
rect 8258 1658 8314 1660
rect 8338 1658 8394 1660
rect 8418 1658 8474 1660
rect 8498 1658 8554 1660
rect 8258 1606 8304 1658
rect 8304 1606 8314 1658
rect 8338 1606 8368 1658
rect 8368 1606 8380 1658
rect 8380 1606 8394 1658
rect 8418 1606 8432 1658
rect 8432 1606 8444 1658
rect 8444 1606 8474 1658
rect 8498 1606 8508 1658
rect 8508 1606 8554 1658
rect 8258 1604 8314 1606
rect 8338 1604 8394 1606
rect 8418 1604 8474 1606
rect 8498 1604 8554 1606
rect 11179 1658 11235 1660
rect 11259 1658 11315 1660
rect 11339 1658 11395 1660
rect 11419 1658 11475 1660
rect 11179 1606 11225 1658
rect 11225 1606 11235 1658
rect 11259 1606 11289 1658
rect 11289 1606 11301 1658
rect 11301 1606 11315 1658
rect 11339 1606 11353 1658
rect 11353 1606 11365 1658
rect 11365 1606 11395 1658
rect 11419 1606 11429 1658
rect 11429 1606 11475 1658
rect 11179 1604 11235 1606
rect 11259 1604 11315 1606
rect 11339 1604 11395 1606
rect 11419 1604 11475 1606
rect 3876 1114 3932 1116
rect 3956 1114 4012 1116
rect 4036 1114 4092 1116
rect 4116 1114 4172 1116
rect 3876 1062 3922 1114
rect 3922 1062 3932 1114
rect 3956 1062 3986 1114
rect 3986 1062 3998 1114
rect 3998 1062 4012 1114
rect 4036 1062 4050 1114
rect 4050 1062 4062 1114
rect 4062 1062 4092 1114
rect 4116 1062 4126 1114
rect 4126 1062 4172 1114
rect 3876 1060 3932 1062
rect 3956 1060 4012 1062
rect 4036 1060 4092 1062
rect 4116 1060 4172 1062
rect 6797 1114 6853 1116
rect 6877 1114 6933 1116
rect 6957 1114 7013 1116
rect 7037 1114 7093 1116
rect 6797 1062 6843 1114
rect 6843 1062 6853 1114
rect 6877 1062 6907 1114
rect 6907 1062 6919 1114
rect 6919 1062 6933 1114
rect 6957 1062 6971 1114
rect 6971 1062 6983 1114
rect 6983 1062 7013 1114
rect 7037 1062 7047 1114
rect 7047 1062 7093 1114
rect 6797 1060 6853 1062
rect 6877 1060 6933 1062
rect 6957 1060 7013 1062
rect 7037 1060 7093 1062
rect 9718 1114 9774 1116
rect 9798 1114 9854 1116
rect 9878 1114 9934 1116
rect 9958 1114 10014 1116
rect 9718 1062 9764 1114
rect 9764 1062 9774 1114
rect 9798 1062 9828 1114
rect 9828 1062 9840 1114
rect 9840 1062 9854 1114
rect 9878 1062 9892 1114
rect 9892 1062 9904 1114
rect 9904 1062 9934 1114
rect 9958 1062 9968 1114
rect 9968 1062 10014 1114
rect 9718 1060 9774 1062
rect 9798 1060 9854 1062
rect 9878 1060 9934 1062
rect 9958 1060 10014 1062
rect 12639 1114 12695 1116
rect 12719 1114 12775 1116
rect 12799 1114 12855 1116
rect 12879 1114 12935 1116
rect 12639 1062 12685 1114
rect 12685 1062 12695 1114
rect 12719 1062 12749 1114
rect 12749 1062 12761 1114
rect 12761 1062 12775 1114
rect 12799 1062 12813 1114
rect 12813 1062 12825 1114
rect 12825 1062 12855 1114
rect 12879 1062 12889 1114
rect 12889 1062 12935 1114
rect 12639 1060 12695 1062
rect 12719 1060 12775 1062
rect 12799 1060 12855 1062
rect 12879 1060 12935 1062
rect 3790 584 3846 640
<< metal3 >>
rect 0 12882 400 12912
rect 4337 12882 4403 12885
rect 0 12880 4403 12882
rect 0 12824 4342 12880
rect 4398 12824 4403 12880
rect 0 12822 4403 12824
rect 0 12792 400 12822
rect 4337 12819 4403 12822
rect 2406 12544 2722 12545
rect 2406 12480 2412 12544
rect 2476 12480 2492 12544
rect 2556 12480 2572 12544
rect 2636 12480 2652 12544
rect 2716 12480 2722 12544
rect 2406 12479 2722 12480
rect 5327 12544 5643 12545
rect 5327 12480 5333 12544
rect 5397 12480 5413 12544
rect 5477 12480 5493 12544
rect 5557 12480 5573 12544
rect 5637 12480 5643 12544
rect 5327 12479 5643 12480
rect 8248 12544 8564 12545
rect 8248 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8494 12544
rect 8558 12480 8564 12544
rect 8248 12479 8564 12480
rect 11169 12544 11485 12545
rect 11169 12480 11175 12544
rect 11239 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11485 12544
rect 11169 12479 11485 12480
rect 0 12066 400 12096
rect 1301 12066 1367 12069
rect 0 12064 1367 12066
rect 0 12008 1306 12064
rect 1362 12008 1367 12064
rect 0 12006 1367 12008
rect 0 11976 400 12006
rect 1301 12003 1367 12006
rect 3866 12000 4182 12001
rect 3866 11936 3872 12000
rect 3936 11936 3952 12000
rect 4016 11936 4032 12000
rect 4096 11936 4112 12000
rect 4176 11936 4182 12000
rect 3866 11935 4182 11936
rect 6787 12000 7103 12001
rect 6787 11936 6793 12000
rect 6857 11936 6873 12000
rect 6937 11936 6953 12000
rect 7017 11936 7033 12000
rect 7097 11936 7103 12000
rect 6787 11935 7103 11936
rect 9708 12000 10024 12001
rect 9708 11936 9714 12000
rect 9778 11936 9794 12000
rect 9858 11936 9874 12000
rect 9938 11936 9954 12000
rect 10018 11936 10024 12000
rect 9708 11935 10024 11936
rect 12629 12000 12945 12001
rect 12629 11936 12635 12000
rect 12699 11936 12715 12000
rect 12779 11936 12795 12000
rect 12859 11936 12875 12000
rect 12939 11936 12945 12000
rect 12629 11935 12945 11936
rect 2406 11456 2722 11457
rect 2406 11392 2412 11456
rect 2476 11392 2492 11456
rect 2556 11392 2572 11456
rect 2636 11392 2652 11456
rect 2716 11392 2722 11456
rect 2406 11391 2722 11392
rect 5327 11456 5643 11457
rect 5327 11392 5333 11456
rect 5397 11392 5413 11456
rect 5477 11392 5493 11456
rect 5557 11392 5573 11456
rect 5637 11392 5643 11456
rect 5327 11391 5643 11392
rect 8248 11456 8564 11457
rect 8248 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8494 11456
rect 8558 11392 8564 11456
rect 8248 11391 8564 11392
rect 11169 11456 11485 11457
rect 11169 11392 11175 11456
rect 11239 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11485 11456
rect 11169 11391 11485 11392
rect 0 11250 400 11280
rect 1301 11250 1367 11253
rect 0 11248 1367 11250
rect 0 11192 1306 11248
rect 1362 11192 1367 11248
rect 0 11190 1367 11192
rect 0 11160 400 11190
rect 1301 11187 1367 11190
rect 3866 10912 4182 10913
rect 3866 10848 3872 10912
rect 3936 10848 3952 10912
rect 4016 10848 4032 10912
rect 4096 10848 4112 10912
rect 4176 10848 4182 10912
rect 3866 10847 4182 10848
rect 6787 10912 7103 10913
rect 6787 10848 6793 10912
rect 6857 10848 6873 10912
rect 6937 10848 6953 10912
rect 7017 10848 7033 10912
rect 7097 10848 7103 10912
rect 6787 10847 7103 10848
rect 9708 10912 10024 10913
rect 9708 10848 9714 10912
rect 9778 10848 9794 10912
rect 9858 10848 9874 10912
rect 9938 10848 9954 10912
rect 10018 10848 10024 10912
rect 9708 10847 10024 10848
rect 12629 10912 12945 10913
rect 12629 10848 12635 10912
rect 12699 10848 12715 10912
rect 12779 10848 12795 10912
rect 12859 10848 12875 10912
rect 12939 10848 12945 10912
rect 12629 10847 12945 10848
rect 0 10434 400 10464
rect 1761 10434 1827 10437
rect 0 10432 1827 10434
rect 0 10376 1766 10432
rect 1822 10376 1827 10432
rect 0 10374 1827 10376
rect 0 10344 400 10374
rect 1761 10371 1827 10374
rect 2406 10368 2722 10369
rect 2406 10304 2412 10368
rect 2476 10304 2492 10368
rect 2556 10304 2572 10368
rect 2636 10304 2652 10368
rect 2716 10304 2722 10368
rect 2406 10303 2722 10304
rect 5327 10368 5643 10369
rect 5327 10304 5333 10368
rect 5397 10304 5413 10368
rect 5477 10304 5493 10368
rect 5557 10304 5573 10368
rect 5637 10304 5643 10368
rect 5327 10303 5643 10304
rect 8248 10368 8564 10369
rect 8248 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8494 10368
rect 8558 10304 8564 10368
rect 8248 10303 8564 10304
rect 11169 10368 11485 10369
rect 11169 10304 11175 10368
rect 11239 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11485 10368
rect 11169 10303 11485 10304
rect 3866 9824 4182 9825
rect 3866 9760 3872 9824
rect 3936 9760 3952 9824
rect 4016 9760 4032 9824
rect 4096 9760 4112 9824
rect 4176 9760 4182 9824
rect 3866 9759 4182 9760
rect 6787 9824 7103 9825
rect 6787 9760 6793 9824
rect 6857 9760 6873 9824
rect 6937 9760 6953 9824
rect 7017 9760 7033 9824
rect 7097 9760 7103 9824
rect 6787 9759 7103 9760
rect 9708 9824 10024 9825
rect 9708 9760 9714 9824
rect 9778 9760 9794 9824
rect 9858 9760 9874 9824
rect 9938 9760 9954 9824
rect 10018 9760 10024 9824
rect 9708 9759 10024 9760
rect 12629 9824 12945 9825
rect 12629 9760 12635 9824
rect 12699 9760 12715 9824
rect 12779 9760 12795 9824
rect 12859 9760 12875 9824
rect 12939 9760 12945 9824
rect 12629 9759 12945 9760
rect 0 9618 400 9648
rect 1761 9618 1827 9621
rect 0 9616 1827 9618
rect 0 9560 1766 9616
rect 1822 9560 1827 9616
rect 0 9558 1827 9560
rect 0 9528 400 9558
rect 1761 9555 1827 9558
rect 2406 9280 2722 9281
rect 2406 9216 2412 9280
rect 2476 9216 2492 9280
rect 2556 9216 2572 9280
rect 2636 9216 2652 9280
rect 2716 9216 2722 9280
rect 2406 9215 2722 9216
rect 5327 9280 5643 9281
rect 5327 9216 5333 9280
rect 5397 9216 5413 9280
rect 5477 9216 5493 9280
rect 5557 9216 5573 9280
rect 5637 9216 5643 9280
rect 5327 9215 5643 9216
rect 8248 9280 8564 9281
rect 8248 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8494 9280
rect 8558 9216 8564 9280
rect 8248 9215 8564 9216
rect 11169 9280 11485 9281
rect 11169 9216 11175 9280
rect 11239 9216 11255 9280
rect 11319 9216 11335 9280
rect 11399 9216 11415 9280
rect 11479 9216 11485 9280
rect 11169 9215 11485 9216
rect 0 8802 400 8832
rect 1301 8802 1367 8805
rect 0 8800 1367 8802
rect 0 8744 1306 8800
rect 1362 8744 1367 8800
rect 0 8742 1367 8744
rect 0 8712 400 8742
rect 1301 8739 1367 8742
rect 3866 8736 4182 8737
rect 3866 8672 3872 8736
rect 3936 8672 3952 8736
rect 4016 8672 4032 8736
rect 4096 8672 4112 8736
rect 4176 8672 4182 8736
rect 3866 8671 4182 8672
rect 6787 8736 7103 8737
rect 6787 8672 6793 8736
rect 6857 8672 6873 8736
rect 6937 8672 6953 8736
rect 7017 8672 7033 8736
rect 7097 8672 7103 8736
rect 6787 8671 7103 8672
rect 9708 8736 10024 8737
rect 9708 8672 9714 8736
rect 9778 8672 9794 8736
rect 9858 8672 9874 8736
rect 9938 8672 9954 8736
rect 10018 8672 10024 8736
rect 9708 8671 10024 8672
rect 12629 8736 12945 8737
rect 12629 8672 12635 8736
rect 12699 8672 12715 8736
rect 12779 8672 12795 8736
rect 12859 8672 12875 8736
rect 12939 8672 12945 8736
rect 12629 8671 12945 8672
rect 2406 8192 2722 8193
rect 2406 8128 2412 8192
rect 2476 8128 2492 8192
rect 2556 8128 2572 8192
rect 2636 8128 2652 8192
rect 2716 8128 2722 8192
rect 2406 8127 2722 8128
rect 5327 8192 5643 8193
rect 5327 8128 5333 8192
rect 5397 8128 5413 8192
rect 5477 8128 5493 8192
rect 5557 8128 5573 8192
rect 5637 8128 5643 8192
rect 5327 8127 5643 8128
rect 8248 8192 8564 8193
rect 8248 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8494 8192
rect 8558 8128 8564 8192
rect 8248 8127 8564 8128
rect 11169 8192 11485 8193
rect 11169 8128 11175 8192
rect 11239 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11485 8192
rect 11169 8127 11485 8128
rect 0 7986 400 8016
rect 1761 7986 1827 7989
rect 0 7984 1827 7986
rect 0 7928 1766 7984
rect 1822 7928 1827 7984
rect 0 7926 1827 7928
rect 0 7896 400 7926
rect 1761 7923 1827 7926
rect 3866 7648 4182 7649
rect 3866 7584 3872 7648
rect 3936 7584 3952 7648
rect 4016 7584 4032 7648
rect 4096 7584 4112 7648
rect 4176 7584 4182 7648
rect 3866 7583 4182 7584
rect 6787 7648 7103 7649
rect 6787 7584 6793 7648
rect 6857 7584 6873 7648
rect 6937 7584 6953 7648
rect 7017 7584 7033 7648
rect 7097 7584 7103 7648
rect 6787 7583 7103 7584
rect 9708 7648 10024 7649
rect 9708 7584 9714 7648
rect 9778 7584 9794 7648
rect 9858 7584 9874 7648
rect 9938 7584 9954 7648
rect 10018 7584 10024 7648
rect 9708 7583 10024 7584
rect 12629 7648 12945 7649
rect 12629 7584 12635 7648
rect 12699 7584 12715 7648
rect 12779 7584 12795 7648
rect 12859 7584 12875 7648
rect 12939 7584 12945 7648
rect 12629 7583 12945 7584
rect 2037 7306 2103 7309
rect 5533 7306 5599 7309
rect 2037 7304 5599 7306
rect 2037 7248 2042 7304
rect 2098 7248 5538 7304
rect 5594 7248 5599 7304
rect 2037 7246 5599 7248
rect 2037 7243 2103 7246
rect 5533 7243 5599 7246
rect 0 7170 400 7200
rect 1761 7170 1827 7173
rect 0 7168 1827 7170
rect 0 7112 1766 7168
rect 1822 7112 1827 7168
rect 0 7110 1827 7112
rect 0 7080 400 7110
rect 1761 7107 1827 7110
rect 2406 7104 2722 7105
rect 2406 7040 2412 7104
rect 2476 7040 2492 7104
rect 2556 7040 2572 7104
rect 2636 7040 2652 7104
rect 2716 7040 2722 7104
rect 2406 7039 2722 7040
rect 5327 7104 5643 7105
rect 5327 7040 5333 7104
rect 5397 7040 5413 7104
rect 5477 7040 5493 7104
rect 5557 7040 5573 7104
rect 5637 7040 5643 7104
rect 5327 7039 5643 7040
rect 8248 7104 8564 7105
rect 8248 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8494 7104
rect 8558 7040 8564 7104
rect 8248 7039 8564 7040
rect 11169 7104 11485 7105
rect 11169 7040 11175 7104
rect 11239 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11485 7104
rect 11169 7039 11485 7040
rect 3866 6560 4182 6561
rect 3866 6496 3872 6560
rect 3936 6496 3952 6560
rect 4016 6496 4032 6560
rect 4096 6496 4112 6560
rect 4176 6496 4182 6560
rect 3866 6495 4182 6496
rect 6787 6560 7103 6561
rect 6787 6496 6793 6560
rect 6857 6496 6873 6560
rect 6937 6496 6953 6560
rect 7017 6496 7033 6560
rect 7097 6496 7103 6560
rect 6787 6495 7103 6496
rect 9708 6560 10024 6561
rect 9708 6496 9714 6560
rect 9778 6496 9794 6560
rect 9858 6496 9874 6560
rect 9938 6496 9954 6560
rect 10018 6496 10024 6560
rect 9708 6495 10024 6496
rect 12629 6560 12945 6561
rect 12629 6496 12635 6560
rect 12699 6496 12715 6560
rect 12779 6496 12795 6560
rect 12859 6496 12875 6560
rect 12939 6496 12945 6560
rect 12629 6495 12945 6496
rect 0 6264 400 6384
rect 2406 6016 2722 6017
rect 2406 5952 2412 6016
rect 2476 5952 2492 6016
rect 2556 5952 2572 6016
rect 2636 5952 2652 6016
rect 2716 5952 2722 6016
rect 2406 5951 2722 5952
rect 5327 6016 5643 6017
rect 5327 5952 5333 6016
rect 5397 5952 5413 6016
rect 5477 5952 5493 6016
rect 5557 5952 5573 6016
rect 5637 5952 5643 6016
rect 5327 5951 5643 5952
rect 8248 6016 8564 6017
rect 8248 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8494 6016
rect 8558 5952 8564 6016
rect 8248 5951 8564 5952
rect 11169 6016 11485 6017
rect 11169 5952 11175 6016
rect 11239 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11485 6016
rect 11169 5951 11485 5952
rect 8293 5674 8359 5677
rect 9213 5674 9279 5677
rect 8293 5672 9279 5674
rect 8293 5616 8298 5672
rect 8354 5616 9218 5672
rect 9274 5616 9279 5672
rect 8293 5614 9279 5616
rect 8293 5611 8359 5614
rect 9213 5611 9279 5614
rect 0 5448 400 5568
rect 3866 5472 4182 5473
rect 3866 5408 3872 5472
rect 3936 5408 3952 5472
rect 4016 5408 4032 5472
rect 4096 5408 4112 5472
rect 4176 5408 4182 5472
rect 3866 5407 4182 5408
rect 6787 5472 7103 5473
rect 6787 5408 6793 5472
rect 6857 5408 6873 5472
rect 6937 5408 6953 5472
rect 7017 5408 7033 5472
rect 7097 5408 7103 5472
rect 6787 5407 7103 5408
rect 9708 5472 10024 5473
rect 9708 5408 9714 5472
rect 9778 5408 9794 5472
rect 9858 5408 9874 5472
rect 9938 5408 9954 5472
rect 10018 5408 10024 5472
rect 9708 5407 10024 5408
rect 12629 5472 12945 5473
rect 12629 5408 12635 5472
rect 12699 5408 12715 5472
rect 12779 5408 12795 5472
rect 12859 5408 12875 5472
rect 12939 5408 12945 5472
rect 12629 5407 12945 5408
rect 2406 4928 2722 4929
rect 2406 4864 2412 4928
rect 2476 4864 2492 4928
rect 2556 4864 2572 4928
rect 2636 4864 2652 4928
rect 2716 4864 2722 4928
rect 2406 4863 2722 4864
rect 5327 4928 5643 4929
rect 5327 4864 5333 4928
rect 5397 4864 5413 4928
rect 5477 4864 5493 4928
rect 5557 4864 5573 4928
rect 5637 4864 5643 4928
rect 5327 4863 5643 4864
rect 8248 4928 8564 4929
rect 8248 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8494 4928
rect 8558 4864 8564 4928
rect 8248 4863 8564 4864
rect 11169 4928 11485 4929
rect 11169 4864 11175 4928
rect 11239 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11485 4928
rect 11169 4863 11485 4864
rect 0 4632 400 4752
rect 3866 4384 4182 4385
rect 3866 4320 3872 4384
rect 3936 4320 3952 4384
rect 4016 4320 4032 4384
rect 4096 4320 4112 4384
rect 4176 4320 4182 4384
rect 3866 4319 4182 4320
rect 6787 4384 7103 4385
rect 6787 4320 6793 4384
rect 6857 4320 6873 4384
rect 6937 4320 6953 4384
rect 7017 4320 7033 4384
rect 7097 4320 7103 4384
rect 6787 4319 7103 4320
rect 9708 4384 10024 4385
rect 9708 4320 9714 4384
rect 9778 4320 9794 4384
rect 9858 4320 9874 4384
rect 9938 4320 9954 4384
rect 10018 4320 10024 4384
rect 9708 4319 10024 4320
rect 12629 4384 12945 4385
rect 12629 4320 12635 4384
rect 12699 4320 12715 4384
rect 12779 4320 12795 4384
rect 12859 4320 12875 4384
rect 12939 4320 12945 4384
rect 12629 4319 12945 4320
rect 3693 4178 3759 4181
rect 5165 4178 5231 4181
rect 3693 4176 5231 4178
rect 3693 4120 3698 4176
rect 3754 4120 5170 4176
rect 5226 4120 5231 4176
rect 3693 4118 5231 4120
rect 3693 4115 3759 4118
rect 5165 4115 5231 4118
rect 0 3816 400 3936
rect 2406 3840 2722 3841
rect 2406 3776 2412 3840
rect 2476 3776 2492 3840
rect 2556 3776 2572 3840
rect 2636 3776 2652 3840
rect 2716 3776 2722 3840
rect 2406 3775 2722 3776
rect 5327 3840 5643 3841
rect 5327 3776 5333 3840
rect 5397 3776 5413 3840
rect 5477 3776 5493 3840
rect 5557 3776 5573 3840
rect 5637 3776 5643 3840
rect 5327 3775 5643 3776
rect 8248 3840 8564 3841
rect 8248 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8494 3840
rect 8558 3776 8564 3840
rect 8248 3775 8564 3776
rect 11169 3840 11485 3841
rect 11169 3776 11175 3840
rect 11239 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11485 3840
rect 11169 3775 11485 3776
rect 3866 3296 4182 3297
rect 3866 3232 3872 3296
rect 3936 3232 3952 3296
rect 4016 3232 4032 3296
rect 4096 3232 4112 3296
rect 4176 3232 4182 3296
rect 3866 3231 4182 3232
rect 6787 3296 7103 3297
rect 6787 3232 6793 3296
rect 6857 3232 6873 3296
rect 6937 3232 6953 3296
rect 7017 3232 7033 3296
rect 7097 3232 7103 3296
rect 6787 3231 7103 3232
rect 9708 3296 10024 3297
rect 9708 3232 9714 3296
rect 9778 3232 9794 3296
rect 9858 3232 9874 3296
rect 9938 3232 9954 3296
rect 10018 3232 10024 3296
rect 9708 3231 10024 3232
rect 12629 3296 12945 3297
rect 12629 3232 12635 3296
rect 12699 3232 12715 3296
rect 12779 3232 12795 3296
rect 12859 3232 12875 3296
rect 12939 3232 12945 3296
rect 12629 3231 12945 3232
rect 0 3000 400 3120
rect 2406 2752 2722 2753
rect 2406 2688 2412 2752
rect 2476 2688 2492 2752
rect 2556 2688 2572 2752
rect 2636 2688 2652 2752
rect 2716 2688 2722 2752
rect 2406 2687 2722 2688
rect 5327 2752 5643 2753
rect 5327 2688 5333 2752
rect 5397 2688 5413 2752
rect 5477 2688 5493 2752
rect 5557 2688 5573 2752
rect 5637 2688 5643 2752
rect 5327 2687 5643 2688
rect 8248 2752 8564 2753
rect 8248 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8494 2752
rect 8558 2688 8564 2752
rect 8248 2687 8564 2688
rect 11169 2752 11485 2753
rect 11169 2688 11175 2752
rect 11239 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11485 2752
rect 11169 2687 11485 2688
rect 0 2184 400 2304
rect 3866 2208 4182 2209
rect 3866 2144 3872 2208
rect 3936 2144 3952 2208
rect 4016 2144 4032 2208
rect 4096 2144 4112 2208
rect 4176 2144 4182 2208
rect 3866 2143 4182 2144
rect 6787 2208 7103 2209
rect 6787 2144 6793 2208
rect 6857 2144 6873 2208
rect 6937 2144 6953 2208
rect 7017 2144 7033 2208
rect 7097 2144 7103 2208
rect 6787 2143 7103 2144
rect 9708 2208 10024 2209
rect 9708 2144 9714 2208
rect 9778 2144 9794 2208
rect 9858 2144 9874 2208
rect 9938 2144 9954 2208
rect 10018 2144 10024 2208
rect 9708 2143 10024 2144
rect 12629 2208 12945 2209
rect 12629 2144 12635 2208
rect 12699 2144 12715 2208
rect 12779 2144 12795 2208
rect 12859 2144 12875 2208
rect 12939 2144 12945 2208
rect 12629 2143 12945 2144
rect 2406 1664 2722 1665
rect 2406 1600 2412 1664
rect 2476 1600 2492 1664
rect 2556 1600 2572 1664
rect 2636 1600 2652 1664
rect 2716 1600 2722 1664
rect 2406 1599 2722 1600
rect 5327 1664 5643 1665
rect 5327 1600 5333 1664
rect 5397 1600 5413 1664
rect 5477 1600 5493 1664
rect 5557 1600 5573 1664
rect 5637 1600 5643 1664
rect 5327 1599 5643 1600
rect 8248 1664 8564 1665
rect 8248 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8494 1664
rect 8558 1600 8564 1664
rect 8248 1599 8564 1600
rect 11169 1664 11485 1665
rect 11169 1600 11175 1664
rect 11239 1600 11255 1664
rect 11319 1600 11335 1664
rect 11399 1600 11415 1664
rect 11479 1600 11485 1664
rect 11169 1599 11485 1600
rect 0 1458 400 1488
rect 749 1458 815 1461
rect 0 1456 815 1458
rect 0 1400 754 1456
rect 810 1400 815 1456
rect 0 1398 815 1400
rect 0 1368 400 1398
rect 749 1395 815 1398
rect 3866 1120 4182 1121
rect 3866 1056 3872 1120
rect 3936 1056 3952 1120
rect 4016 1056 4032 1120
rect 4096 1056 4112 1120
rect 4176 1056 4182 1120
rect 3866 1055 4182 1056
rect 6787 1120 7103 1121
rect 6787 1056 6793 1120
rect 6857 1056 6873 1120
rect 6937 1056 6953 1120
rect 7017 1056 7033 1120
rect 7097 1056 7103 1120
rect 6787 1055 7103 1056
rect 9708 1120 10024 1121
rect 9708 1056 9714 1120
rect 9778 1056 9794 1120
rect 9858 1056 9874 1120
rect 9938 1056 9954 1120
rect 10018 1056 10024 1120
rect 9708 1055 10024 1056
rect 12629 1120 12945 1121
rect 12629 1056 12635 1120
rect 12699 1056 12715 1120
rect 12779 1056 12795 1120
rect 12859 1056 12875 1120
rect 12939 1056 12945 1120
rect 12629 1055 12945 1056
rect 0 642 400 672
rect 3785 642 3851 645
rect 0 640 3851 642
rect 0 584 3790 640
rect 3846 584 3851 640
rect 0 582 3851 584
rect 0 552 400 582
rect 3785 579 3851 582
<< via3 >>
rect 2412 12540 2476 12544
rect 2412 12484 2416 12540
rect 2416 12484 2472 12540
rect 2472 12484 2476 12540
rect 2412 12480 2476 12484
rect 2492 12540 2556 12544
rect 2492 12484 2496 12540
rect 2496 12484 2552 12540
rect 2552 12484 2556 12540
rect 2492 12480 2556 12484
rect 2572 12540 2636 12544
rect 2572 12484 2576 12540
rect 2576 12484 2632 12540
rect 2632 12484 2636 12540
rect 2572 12480 2636 12484
rect 2652 12540 2716 12544
rect 2652 12484 2656 12540
rect 2656 12484 2712 12540
rect 2712 12484 2716 12540
rect 2652 12480 2716 12484
rect 5333 12540 5397 12544
rect 5333 12484 5337 12540
rect 5337 12484 5393 12540
rect 5393 12484 5397 12540
rect 5333 12480 5397 12484
rect 5413 12540 5477 12544
rect 5413 12484 5417 12540
rect 5417 12484 5473 12540
rect 5473 12484 5477 12540
rect 5413 12480 5477 12484
rect 5493 12540 5557 12544
rect 5493 12484 5497 12540
rect 5497 12484 5553 12540
rect 5553 12484 5557 12540
rect 5493 12480 5557 12484
rect 5573 12540 5637 12544
rect 5573 12484 5577 12540
rect 5577 12484 5633 12540
rect 5633 12484 5637 12540
rect 5573 12480 5637 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 8494 12540 8558 12544
rect 8494 12484 8498 12540
rect 8498 12484 8554 12540
rect 8554 12484 8558 12540
rect 8494 12480 8558 12484
rect 11175 12540 11239 12544
rect 11175 12484 11179 12540
rect 11179 12484 11235 12540
rect 11235 12484 11239 12540
rect 11175 12480 11239 12484
rect 11255 12540 11319 12544
rect 11255 12484 11259 12540
rect 11259 12484 11315 12540
rect 11315 12484 11319 12540
rect 11255 12480 11319 12484
rect 11335 12540 11399 12544
rect 11335 12484 11339 12540
rect 11339 12484 11395 12540
rect 11395 12484 11399 12540
rect 11335 12480 11399 12484
rect 11415 12540 11479 12544
rect 11415 12484 11419 12540
rect 11419 12484 11475 12540
rect 11475 12484 11479 12540
rect 11415 12480 11479 12484
rect 3872 11996 3936 12000
rect 3872 11940 3876 11996
rect 3876 11940 3932 11996
rect 3932 11940 3936 11996
rect 3872 11936 3936 11940
rect 3952 11996 4016 12000
rect 3952 11940 3956 11996
rect 3956 11940 4012 11996
rect 4012 11940 4016 11996
rect 3952 11936 4016 11940
rect 4032 11996 4096 12000
rect 4032 11940 4036 11996
rect 4036 11940 4092 11996
rect 4092 11940 4096 11996
rect 4032 11936 4096 11940
rect 4112 11996 4176 12000
rect 4112 11940 4116 11996
rect 4116 11940 4172 11996
rect 4172 11940 4176 11996
rect 4112 11936 4176 11940
rect 6793 11996 6857 12000
rect 6793 11940 6797 11996
rect 6797 11940 6853 11996
rect 6853 11940 6857 11996
rect 6793 11936 6857 11940
rect 6873 11996 6937 12000
rect 6873 11940 6877 11996
rect 6877 11940 6933 11996
rect 6933 11940 6937 11996
rect 6873 11936 6937 11940
rect 6953 11996 7017 12000
rect 6953 11940 6957 11996
rect 6957 11940 7013 11996
rect 7013 11940 7017 11996
rect 6953 11936 7017 11940
rect 7033 11996 7097 12000
rect 7033 11940 7037 11996
rect 7037 11940 7093 11996
rect 7093 11940 7097 11996
rect 7033 11936 7097 11940
rect 9714 11996 9778 12000
rect 9714 11940 9718 11996
rect 9718 11940 9774 11996
rect 9774 11940 9778 11996
rect 9714 11936 9778 11940
rect 9794 11996 9858 12000
rect 9794 11940 9798 11996
rect 9798 11940 9854 11996
rect 9854 11940 9858 11996
rect 9794 11936 9858 11940
rect 9874 11996 9938 12000
rect 9874 11940 9878 11996
rect 9878 11940 9934 11996
rect 9934 11940 9938 11996
rect 9874 11936 9938 11940
rect 9954 11996 10018 12000
rect 9954 11940 9958 11996
rect 9958 11940 10014 11996
rect 10014 11940 10018 11996
rect 9954 11936 10018 11940
rect 12635 11996 12699 12000
rect 12635 11940 12639 11996
rect 12639 11940 12695 11996
rect 12695 11940 12699 11996
rect 12635 11936 12699 11940
rect 12715 11996 12779 12000
rect 12715 11940 12719 11996
rect 12719 11940 12775 11996
rect 12775 11940 12779 11996
rect 12715 11936 12779 11940
rect 12795 11996 12859 12000
rect 12795 11940 12799 11996
rect 12799 11940 12855 11996
rect 12855 11940 12859 11996
rect 12795 11936 12859 11940
rect 12875 11996 12939 12000
rect 12875 11940 12879 11996
rect 12879 11940 12935 11996
rect 12935 11940 12939 11996
rect 12875 11936 12939 11940
rect 2412 11452 2476 11456
rect 2412 11396 2416 11452
rect 2416 11396 2472 11452
rect 2472 11396 2476 11452
rect 2412 11392 2476 11396
rect 2492 11452 2556 11456
rect 2492 11396 2496 11452
rect 2496 11396 2552 11452
rect 2552 11396 2556 11452
rect 2492 11392 2556 11396
rect 2572 11452 2636 11456
rect 2572 11396 2576 11452
rect 2576 11396 2632 11452
rect 2632 11396 2636 11452
rect 2572 11392 2636 11396
rect 2652 11452 2716 11456
rect 2652 11396 2656 11452
rect 2656 11396 2712 11452
rect 2712 11396 2716 11452
rect 2652 11392 2716 11396
rect 5333 11452 5397 11456
rect 5333 11396 5337 11452
rect 5337 11396 5393 11452
rect 5393 11396 5397 11452
rect 5333 11392 5397 11396
rect 5413 11452 5477 11456
rect 5413 11396 5417 11452
rect 5417 11396 5473 11452
rect 5473 11396 5477 11452
rect 5413 11392 5477 11396
rect 5493 11452 5557 11456
rect 5493 11396 5497 11452
rect 5497 11396 5553 11452
rect 5553 11396 5557 11452
rect 5493 11392 5557 11396
rect 5573 11452 5637 11456
rect 5573 11396 5577 11452
rect 5577 11396 5633 11452
rect 5633 11396 5637 11452
rect 5573 11392 5637 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 8494 11452 8558 11456
rect 8494 11396 8498 11452
rect 8498 11396 8554 11452
rect 8554 11396 8558 11452
rect 8494 11392 8558 11396
rect 11175 11452 11239 11456
rect 11175 11396 11179 11452
rect 11179 11396 11235 11452
rect 11235 11396 11239 11452
rect 11175 11392 11239 11396
rect 11255 11452 11319 11456
rect 11255 11396 11259 11452
rect 11259 11396 11315 11452
rect 11315 11396 11319 11452
rect 11255 11392 11319 11396
rect 11335 11452 11399 11456
rect 11335 11396 11339 11452
rect 11339 11396 11395 11452
rect 11395 11396 11399 11452
rect 11335 11392 11399 11396
rect 11415 11452 11479 11456
rect 11415 11396 11419 11452
rect 11419 11396 11475 11452
rect 11475 11396 11479 11452
rect 11415 11392 11479 11396
rect 3872 10908 3936 10912
rect 3872 10852 3876 10908
rect 3876 10852 3932 10908
rect 3932 10852 3936 10908
rect 3872 10848 3936 10852
rect 3952 10908 4016 10912
rect 3952 10852 3956 10908
rect 3956 10852 4012 10908
rect 4012 10852 4016 10908
rect 3952 10848 4016 10852
rect 4032 10908 4096 10912
rect 4032 10852 4036 10908
rect 4036 10852 4092 10908
rect 4092 10852 4096 10908
rect 4032 10848 4096 10852
rect 4112 10908 4176 10912
rect 4112 10852 4116 10908
rect 4116 10852 4172 10908
rect 4172 10852 4176 10908
rect 4112 10848 4176 10852
rect 6793 10908 6857 10912
rect 6793 10852 6797 10908
rect 6797 10852 6853 10908
rect 6853 10852 6857 10908
rect 6793 10848 6857 10852
rect 6873 10908 6937 10912
rect 6873 10852 6877 10908
rect 6877 10852 6933 10908
rect 6933 10852 6937 10908
rect 6873 10848 6937 10852
rect 6953 10908 7017 10912
rect 6953 10852 6957 10908
rect 6957 10852 7013 10908
rect 7013 10852 7017 10908
rect 6953 10848 7017 10852
rect 7033 10908 7097 10912
rect 7033 10852 7037 10908
rect 7037 10852 7093 10908
rect 7093 10852 7097 10908
rect 7033 10848 7097 10852
rect 9714 10908 9778 10912
rect 9714 10852 9718 10908
rect 9718 10852 9774 10908
rect 9774 10852 9778 10908
rect 9714 10848 9778 10852
rect 9794 10908 9858 10912
rect 9794 10852 9798 10908
rect 9798 10852 9854 10908
rect 9854 10852 9858 10908
rect 9794 10848 9858 10852
rect 9874 10908 9938 10912
rect 9874 10852 9878 10908
rect 9878 10852 9934 10908
rect 9934 10852 9938 10908
rect 9874 10848 9938 10852
rect 9954 10908 10018 10912
rect 9954 10852 9958 10908
rect 9958 10852 10014 10908
rect 10014 10852 10018 10908
rect 9954 10848 10018 10852
rect 12635 10908 12699 10912
rect 12635 10852 12639 10908
rect 12639 10852 12695 10908
rect 12695 10852 12699 10908
rect 12635 10848 12699 10852
rect 12715 10908 12779 10912
rect 12715 10852 12719 10908
rect 12719 10852 12775 10908
rect 12775 10852 12779 10908
rect 12715 10848 12779 10852
rect 12795 10908 12859 10912
rect 12795 10852 12799 10908
rect 12799 10852 12855 10908
rect 12855 10852 12859 10908
rect 12795 10848 12859 10852
rect 12875 10908 12939 10912
rect 12875 10852 12879 10908
rect 12879 10852 12935 10908
rect 12935 10852 12939 10908
rect 12875 10848 12939 10852
rect 2412 10364 2476 10368
rect 2412 10308 2416 10364
rect 2416 10308 2472 10364
rect 2472 10308 2476 10364
rect 2412 10304 2476 10308
rect 2492 10364 2556 10368
rect 2492 10308 2496 10364
rect 2496 10308 2552 10364
rect 2552 10308 2556 10364
rect 2492 10304 2556 10308
rect 2572 10364 2636 10368
rect 2572 10308 2576 10364
rect 2576 10308 2632 10364
rect 2632 10308 2636 10364
rect 2572 10304 2636 10308
rect 2652 10364 2716 10368
rect 2652 10308 2656 10364
rect 2656 10308 2712 10364
rect 2712 10308 2716 10364
rect 2652 10304 2716 10308
rect 5333 10364 5397 10368
rect 5333 10308 5337 10364
rect 5337 10308 5393 10364
rect 5393 10308 5397 10364
rect 5333 10304 5397 10308
rect 5413 10364 5477 10368
rect 5413 10308 5417 10364
rect 5417 10308 5473 10364
rect 5473 10308 5477 10364
rect 5413 10304 5477 10308
rect 5493 10364 5557 10368
rect 5493 10308 5497 10364
rect 5497 10308 5553 10364
rect 5553 10308 5557 10364
rect 5493 10304 5557 10308
rect 5573 10364 5637 10368
rect 5573 10308 5577 10364
rect 5577 10308 5633 10364
rect 5633 10308 5637 10364
rect 5573 10304 5637 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 8494 10364 8558 10368
rect 8494 10308 8498 10364
rect 8498 10308 8554 10364
rect 8554 10308 8558 10364
rect 8494 10304 8558 10308
rect 11175 10364 11239 10368
rect 11175 10308 11179 10364
rect 11179 10308 11235 10364
rect 11235 10308 11239 10364
rect 11175 10304 11239 10308
rect 11255 10364 11319 10368
rect 11255 10308 11259 10364
rect 11259 10308 11315 10364
rect 11315 10308 11319 10364
rect 11255 10304 11319 10308
rect 11335 10364 11399 10368
rect 11335 10308 11339 10364
rect 11339 10308 11395 10364
rect 11395 10308 11399 10364
rect 11335 10304 11399 10308
rect 11415 10364 11479 10368
rect 11415 10308 11419 10364
rect 11419 10308 11475 10364
rect 11475 10308 11479 10364
rect 11415 10304 11479 10308
rect 3872 9820 3936 9824
rect 3872 9764 3876 9820
rect 3876 9764 3932 9820
rect 3932 9764 3936 9820
rect 3872 9760 3936 9764
rect 3952 9820 4016 9824
rect 3952 9764 3956 9820
rect 3956 9764 4012 9820
rect 4012 9764 4016 9820
rect 3952 9760 4016 9764
rect 4032 9820 4096 9824
rect 4032 9764 4036 9820
rect 4036 9764 4092 9820
rect 4092 9764 4096 9820
rect 4032 9760 4096 9764
rect 4112 9820 4176 9824
rect 4112 9764 4116 9820
rect 4116 9764 4172 9820
rect 4172 9764 4176 9820
rect 4112 9760 4176 9764
rect 6793 9820 6857 9824
rect 6793 9764 6797 9820
rect 6797 9764 6853 9820
rect 6853 9764 6857 9820
rect 6793 9760 6857 9764
rect 6873 9820 6937 9824
rect 6873 9764 6877 9820
rect 6877 9764 6933 9820
rect 6933 9764 6937 9820
rect 6873 9760 6937 9764
rect 6953 9820 7017 9824
rect 6953 9764 6957 9820
rect 6957 9764 7013 9820
rect 7013 9764 7017 9820
rect 6953 9760 7017 9764
rect 7033 9820 7097 9824
rect 7033 9764 7037 9820
rect 7037 9764 7093 9820
rect 7093 9764 7097 9820
rect 7033 9760 7097 9764
rect 9714 9820 9778 9824
rect 9714 9764 9718 9820
rect 9718 9764 9774 9820
rect 9774 9764 9778 9820
rect 9714 9760 9778 9764
rect 9794 9820 9858 9824
rect 9794 9764 9798 9820
rect 9798 9764 9854 9820
rect 9854 9764 9858 9820
rect 9794 9760 9858 9764
rect 9874 9820 9938 9824
rect 9874 9764 9878 9820
rect 9878 9764 9934 9820
rect 9934 9764 9938 9820
rect 9874 9760 9938 9764
rect 9954 9820 10018 9824
rect 9954 9764 9958 9820
rect 9958 9764 10014 9820
rect 10014 9764 10018 9820
rect 9954 9760 10018 9764
rect 12635 9820 12699 9824
rect 12635 9764 12639 9820
rect 12639 9764 12695 9820
rect 12695 9764 12699 9820
rect 12635 9760 12699 9764
rect 12715 9820 12779 9824
rect 12715 9764 12719 9820
rect 12719 9764 12775 9820
rect 12775 9764 12779 9820
rect 12715 9760 12779 9764
rect 12795 9820 12859 9824
rect 12795 9764 12799 9820
rect 12799 9764 12855 9820
rect 12855 9764 12859 9820
rect 12795 9760 12859 9764
rect 12875 9820 12939 9824
rect 12875 9764 12879 9820
rect 12879 9764 12935 9820
rect 12935 9764 12939 9820
rect 12875 9760 12939 9764
rect 2412 9276 2476 9280
rect 2412 9220 2416 9276
rect 2416 9220 2472 9276
rect 2472 9220 2476 9276
rect 2412 9216 2476 9220
rect 2492 9276 2556 9280
rect 2492 9220 2496 9276
rect 2496 9220 2552 9276
rect 2552 9220 2556 9276
rect 2492 9216 2556 9220
rect 2572 9276 2636 9280
rect 2572 9220 2576 9276
rect 2576 9220 2632 9276
rect 2632 9220 2636 9276
rect 2572 9216 2636 9220
rect 2652 9276 2716 9280
rect 2652 9220 2656 9276
rect 2656 9220 2712 9276
rect 2712 9220 2716 9276
rect 2652 9216 2716 9220
rect 5333 9276 5397 9280
rect 5333 9220 5337 9276
rect 5337 9220 5393 9276
rect 5393 9220 5397 9276
rect 5333 9216 5397 9220
rect 5413 9276 5477 9280
rect 5413 9220 5417 9276
rect 5417 9220 5473 9276
rect 5473 9220 5477 9276
rect 5413 9216 5477 9220
rect 5493 9276 5557 9280
rect 5493 9220 5497 9276
rect 5497 9220 5553 9276
rect 5553 9220 5557 9276
rect 5493 9216 5557 9220
rect 5573 9276 5637 9280
rect 5573 9220 5577 9276
rect 5577 9220 5633 9276
rect 5633 9220 5637 9276
rect 5573 9216 5637 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 8494 9276 8558 9280
rect 8494 9220 8498 9276
rect 8498 9220 8554 9276
rect 8554 9220 8558 9276
rect 8494 9216 8558 9220
rect 11175 9276 11239 9280
rect 11175 9220 11179 9276
rect 11179 9220 11235 9276
rect 11235 9220 11239 9276
rect 11175 9216 11239 9220
rect 11255 9276 11319 9280
rect 11255 9220 11259 9276
rect 11259 9220 11315 9276
rect 11315 9220 11319 9276
rect 11255 9216 11319 9220
rect 11335 9276 11399 9280
rect 11335 9220 11339 9276
rect 11339 9220 11395 9276
rect 11395 9220 11399 9276
rect 11335 9216 11399 9220
rect 11415 9276 11479 9280
rect 11415 9220 11419 9276
rect 11419 9220 11475 9276
rect 11475 9220 11479 9276
rect 11415 9216 11479 9220
rect 3872 8732 3936 8736
rect 3872 8676 3876 8732
rect 3876 8676 3932 8732
rect 3932 8676 3936 8732
rect 3872 8672 3936 8676
rect 3952 8732 4016 8736
rect 3952 8676 3956 8732
rect 3956 8676 4012 8732
rect 4012 8676 4016 8732
rect 3952 8672 4016 8676
rect 4032 8732 4096 8736
rect 4032 8676 4036 8732
rect 4036 8676 4092 8732
rect 4092 8676 4096 8732
rect 4032 8672 4096 8676
rect 4112 8732 4176 8736
rect 4112 8676 4116 8732
rect 4116 8676 4172 8732
rect 4172 8676 4176 8732
rect 4112 8672 4176 8676
rect 6793 8732 6857 8736
rect 6793 8676 6797 8732
rect 6797 8676 6853 8732
rect 6853 8676 6857 8732
rect 6793 8672 6857 8676
rect 6873 8732 6937 8736
rect 6873 8676 6877 8732
rect 6877 8676 6933 8732
rect 6933 8676 6937 8732
rect 6873 8672 6937 8676
rect 6953 8732 7017 8736
rect 6953 8676 6957 8732
rect 6957 8676 7013 8732
rect 7013 8676 7017 8732
rect 6953 8672 7017 8676
rect 7033 8732 7097 8736
rect 7033 8676 7037 8732
rect 7037 8676 7093 8732
rect 7093 8676 7097 8732
rect 7033 8672 7097 8676
rect 9714 8732 9778 8736
rect 9714 8676 9718 8732
rect 9718 8676 9774 8732
rect 9774 8676 9778 8732
rect 9714 8672 9778 8676
rect 9794 8732 9858 8736
rect 9794 8676 9798 8732
rect 9798 8676 9854 8732
rect 9854 8676 9858 8732
rect 9794 8672 9858 8676
rect 9874 8732 9938 8736
rect 9874 8676 9878 8732
rect 9878 8676 9934 8732
rect 9934 8676 9938 8732
rect 9874 8672 9938 8676
rect 9954 8732 10018 8736
rect 9954 8676 9958 8732
rect 9958 8676 10014 8732
rect 10014 8676 10018 8732
rect 9954 8672 10018 8676
rect 12635 8732 12699 8736
rect 12635 8676 12639 8732
rect 12639 8676 12695 8732
rect 12695 8676 12699 8732
rect 12635 8672 12699 8676
rect 12715 8732 12779 8736
rect 12715 8676 12719 8732
rect 12719 8676 12775 8732
rect 12775 8676 12779 8732
rect 12715 8672 12779 8676
rect 12795 8732 12859 8736
rect 12795 8676 12799 8732
rect 12799 8676 12855 8732
rect 12855 8676 12859 8732
rect 12795 8672 12859 8676
rect 12875 8732 12939 8736
rect 12875 8676 12879 8732
rect 12879 8676 12935 8732
rect 12935 8676 12939 8732
rect 12875 8672 12939 8676
rect 2412 8188 2476 8192
rect 2412 8132 2416 8188
rect 2416 8132 2472 8188
rect 2472 8132 2476 8188
rect 2412 8128 2476 8132
rect 2492 8188 2556 8192
rect 2492 8132 2496 8188
rect 2496 8132 2552 8188
rect 2552 8132 2556 8188
rect 2492 8128 2556 8132
rect 2572 8188 2636 8192
rect 2572 8132 2576 8188
rect 2576 8132 2632 8188
rect 2632 8132 2636 8188
rect 2572 8128 2636 8132
rect 2652 8188 2716 8192
rect 2652 8132 2656 8188
rect 2656 8132 2712 8188
rect 2712 8132 2716 8188
rect 2652 8128 2716 8132
rect 5333 8188 5397 8192
rect 5333 8132 5337 8188
rect 5337 8132 5393 8188
rect 5393 8132 5397 8188
rect 5333 8128 5397 8132
rect 5413 8188 5477 8192
rect 5413 8132 5417 8188
rect 5417 8132 5473 8188
rect 5473 8132 5477 8188
rect 5413 8128 5477 8132
rect 5493 8188 5557 8192
rect 5493 8132 5497 8188
rect 5497 8132 5553 8188
rect 5553 8132 5557 8188
rect 5493 8128 5557 8132
rect 5573 8188 5637 8192
rect 5573 8132 5577 8188
rect 5577 8132 5633 8188
rect 5633 8132 5637 8188
rect 5573 8128 5637 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 8494 8188 8558 8192
rect 8494 8132 8498 8188
rect 8498 8132 8554 8188
rect 8554 8132 8558 8188
rect 8494 8128 8558 8132
rect 11175 8188 11239 8192
rect 11175 8132 11179 8188
rect 11179 8132 11235 8188
rect 11235 8132 11239 8188
rect 11175 8128 11239 8132
rect 11255 8188 11319 8192
rect 11255 8132 11259 8188
rect 11259 8132 11315 8188
rect 11315 8132 11319 8188
rect 11255 8128 11319 8132
rect 11335 8188 11399 8192
rect 11335 8132 11339 8188
rect 11339 8132 11395 8188
rect 11395 8132 11399 8188
rect 11335 8128 11399 8132
rect 11415 8188 11479 8192
rect 11415 8132 11419 8188
rect 11419 8132 11475 8188
rect 11475 8132 11479 8188
rect 11415 8128 11479 8132
rect 3872 7644 3936 7648
rect 3872 7588 3876 7644
rect 3876 7588 3932 7644
rect 3932 7588 3936 7644
rect 3872 7584 3936 7588
rect 3952 7644 4016 7648
rect 3952 7588 3956 7644
rect 3956 7588 4012 7644
rect 4012 7588 4016 7644
rect 3952 7584 4016 7588
rect 4032 7644 4096 7648
rect 4032 7588 4036 7644
rect 4036 7588 4092 7644
rect 4092 7588 4096 7644
rect 4032 7584 4096 7588
rect 4112 7644 4176 7648
rect 4112 7588 4116 7644
rect 4116 7588 4172 7644
rect 4172 7588 4176 7644
rect 4112 7584 4176 7588
rect 6793 7644 6857 7648
rect 6793 7588 6797 7644
rect 6797 7588 6853 7644
rect 6853 7588 6857 7644
rect 6793 7584 6857 7588
rect 6873 7644 6937 7648
rect 6873 7588 6877 7644
rect 6877 7588 6933 7644
rect 6933 7588 6937 7644
rect 6873 7584 6937 7588
rect 6953 7644 7017 7648
rect 6953 7588 6957 7644
rect 6957 7588 7013 7644
rect 7013 7588 7017 7644
rect 6953 7584 7017 7588
rect 7033 7644 7097 7648
rect 7033 7588 7037 7644
rect 7037 7588 7093 7644
rect 7093 7588 7097 7644
rect 7033 7584 7097 7588
rect 9714 7644 9778 7648
rect 9714 7588 9718 7644
rect 9718 7588 9774 7644
rect 9774 7588 9778 7644
rect 9714 7584 9778 7588
rect 9794 7644 9858 7648
rect 9794 7588 9798 7644
rect 9798 7588 9854 7644
rect 9854 7588 9858 7644
rect 9794 7584 9858 7588
rect 9874 7644 9938 7648
rect 9874 7588 9878 7644
rect 9878 7588 9934 7644
rect 9934 7588 9938 7644
rect 9874 7584 9938 7588
rect 9954 7644 10018 7648
rect 9954 7588 9958 7644
rect 9958 7588 10014 7644
rect 10014 7588 10018 7644
rect 9954 7584 10018 7588
rect 12635 7644 12699 7648
rect 12635 7588 12639 7644
rect 12639 7588 12695 7644
rect 12695 7588 12699 7644
rect 12635 7584 12699 7588
rect 12715 7644 12779 7648
rect 12715 7588 12719 7644
rect 12719 7588 12775 7644
rect 12775 7588 12779 7644
rect 12715 7584 12779 7588
rect 12795 7644 12859 7648
rect 12795 7588 12799 7644
rect 12799 7588 12855 7644
rect 12855 7588 12859 7644
rect 12795 7584 12859 7588
rect 12875 7644 12939 7648
rect 12875 7588 12879 7644
rect 12879 7588 12935 7644
rect 12935 7588 12939 7644
rect 12875 7584 12939 7588
rect 2412 7100 2476 7104
rect 2412 7044 2416 7100
rect 2416 7044 2472 7100
rect 2472 7044 2476 7100
rect 2412 7040 2476 7044
rect 2492 7100 2556 7104
rect 2492 7044 2496 7100
rect 2496 7044 2552 7100
rect 2552 7044 2556 7100
rect 2492 7040 2556 7044
rect 2572 7100 2636 7104
rect 2572 7044 2576 7100
rect 2576 7044 2632 7100
rect 2632 7044 2636 7100
rect 2572 7040 2636 7044
rect 2652 7100 2716 7104
rect 2652 7044 2656 7100
rect 2656 7044 2712 7100
rect 2712 7044 2716 7100
rect 2652 7040 2716 7044
rect 5333 7100 5397 7104
rect 5333 7044 5337 7100
rect 5337 7044 5393 7100
rect 5393 7044 5397 7100
rect 5333 7040 5397 7044
rect 5413 7100 5477 7104
rect 5413 7044 5417 7100
rect 5417 7044 5473 7100
rect 5473 7044 5477 7100
rect 5413 7040 5477 7044
rect 5493 7100 5557 7104
rect 5493 7044 5497 7100
rect 5497 7044 5553 7100
rect 5553 7044 5557 7100
rect 5493 7040 5557 7044
rect 5573 7100 5637 7104
rect 5573 7044 5577 7100
rect 5577 7044 5633 7100
rect 5633 7044 5637 7100
rect 5573 7040 5637 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 8494 7100 8558 7104
rect 8494 7044 8498 7100
rect 8498 7044 8554 7100
rect 8554 7044 8558 7100
rect 8494 7040 8558 7044
rect 11175 7100 11239 7104
rect 11175 7044 11179 7100
rect 11179 7044 11235 7100
rect 11235 7044 11239 7100
rect 11175 7040 11239 7044
rect 11255 7100 11319 7104
rect 11255 7044 11259 7100
rect 11259 7044 11315 7100
rect 11315 7044 11319 7100
rect 11255 7040 11319 7044
rect 11335 7100 11399 7104
rect 11335 7044 11339 7100
rect 11339 7044 11395 7100
rect 11395 7044 11399 7100
rect 11335 7040 11399 7044
rect 11415 7100 11479 7104
rect 11415 7044 11419 7100
rect 11419 7044 11475 7100
rect 11475 7044 11479 7100
rect 11415 7040 11479 7044
rect 3872 6556 3936 6560
rect 3872 6500 3876 6556
rect 3876 6500 3932 6556
rect 3932 6500 3936 6556
rect 3872 6496 3936 6500
rect 3952 6556 4016 6560
rect 3952 6500 3956 6556
rect 3956 6500 4012 6556
rect 4012 6500 4016 6556
rect 3952 6496 4016 6500
rect 4032 6556 4096 6560
rect 4032 6500 4036 6556
rect 4036 6500 4092 6556
rect 4092 6500 4096 6556
rect 4032 6496 4096 6500
rect 4112 6556 4176 6560
rect 4112 6500 4116 6556
rect 4116 6500 4172 6556
rect 4172 6500 4176 6556
rect 4112 6496 4176 6500
rect 6793 6556 6857 6560
rect 6793 6500 6797 6556
rect 6797 6500 6853 6556
rect 6853 6500 6857 6556
rect 6793 6496 6857 6500
rect 6873 6556 6937 6560
rect 6873 6500 6877 6556
rect 6877 6500 6933 6556
rect 6933 6500 6937 6556
rect 6873 6496 6937 6500
rect 6953 6556 7017 6560
rect 6953 6500 6957 6556
rect 6957 6500 7013 6556
rect 7013 6500 7017 6556
rect 6953 6496 7017 6500
rect 7033 6556 7097 6560
rect 7033 6500 7037 6556
rect 7037 6500 7093 6556
rect 7093 6500 7097 6556
rect 7033 6496 7097 6500
rect 9714 6556 9778 6560
rect 9714 6500 9718 6556
rect 9718 6500 9774 6556
rect 9774 6500 9778 6556
rect 9714 6496 9778 6500
rect 9794 6556 9858 6560
rect 9794 6500 9798 6556
rect 9798 6500 9854 6556
rect 9854 6500 9858 6556
rect 9794 6496 9858 6500
rect 9874 6556 9938 6560
rect 9874 6500 9878 6556
rect 9878 6500 9934 6556
rect 9934 6500 9938 6556
rect 9874 6496 9938 6500
rect 9954 6556 10018 6560
rect 9954 6500 9958 6556
rect 9958 6500 10014 6556
rect 10014 6500 10018 6556
rect 9954 6496 10018 6500
rect 12635 6556 12699 6560
rect 12635 6500 12639 6556
rect 12639 6500 12695 6556
rect 12695 6500 12699 6556
rect 12635 6496 12699 6500
rect 12715 6556 12779 6560
rect 12715 6500 12719 6556
rect 12719 6500 12775 6556
rect 12775 6500 12779 6556
rect 12715 6496 12779 6500
rect 12795 6556 12859 6560
rect 12795 6500 12799 6556
rect 12799 6500 12855 6556
rect 12855 6500 12859 6556
rect 12795 6496 12859 6500
rect 12875 6556 12939 6560
rect 12875 6500 12879 6556
rect 12879 6500 12935 6556
rect 12935 6500 12939 6556
rect 12875 6496 12939 6500
rect 2412 6012 2476 6016
rect 2412 5956 2416 6012
rect 2416 5956 2472 6012
rect 2472 5956 2476 6012
rect 2412 5952 2476 5956
rect 2492 6012 2556 6016
rect 2492 5956 2496 6012
rect 2496 5956 2552 6012
rect 2552 5956 2556 6012
rect 2492 5952 2556 5956
rect 2572 6012 2636 6016
rect 2572 5956 2576 6012
rect 2576 5956 2632 6012
rect 2632 5956 2636 6012
rect 2572 5952 2636 5956
rect 2652 6012 2716 6016
rect 2652 5956 2656 6012
rect 2656 5956 2712 6012
rect 2712 5956 2716 6012
rect 2652 5952 2716 5956
rect 5333 6012 5397 6016
rect 5333 5956 5337 6012
rect 5337 5956 5393 6012
rect 5393 5956 5397 6012
rect 5333 5952 5397 5956
rect 5413 6012 5477 6016
rect 5413 5956 5417 6012
rect 5417 5956 5473 6012
rect 5473 5956 5477 6012
rect 5413 5952 5477 5956
rect 5493 6012 5557 6016
rect 5493 5956 5497 6012
rect 5497 5956 5553 6012
rect 5553 5956 5557 6012
rect 5493 5952 5557 5956
rect 5573 6012 5637 6016
rect 5573 5956 5577 6012
rect 5577 5956 5633 6012
rect 5633 5956 5637 6012
rect 5573 5952 5637 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 8494 6012 8558 6016
rect 8494 5956 8498 6012
rect 8498 5956 8554 6012
rect 8554 5956 8558 6012
rect 8494 5952 8558 5956
rect 11175 6012 11239 6016
rect 11175 5956 11179 6012
rect 11179 5956 11235 6012
rect 11235 5956 11239 6012
rect 11175 5952 11239 5956
rect 11255 6012 11319 6016
rect 11255 5956 11259 6012
rect 11259 5956 11315 6012
rect 11315 5956 11319 6012
rect 11255 5952 11319 5956
rect 11335 6012 11399 6016
rect 11335 5956 11339 6012
rect 11339 5956 11395 6012
rect 11395 5956 11399 6012
rect 11335 5952 11399 5956
rect 11415 6012 11479 6016
rect 11415 5956 11419 6012
rect 11419 5956 11475 6012
rect 11475 5956 11479 6012
rect 11415 5952 11479 5956
rect 3872 5468 3936 5472
rect 3872 5412 3876 5468
rect 3876 5412 3932 5468
rect 3932 5412 3936 5468
rect 3872 5408 3936 5412
rect 3952 5468 4016 5472
rect 3952 5412 3956 5468
rect 3956 5412 4012 5468
rect 4012 5412 4016 5468
rect 3952 5408 4016 5412
rect 4032 5468 4096 5472
rect 4032 5412 4036 5468
rect 4036 5412 4092 5468
rect 4092 5412 4096 5468
rect 4032 5408 4096 5412
rect 4112 5468 4176 5472
rect 4112 5412 4116 5468
rect 4116 5412 4172 5468
rect 4172 5412 4176 5468
rect 4112 5408 4176 5412
rect 6793 5468 6857 5472
rect 6793 5412 6797 5468
rect 6797 5412 6853 5468
rect 6853 5412 6857 5468
rect 6793 5408 6857 5412
rect 6873 5468 6937 5472
rect 6873 5412 6877 5468
rect 6877 5412 6933 5468
rect 6933 5412 6937 5468
rect 6873 5408 6937 5412
rect 6953 5468 7017 5472
rect 6953 5412 6957 5468
rect 6957 5412 7013 5468
rect 7013 5412 7017 5468
rect 6953 5408 7017 5412
rect 7033 5468 7097 5472
rect 7033 5412 7037 5468
rect 7037 5412 7093 5468
rect 7093 5412 7097 5468
rect 7033 5408 7097 5412
rect 9714 5468 9778 5472
rect 9714 5412 9718 5468
rect 9718 5412 9774 5468
rect 9774 5412 9778 5468
rect 9714 5408 9778 5412
rect 9794 5468 9858 5472
rect 9794 5412 9798 5468
rect 9798 5412 9854 5468
rect 9854 5412 9858 5468
rect 9794 5408 9858 5412
rect 9874 5468 9938 5472
rect 9874 5412 9878 5468
rect 9878 5412 9934 5468
rect 9934 5412 9938 5468
rect 9874 5408 9938 5412
rect 9954 5468 10018 5472
rect 9954 5412 9958 5468
rect 9958 5412 10014 5468
rect 10014 5412 10018 5468
rect 9954 5408 10018 5412
rect 12635 5468 12699 5472
rect 12635 5412 12639 5468
rect 12639 5412 12695 5468
rect 12695 5412 12699 5468
rect 12635 5408 12699 5412
rect 12715 5468 12779 5472
rect 12715 5412 12719 5468
rect 12719 5412 12775 5468
rect 12775 5412 12779 5468
rect 12715 5408 12779 5412
rect 12795 5468 12859 5472
rect 12795 5412 12799 5468
rect 12799 5412 12855 5468
rect 12855 5412 12859 5468
rect 12795 5408 12859 5412
rect 12875 5468 12939 5472
rect 12875 5412 12879 5468
rect 12879 5412 12935 5468
rect 12935 5412 12939 5468
rect 12875 5408 12939 5412
rect 2412 4924 2476 4928
rect 2412 4868 2416 4924
rect 2416 4868 2472 4924
rect 2472 4868 2476 4924
rect 2412 4864 2476 4868
rect 2492 4924 2556 4928
rect 2492 4868 2496 4924
rect 2496 4868 2552 4924
rect 2552 4868 2556 4924
rect 2492 4864 2556 4868
rect 2572 4924 2636 4928
rect 2572 4868 2576 4924
rect 2576 4868 2632 4924
rect 2632 4868 2636 4924
rect 2572 4864 2636 4868
rect 2652 4924 2716 4928
rect 2652 4868 2656 4924
rect 2656 4868 2712 4924
rect 2712 4868 2716 4924
rect 2652 4864 2716 4868
rect 5333 4924 5397 4928
rect 5333 4868 5337 4924
rect 5337 4868 5393 4924
rect 5393 4868 5397 4924
rect 5333 4864 5397 4868
rect 5413 4924 5477 4928
rect 5413 4868 5417 4924
rect 5417 4868 5473 4924
rect 5473 4868 5477 4924
rect 5413 4864 5477 4868
rect 5493 4924 5557 4928
rect 5493 4868 5497 4924
rect 5497 4868 5553 4924
rect 5553 4868 5557 4924
rect 5493 4864 5557 4868
rect 5573 4924 5637 4928
rect 5573 4868 5577 4924
rect 5577 4868 5633 4924
rect 5633 4868 5637 4924
rect 5573 4864 5637 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 8494 4924 8558 4928
rect 8494 4868 8498 4924
rect 8498 4868 8554 4924
rect 8554 4868 8558 4924
rect 8494 4864 8558 4868
rect 11175 4924 11239 4928
rect 11175 4868 11179 4924
rect 11179 4868 11235 4924
rect 11235 4868 11239 4924
rect 11175 4864 11239 4868
rect 11255 4924 11319 4928
rect 11255 4868 11259 4924
rect 11259 4868 11315 4924
rect 11315 4868 11319 4924
rect 11255 4864 11319 4868
rect 11335 4924 11399 4928
rect 11335 4868 11339 4924
rect 11339 4868 11395 4924
rect 11395 4868 11399 4924
rect 11335 4864 11399 4868
rect 11415 4924 11479 4928
rect 11415 4868 11419 4924
rect 11419 4868 11475 4924
rect 11475 4868 11479 4924
rect 11415 4864 11479 4868
rect 3872 4380 3936 4384
rect 3872 4324 3876 4380
rect 3876 4324 3932 4380
rect 3932 4324 3936 4380
rect 3872 4320 3936 4324
rect 3952 4380 4016 4384
rect 3952 4324 3956 4380
rect 3956 4324 4012 4380
rect 4012 4324 4016 4380
rect 3952 4320 4016 4324
rect 4032 4380 4096 4384
rect 4032 4324 4036 4380
rect 4036 4324 4092 4380
rect 4092 4324 4096 4380
rect 4032 4320 4096 4324
rect 4112 4380 4176 4384
rect 4112 4324 4116 4380
rect 4116 4324 4172 4380
rect 4172 4324 4176 4380
rect 4112 4320 4176 4324
rect 6793 4380 6857 4384
rect 6793 4324 6797 4380
rect 6797 4324 6853 4380
rect 6853 4324 6857 4380
rect 6793 4320 6857 4324
rect 6873 4380 6937 4384
rect 6873 4324 6877 4380
rect 6877 4324 6933 4380
rect 6933 4324 6937 4380
rect 6873 4320 6937 4324
rect 6953 4380 7017 4384
rect 6953 4324 6957 4380
rect 6957 4324 7013 4380
rect 7013 4324 7017 4380
rect 6953 4320 7017 4324
rect 7033 4380 7097 4384
rect 7033 4324 7037 4380
rect 7037 4324 7093 4380
rect 7093 4324 7097 4380
rect 7033 4320 7097 4324
rect 9714 4380 9778 4384
rect 9714 4324 9718 4380
rect 9718 4324 9774 4380
rect 9774 4324 9778 4380
rect 9714 4320 9778 4324
rect 9794 4380 9858 4384
rect 9794 4324 9798 4380
rect 9798 4324 9854 4380
rect 9854 4324 9858 4380
rect 9794 4320 9858 4324
rect 9874 4380 9938 4384
rect 9874 4324 9878 4380
rect 9878 4324 9934 4380
rect 9934 4324 9938 4380
rect 9874 4320 9938 4324
rect 9954 4380 10018 4384
rect 9954 4324 9958 4380
rect 9958 4324 10014 4380
rect 10014 4324 10018 4380
rect 9954 4320 10018 4324
rect 12635 4380 12699 4384
rect 12635 4324 12639 4380
rect 12639 4324 12695 4380
rect 12695 4324 12699 4380
rect 12635 4320 12699 4324
rect 12715 4380 12779 4384
rect 12715 4324 12719 4380
rect 12719 4324 12775 4380
rect 12775 4324 12779 4380
rect 12715 4320 12779 4324
rect 12795 4380 12859 4384
rect 12795 4324 12799 4380
rect 12799 4324 12855 4380
rect 12855 4324 12859 4380
rect 12795 4320 12859 4324
rect 12875 4380 12939 4384
rect 12875 4324 12879 4380
rect 12879 4324 12935 4380
rect 12935 4324 12939 4380
rect 12875 4320 12939 4324
rect 2412 3836 2476 3840
rect 2412 3780 2416 3836
rect 2416 3780 2472 3836
rect 2472 3780 2476 3836
rect 2412 3776 2476 3780
rect 2492 3836 2556 3840
rect 2492 3780 2496 3836
rect 2496 3780 2552 3836
rect 2552 3780 2556 3836
rect 2492 3776 2556 3780
rect 2572 3836 2636 3840
rect 2572 3780 2576 3836
rect 2576 3780 2632 3836
rect 2632 3780 2636 3836
rect 2572 3776 2636 3780
rect 2652 3836 2716 3840
rect 2652 3780 2656 3836
rect 2656 3780 2712 3836
rect 2712 3780 2716 3836
rect 2652 3776 2716 3780
rect 5333 3836 5397 3840
rect 5333 3780 5337 3836
rect 5337 3780 5393 3836
rect 5393 3780 5397 3836
rect 5333 3776 5397 3780
rect 5413 3836 5477 3840
rect 5413 3780 5417 3836
rect 5417 3780 5473 3836
rect 5473 3780 5477 3836
rect 5413 3776 5477 3780
rect 5493 3836 5557 3840
rect 5493 3780 5497 3836
rect 5497 3780 5553 3836
rect 5553 3780 5557 3836
rect 5493 3776 5557 3780
rect 5573 3836 5637 3840
rect 5573 3780 5577 3836
rect 5577 3780 5633 3836
rect 5633 3780 5637 3836
rect 5573 3776 5637 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 8494 3836 8558 3840
rect 8494 3780 8498 3836
rect 8498 3780 8554 3836
rect 8554 3780 8558 3836
rect 8494 3776 8558 3780
rect 11175 3836 11239 3840
rect 11175 3780 11179 3836
rect 11179 3780 11235 3836
rect 11235 3780 11239 3836
rect 11175 3776 11239 3780
rect 11255 3836 11319 3840
rect 11255 3780 11259 3836
rect 11259 3780 11315 3836
rect 11315 3780 11319 3836
rect 11255 3776 11319 3780
rect 11335 3836 11399 3840
rect 11335 3780 11339 3836
rect 11339 3780 11395 3836
rect 11395 3780 11399 3836
rect 11335 3776 11399 3780
rect 11415 3836 11479 3840
rect 11415 3780 11419 3836
rect 11419 3780 11475 3836
rect 11475 3780 11479 3836
rect 11415 3776 11479 3780
rect 3872 3292 3936 3296
rect 3872 3236 3876 3292
rect 3876 3236 3932 3292
rect 3932 3236 3936 3292
rect 3872 3232 3936 3236
rect 3952 3292 4016 3296
rect 3952 3236 3956 3292
rect 3956 3236 4012 3292
rect 4012 3236 4016 3292
rect 3952 3232 4016 3236
rect 4032 3292 4096 3296
rect 4032 3236 4036 3292
rect 4036 3236 4092 3292
rect 4092 3236 4096 3292
rect 4032 3232 4096 3236
rect 4112 3292 4176 3296
rect 4112 3236 4116 3292
rect 4116 3236 4172 3292
rect 4172 3236 4176 3292
rect 4112 3232 4176 3236
rect 6793 3292 6857 3296
rect 6793 3236 6797 3292
rect 6797 3236 6853 3292
rect 6853 3236 6857 3292
rect 6793 3232 6857 3236
rect 6873 3292 6937 3296
rect 6873 3236 6877 3292
rect 6877 3236 6933 3292
rect 6933 3236 6937 3292
rect 6873 3232 6937 3236
rect 6953 3292 7017 3296
rect 6953 3236 6957 3292
rect 6957 3236 7013 3292
rect 7013 3236 7017 3292
rect 6953 3232 7017 3236
rect 7033 3292 7097 3296
rect 7033 3236 7037 3292
rect 7037 3236 7093 3292
rect 7093 3236 7097 3292
rect 7033 3232 7097 3236
rect 9714 3292 9778 3296
rect 9714 3236 9718 3292
rect 9718 3236 9774 3292
rect 9774 3236 9778 3292
rect 9714 3232 9778 3236
rect 9794 3292 9858 3296
rect 9794 3236 9798 3292
rect 9798 3236 9854 3292
rect 9854 3236 9858 3292
rect 9794 3232 9858 3236
rect 9874 3292 9938 3296
rect 9874 3236 9878 3292
rect 9878 3236 9934 3292
rect 9934 3236 9938 3292
rect 9874 3232 9938 3236
rect 9954 3292 10018 3296
rect 9954 3236 9958 3292
rect 9958 3236 10014 3292
rect 10014 3236 10018 3292
rect 9954 3232 10018 3236
rect 12635 3292 12699 3296
rect 12635 3236 12639 3292
rect 12639 3236 12695 3292
rect 12695 3236 12699 3292
rect 12635 3232 12699 3236
rect 12715 3292 12779 3296
rect 12715 3236 12719 3292
rect 12719 3236 12775 3292
rect 12775 3236 12779 3292
rect 12715 3232 12779 3236
rect 12795 3292 12859 3296
rect 12795 3236 12799 3292
rect 12799 3236 12855 3292
rect 12855 3236 12859 3292
rect 12795 3232 12859 3236
rect 12875 3292 12939 3296
rect 12875 3236 12879 3292
rect 12879 3236 12935 3292
rect 12935 3236 12939 3292
rect 12875 3232 12939 3236
rect 2412 2748 2476 2752
rect 2412 2692 2416 2748
rect 2416 2692 2472 2748
rect 2472 2692 2476 2748
rect 2412 2688 2476 2692
rect 2492 2748 2556 2752
rect 2492 2692 2496 2748
rect 2496 2692 2552 2748
rect 2552 2692 2556 2748
rect 2492 2688 2556 2692
rect 2572 2748 2636 2752
rect 2572 2692 2576 2748
rect 2576 2692 2632 2748
rect 2632 2692 2636 2748
rect 2572 2688 2636 2692
rect 2652 2748 2716 2752
rect 2652 2692 2656 2748
rect 2656 2692 2712 2748
rect 2712 2692 2716 2748
rect 2652 2688 2716 2692
rect 5333 2748 5397 2752
rect 5333 2692 5337 2748
rect 5337 2692 5393 2748
rect 5393 2692 5397 2748
rect 5333 2688 5397 2692
rect 5413 2748 5477 2752
rect 5413 2692 5417 2748
rect 5417 2692 5473 2748
rect 5473 2692 5477 2748
rect 5413 2688 5477 2692
rect 5493 2748 5557 2752
rect 5493 2692 5497 2748
rect 5497 2692 5553 2748
rect 5553 2692 5557 2748
rect 5493 2688 5557 2692
rect 5573 2748 5637 2752
rect 5573 2692 5577 2748
rect 5577 2692 5633 2748
rect 5633 2692 5637 2748
rect 5573 2688 5637 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 8494 2748 8558 2752
rect 8494 2692 8498 2748
rect 8498 2692 8554 2748
rect 8554 2692 8558 2748
rect 8494 2688 8558 2692
rect 11175 2748 11239 2752
rect 11175 2692 11179 2748
rect 11179 2692 11235 2748
rect 11235 2692 11239 2748
rect 11175 2688 11239 2692
rect 11255 2748 11319 2752
rect 11255 2692 11259 2748
rect 11259 2692 11315 2748
rect 11315 2692 11319 2748
rect 11255 2688 11319 2692
rect 11335 2748 11399 2752
rect 11335 2692 11339 2748
rect 11339 2692 11395 2748
rect 11395 2692 11399 2748
rect 11335 2688 11399 2692
rect 11415 2748 11479 2752
rect 11415 2692 11419 2748
rect 11419 2692 11475 2748
rect 11475 2692 11479 2748
rect 11415 2688 11479 2692
rect 3872 2204 3936 2208
rect 3872 2148 3876 2204
rect 3876 2148 3932 2204
rect 3932 2148 3936 2204
rect 3872 2144 3936 2148
rect 3952 2204 4016 2208
rect 3952 2148 3956 2204
rect 3956 2148 4012 2204
rect 4012 2148 4016 2204
rect 3952 2144 4016 2148
rect 4032 2204 4096 2208
rect 4032 2148 4036 2204
rect 4036 2148 4092 2204
rect 4092 2148 4096 2204
rect 4032 2144 4096 2148
rect 4112 2204 4176 2208
rect 4112 2148 4116 2204
rect 4116 2148 4172 2204
rect 4172 2148 4176 2204
rect 4112 2144 4176 2148
rect 6793 2204 6857 2208
rect 6793 2148 6797 2204
rect 6797 2148 6853 2204
rect 6853 2148 6857 2204
rect 6793 2144 6857 2148
rect 6873 2204 6937 2208
rect 6873 2148 6877 2204
rect 6877 2148 6933 2204
rect 6933 2148 6937 2204
rect 6873 2144 6937 2148
rect 6953 2204 7017 2208
rect 6953 2148 6957 2204
rect 6957 2148 7013 2204
rect 7013 2148 7017 2204
rect 6953 2144 7017 2148
rect 7033 2204 7097 2208
rect 7033 2148 7037 2204
rect 7037 2148 7093 2204
rect 7093 2148 7097 2204
rect 7033 2144 7097 2148
rect 9714 2204 9778 2208
rect 9714 2148 9718 2204
rect 9718 2148 9774 2204
rect 9774 2148 9778 2204
rect 9714 2144 9778 2148
rect 9794 2204 9858 2208
rect 9794 2148 9798 2204
rect 9798 2148 9854 2204
rect 9854 2148 9858 2204
rect 9794 2144 9858 2148
rect 9874 2204 9938 2208
rect 9874 2148 9878 2204
rect 9878 2148 9934 2204
rect 9934 2148 9938 2204
rect 9874 2144 9938 2148
rect 9954 2204 10018 2208
rect 9954 2148 9958 2204
rect 9958 2148 10014 2204
rect 10014 2148 10018 2204
rect 9954 2144 10018 2148
rect 12635 2204 12699 2208
rect 12635 2148 12639 2204
rect 12639 2148 12695 2204
rect 12695 2148 12699 2204
rect 12635 2144 12699 2148
rect 12715 2204 12779 2208
rect 12715 2148 12719 2204
rect 12719 2148 12775 2204
rect 12775 2148 12779 2204
rect 12715 2144 12779 2148
rect 12795 2204 12859 2208
rect 12795 2148 12799 2204
rect 12799 2148 12855 2204
rect 12855 2148 12859 2204
rect 12795 2144 12859 2148
rect 12875 2204 12939 2208
rect 12875 2148 12879 2204
rect 12879 2148 12935 2204
rect 12935 2148 12939 2204
rect 12875 2144 12939 2148
rect 2412 1660 2476 1664
rect 2412 1604 2416 1660
rect 2416 1604 2472 1660
rect 2472 1604 2476 1660
rect 2412 1600 2476 1604
rect 2492 1660 2556 1664
rect 2492 1604 2496 1660
rect 2496 1604 2552 1660
rect 2552 1604 2556 1660
rect 2492 1600 2556 1604
rect 2572 1660 2636 1664
rect 2572 1604 2576 1660
rect 2576 1604 2632 1660
rect 2632 1604 2636 1660
rect 2572 1600 2636 1604
rect 2652 1660 2716 1664
rect 2652 1604 2656 1660
rect 2656 1604 2712 1660
rect 2712 1604 2716 1660
rect 2652 1600 2716 1604
rect 5333 1660 5397 1664
rect 5333 1604 5337 1660
rect 5337 1604 5393 1660
rect 5393 1604 5397 1660
rect 5333 1600 5397 1604
rect 5413 1660 5477 1664
rect 5413 1604 5417 1660
rect 5417 1604 5473 1660
rect 5473 1604 5477 1660
rect 5413 1600 5477 1604
rect 5493 1660 5557 1664
rect 5493 1604 5497 1660
rect 5497 1604 5553 1660
rect 5553 1604 5557 1660
rect 5493 1600 5557 1604
rect 5573 1660 5637 1664
rect 5573 1604 5577 1660
rect 5577 1604 5633 1660
rect 5633 1604 5637 1660
rect 5573 1600 5637 1604
rect 8254 1660 8318 1664
rect 8254 1604 8258 1660
rect 8258 1604 8314 1660
rect 8314 1604 8318 1660
rect 8254 1600 8318 1604
rect 8334 1660 8398 1664
rect 8334 1604 8338 1660
rect 8338 1604 8394 1660
rect 8394 1604 8398 1660
rect 8334 1600 8398 1604
rect 8414 1660 8478 1664
rect 8414 1604 8418 1660
rect 8418 1604 8474 1660
rect 8474 1604 8478 1660
rect 8414 1600 8478 1604
rect 8494 1660 8558 1664
rect 8494 1604 8498 1660
rect 8498 1604 8554 1660
rect 8554 1604 8558 1660
rect 8494 1600 8558 1604
rect 11175 1660 11239 1664
rect 11175 1604 11179 1660
rect 11179 1604 11235 1660
rect 11235 1604 11239 1660
rect 11175 1600 11239 1604
rect 11255 1660 11319 1664
rect 11255 1604 11259 1660
rect 11259 1604 11315 1660
rect 11315 1604 11319 1660
rect 11255 1600 11319 1604
rect 11335 1660 11399 1664
rect 11335 1604 11339 1660
rect 11339 1604 11395 1660
rect 11395 1604 11399 1660
rect 11335 1600 11399 1604
rect 11415 1660 11479 1664
rect 11415 1604 11419 1660
rect 11419 1604 11475 1660
rect 11475 1604 11479 1660
rect 11415 1600 11479 1604
rect 3872 1116 3936 1120
rect 3872 1060 3876 1116
rect 3876 1060 3932 1116
rect 3932 1060 3936 1116
rect 3872 1056 3936 1060
rect 3952 1116 4016 1120
rect 3952 1060 3956 1116
rect 3956 1060 4012 1116
rect 4012 1060 4016 1116
rect 3952 1056 4016 1060
rect 4032 1116 4096 1120
rect 4032 1060 4036 1116
rect 4036 1060 4092 1116
rect 4092 1060 4096 1116
rect 4032 1056 4096 1060
rect 4112 1116 4176 1120
rect 4112 1060 4116 1116
rect 4116 1060 4172 1116
rect 4172 1060 4176 1116
rect 4112 1056 4176 1060
rect 6793 1116 6857 1120
rect 6793 1060 6797 1116
rect 6797 1060 6853 1116
rect 6853 1060 6857 1116
rect 6793 1056 6857 1060
rect 6873 1116 6937 1120
rect 6873 1060 6877 1116
rect 6877 1060 6933 1116
rect 6933 1060 6937 1116
rect 6873 1056 6937 1060
rect 6953 1116 7017 1120
rect 6953 1060 6957 1116
rect 6957 1060 7013 1116
rect 7013 1060 7017 1116
rect 6953 1056 7017 1060
rect 7033 1116 7097 1120
rect 7033 1060 7037 1116
rect 7037 1060 7093 1116
rect 7093 1060 7097 1116
rect 7033 1056 7097 1060
rect 9714 1116 9778 1120
rect 9714 1060 9718 1116
rect 9718 1060 9774 1116
rect 9774 1060 9778 1116
rect 9714 1056 9778 1060
rect 9794 1116 9858 1120
rect 9794 1060 9798 1116
rect 9798 1060 9854 1116
rect 9854 1060 9858 1116
rect 9794 1056 9858 1060
rect 9874 1116 9938 1120
rect 9874 1060 9878 1116
rect 9878 1060 9934 1116
rect 9934 1060 9938 1116
rect 9874 1056 9938 1060
rect 9954 1116 10018 1120
rect 9954 1060 9958 1116
rect 9958 1060 10014 1116
rect 10014 1060 10018 1116
rect 9954 1056 10018 1060
rect 12635 1116 12699 1120
rect 12635 1060 12639 1116
rect 12639 1060 12695 1116
rect 12695 1060 12699 1116
rect 12635 1056 12699 1060
rect 12715 1116 12779 1120
rect 12715 1060 12719 1116
rect 12719 1060 12775 1116
rect 12775 1060 12779 1116
rect 12715 1056 12779 1060
rect 12795 1116 12859 1120
rect 12795 1060 12799 1116
rect 12799 1060 12855 1116
rect 12855 1060 12859 1116
rect 12795 1056 12859 1060
rect 12875 1116 12939 1120
rect 12875 1060 12879 1116
rect 12879 1060 12935 1116
rect 12935 1060 12939 1116
rect 12875 1056 12939 1060
<< metal4 >>
rect 2404 12544 2724 12560
rect 2404 12480 2412 12544
rect 2476 12480 2492 12544
rect 2556 12480 2572 12544
rect 2636 12480 2652 12544
rect 2716 12480 2724 12544
rect 2404 11456 2724 12480
rect 2404 11392 2412 11456
rect 2476 11392 2492 11456
rect 2556 11392 2572 11456
rect 2636 11392 2652 11456
rect 2716 11392 2724 11456
rect 2404 10368 2724 11392
rect 2404 10304 2412 10368
rect 2476 10304 2492 10368
rect 2556 10304 2572 10368
rect 2636 10304 2652 10368
rect 2716 10304 2724 10368
rect 2404 9280 2724 10304
rect 2404 9216 2412 9280
rect 2476 9216 2492 9280
rect 2556 9216 2572 9280
rect 2636 9216 2652 9280
rect 2716 9216 2724 9280
rect 2404 8192 2724 9216
rect 2404 8128 2412 8192
rect 2476 8128 2492 8192
rect 2556 8128 2572 8192
rect 2636 8128 2652 8192
rect 2716 8128 2724 8192
rect 2404 7104 2724 8128
rect 2404 7040 2412 7104
rect 2476 7040 2492 7104
rect 2556 7040 2572 7104
rect 2636 7040 2652 7104
rect 2716 7040 2724 7104
rect 2404 6016 2724 7040
rect 2404 5952 2412 6016
rect 2476 5952 2492 6016
rect 2556 5952 2572 6016
rect 2636 5952 2652 6016
rect 2716 5952 2724 6016
rect 2404 4928 2724 5952
rect 2404 4864 2412 4928
rect 2476 4864 2492 4928
rect 2556 4864 2572 4928
rect 2636 4864 2652 4928
rect 2716 4864 2724 4928
rect 2404 3840 2724 4864
rect 2404 3776 2412 3840
rect 2476 3776 2492 3840
rect 2556 3776 2572 3840
rect 2636 3776 2652 3840
rect 2716 3776 2724 3840
rect 2404 2752 2724 3776
rect 2404 2688 2412 2752
rect 2476 2688 2492 2752
rect 2556 2688 2572 2752
rect 2636 2688 2652 2752
rect 2716 2688 2724 2752
rect 2404 1664 2724 2688
rect 2404 1600 2412 1664
rect 2476 1600 2492 1664
rect 2556 1600 2572 1664
rect 2636 1600 2652 1664
rect 2716 1600 2724 1664
rect 2404 1040 2724 1600
rect 3864 12000 4184 12560
rect 3864 11936 3872 12000
rect 3936 11936 3952 12000
rect 4016 11936 4032 12000
rect 4096 11936 4112 12000
rect 4176 11936 4184 12000
rect 3864 10912 4184 11936
rect 3864 10848 3872 10912
rect 3936 10848 3952 10912
rect 4016 10848 4032 10912
rect 4096 10848 4112 10912
rect 4176 10848 4184 10912
rect 3864 9824 4184 10848
rect 3864 9760 3872 9824
rect 3936 9760 3952 9824
rect 4016 9760 4032 9824
rect 4096 9760 4112 9824
rect 4176 9760 4184 9824
rect 3864 8736 4184 9760
rect 3864 8672 3872 8736
rect 3936 8672 3952 8736
rect 4016 8672 4032 8736
rect 4096 8672 4112 8736
rect 4176 8672 4184 8736
rect 3864 7648 4184 8672
rect 3864 7584 3872 7648
rect 3936 7584 3952 7648
rect 4016 7584 4032 7648
rect 4096 7584 4112 7648
rect 4176 7584 4184 7648
rect 3864 6560 4184 7584
rect 3864 6496 3872 6560
rect 3936 6496 3952 6560
rect 4016 6496 4032 6560
rect 4096 6496 4112 6560
rect 4176 6496 4184 6560
rect 3864 5472 4184 6496
rect 3864 5408 3872 5472
rect 3936 5408 3952 5472
rect 4016 5408 4032 5472
rect 4096 5408 4112 5472
rect 4176 5408 4184 5472
rect 3864 4384 4184 5408
rect 3864 4320 3872 4384
rect 3936 4320 3952 4384
rect 4016 4320 4032 4384
rect 4096 4320 4112 4384
rect 4176 4320 4184 4384
rect 3864 3296 4184 4320
rect 3864 3232 3872 3296
rect 3936 3232 3952 3296
rect 4016 3232 4032 3296
rect 4096 3232 4112 3296
rect 4176 3232 4184 3296
rect 3864 2208 4184 3232
rect 3864 2144 3872 2208
rect 3936 2144 3952 2208
rect 4016 2144 4032 2208
rect 4096 2144 4112 2208
rect 4176 2144 4184 2208
rect 3864 1120 4184 2144
rect 3864 1056 3872 1120
rect 3936 1056 3952 1120
rect 4016 1056 4032 1120
rect 4096 1056 4112 1120
rect 4176 1056 4184 1120
rect 3864 1040 4184 1056
rect 5325 12544 5645 12560
rect 5325 12480 5333 12544
rect 5397 12480 5413 12544
rect 5477 12480 5493 12544
rect 5557 12480 5573 12544
rect 5637 12480 5645 12544
rect 5325 11456 5645 12480
rect 5325 11392 5333 11456
rect 5397 11392 5413 11456
rect 5477 11392 5493 11456
rect 5557 11392 5573 11456
rect 5637 11392 5645 11456
rect 5325 10368 5645 11392
rect 5325 10304 5333 10368
rect 5397 10304 5413 10368
rect 5477 10304 5493 10368
rect 5557 10304 5573 10368
rect 5637 10304 5645 10368
rect 5325 9280 5645 10304
rect 5325 9216 5333 9280
rect 5397 9216 5413 9280
rect 5477 9216 5493 9280
rect 5557 9216 5573 9280
rect 5637 9216 5645 9280
rect 5325 8192 5645 9216
rect 5325 8128 5333 8192
rect 5397 8128 5413 8192
rect 5477 8128 5493 8192
rect 5557 8128 5573 8192
rect 5637 8128 5645 8192
rect 5325 7104 5645 8128
rect 5325 7040 5333 7104
rect 5397 7040 5413 7104
rect 5477 7040 5493 7104
rect 5557 7040 5573 7104
rect 5637 7040 5645 7104
rect 5325 6016 5645 7040
rect 5325 5952 5333 6016
rect 5397 5952 5413 6016
rect 5477 5952 5493 6016
rect 5557 5952 5573 6016
rect 5637 5952 5645 6016
rect 5325 4928 5645 5952
rect 5325 4864 5333 4928
rect 5397 4864 5413 4928
rect 5477 4864 5493 4928
rect 5557 4864 5573 4928
rect 5637 4864 5645 4928
rect 5325 3840 5645 4864
rect 5325 3776 5333 3840
rect 5397 3776 5413 3840
rect 5477 3776 5493 3840
rect 5557 3776 5573 3840
rect 5637 3776 5645 3840
rect 5325 2752 5645 3776
rect 5325 2688 5333 2752
rect 5397 2688 5413 2752
rect 5477 2688 5493 2752
rect 5557 2688 5573 2752
rect 5637 2688 5645 2752
rect 5325 1664 5645 2688
rect 5325 1600 5333 1664
rect 5397 1600 5413 1664
rect 5477 1600 5493 1664
rect 5557 1600 5573 1664
rect 5637 1600 5645 1664
rect 5325 1040 5645 1600
rect 6785 12000 7105 12560
rect 6785 11936 6793 12000
rect 6857 11936 6873 12000
rect 6937 11936 6953 12000
rect 7017 11936 7033 12000
rect 7097 11936 7105 12000
rect 6785 10912 7105 11936
rect 6785 10848 6793 10912
rect 6857 10848 6873 10912
rect 6937 10848 6953 10912
rect 7017 10848 7033 10912
rect 7097 10848 7105 10912
rect 6785 9824 7105 10848
rect 6785 9760 6793 9824
rect 6857 9760 6873 9824
rect 6937 9760 6953 9824
rect 7017 9760 7033 9824
rect 7097 9760 7105 9824
rect 6785 8736 7105 9760
rect 6785 8672 6793 8736
rect 6857 8672 6873 8736
rect 6937 8672 6953 8736
rect 7017 8672 7033 8736
rect 7097 8672 7105 8736
rect 6785 7648 7105 8672
rect 6785 7584 6793 7648
rect 6857 7584 6873 7648
rect 6937 7584 6953 7648
rect 7017 7584 7033 7648
rect 7097 7584 7105 7648
rect 6785 6560 7105 7584
rect 6785 6496 6793 6560
rect 6857 6496 6873 6560
rect 6937 6496 6953 6560
rect 7017 6496 7033 6560
rect 7097 6496 7105 6560
rect 6785 5472 7105 6496
rect 6785 5408 6793 5472
rect 6857 5408 6873 5472
rect 6937 5408 6953 5472
rect 7017 5408 7033 5472
rect 7097 5408 7105 5472
rect 6785 4384 7105 5408
rect 6785 4320 6793 4384
rect 6857 4320 6873 4384
rect 6937 4320 6953 4384
rect 7017 4320 7033 4384
rect 7097 4320 7105 4384
rect 6785 3296 7105 4320
rect 6785 3232 6793 3296
rect 6857 3232 6873 3296
rect 6937 3232 6953 3296
rect 7017 3232 7033 3296
rect 7097 3232 7105 3296
rect 6785 2208 7105 3232
rect 6785 2144 6793 2208
rect 6857 2144 6873 2208
rect 6937 2144 6953 2208
rect 7017 2144 7033 2208
rect 7097 2144 7105 2208
rect 6785 1120 7105 2144
rect 6785 1056 6793 1120
rect 6857 1056 6873 1120
rect 6937 1056 6953 1120
rect 7017 1056 7033 1120
rect 7097 1056 7105 1120
rect 6785 1040 7105 1056
rect 8246 12544 8566 12560
rect 8246 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8494 12544
rect 8558 12480 8566 12544
rect 8246 11456 8566 12480
rect 8246 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8494 11456
rect 8558 11392 8566 11456
rect 8246 10368 8566 11392
rect 8246 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8494 10368
rect 8558 10304 8566 10368
rect 8246 9280 8566 10304
rect 8246 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8494 9280
rect 8558 9216 8566 9280
rect 8246 8192 8566 9216
rect 8246 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8494 8192
rect 8558 8128 8566 8192
rect 8246 7104 8566 8128
rect 8246 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8494 7104
rect 8558 7040 8566 7104
rect 8246 6016 8566 7040
rect 8246 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8494 6016
rect 8558 5952 8566 6016
rect 8246 4928 8566 5952
rect 8246 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8494 4928
rect 8558 4864 8566 4928
rect 8246 3840 8566 4864
rect 8246 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8494 3840
rect 8558 3776 8566 3840
rect 8246 2752 8566 3776
rect 8246 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8494 2752
rect 8558 2688 8566 2752
rect 8246 1664 8566 2688
rect 8246 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8494 1664
rect 8558 1600 8566 1664
rect 8246 1040 8566 1600
rect 9706 12000 10026 12560
rect 9706 11936 9714 12000
rect 9778 11936 9794 12000
rect 9858 11936 9874 12000
rect 9938 11936 9954 12000
rect 10018 11936 10026 12000
rect 9706 10912 10026 11936
rect 9706 10848 9714 10912
rect 9778 10848 9794 10912
rect 9858 10848 9874 10912
rect 9938 10848 9954 10912
rect 10018 10848 10026 10912
rect 9706 9824 10026 10848
rect 9706 9760 9714 9824
rect 9778 9760 9794 9824
rect 9858 9760 9874 9824
rect 9938 9760 9954 9824
rect 10018 9760 10026 9824
rect 9706 8736 10026 9760
rect 9706 8672 9714 8736
rect 9778 8672 9794 8736
rect 9858 8672 9874 8736
rect 9938 8672 9954 8736
rect 10018 8672 10026 8736
rect 9706 7648 10026 8672
rect 9706 7584 9714 7648
rect 9778 7584 9794 7648
rect 9858 7584 9874 7648
rect 9938 7584 9954 7648
rect 10018 7584 10026 7648
rect 9706 6560 10026 7584
rect 9706 6496 9714 6560
rect 9778 6496 9794 6560
rect 9858 6496 9874 6560
rect 9938 6496 9954 6560
rect 10018 6496 10026 6560
rect 9706 5472 10026 6496
rect 9706 5408 9714 5472
rect 9778 5408 9794 5472
rect 9858 5408 9874 5472
rect 9938 5408 9954 5472
rect 10018 5408 10026 5472
rect 9706 4384 10026 5408
rect 9706 4320 9714 4384
rect 9778 4320 9794 4384
rect 9858 4320 9874 4384
rect 9938 4320 9954 4384
rect 10018 4320 10026 4384
rect 9706 3296 10026 4320
rect 9706 3232 9714 3296
rect 9778 3232 9794 3296
rect 9858 3232 9874 3296
rect 9938 3232 9954 3296
rect 10018 3232 10026 3296
rect 9706 2208 10026 3232
rect 9706 2144 9714 2208
rect 9778 2144 9794 2208
rect 9858 2144 9874 2208
rect 9938 2144 9954 2208
rect 10018 2144 10026 2208
rect 9706 1120 10026 2144
rect 9706 1056 9714 1120
rect 9778 1056 9794 1120
rect 9858 1056 9874 1120
rect 9938 1056 9954 1120
rect 10018 1056 10026 1120
rect 9706 1040 10026 1056
rect 11167 12544 11487 12560
rect 11167 12480 11175 12544
rect 11239 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11487 12544
rect 11167 11456 11487 12480
rect 11167 11392 11175 11456
rect 11239 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11487 11456
rect 11167 10368 11487 11392
rect 11167 10304 11175 10368
rect 11239 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11487 10368
rect 11167 9280 11487 10304
rect 11167 9216 11175 9280
rect 11239 9216 11255 9280
rect 11319 9216 11335 9280
rect 11399 9216 11415 9280
rect 11479 9216 11487 9280
rect 11167 8192 11487 9216
rect 11167 8128 11175 8192
rect 11239 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11487 8192
rect 11167 7104 11487 8128
rect 11167 7040 11175 7104
rect 11239 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11487 7104
rect 11167 6016 11487 7040
rect 11167 5952 11175 6016
rect 11239 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11487 6016
rect 11167 4928 11487 5952
rect 11167 4864 11175 4928
rect 11239 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11487 4928
rect 11167 3840 11487 4864
rect 11167 3776 11175 3840
rect 11239 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11487 3840
rect 11167 2752 11487 3776
rect 11167 2688 11175 2752
rect 11239 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11487 2752
rect 11167 1664 11487 2688
rect 11167 1600 11175 1664
rect 11239 1600 11255 1664
rect 11319 1600 11335 1664
rect 11399 1600 11415 1664
rect 11479 1600 11487 1664
rect 11167 1040 11487 1600
rect 12627 12000 12947 12560
rect 12627 11936 12635 12000
rect 12699 11936 12715 12000
rect 12779 11936 12795 12000
rect 12859 11936 12875 12000
rect 12939 11936 12947 12000
rect 12627 10912 12947 11936
rect 12627 10848 12635 10912
rect 12699 10848 12715 10912
rect 12779 10848 12795 10912
rect 12859 10848 12875 10912
rect 12939 10848 12947 10912
rect 12627 9824 12947 10848
rect 12627 9760 12635 9824
rect 12699 9760 12715 9824
rect 12779 9760 12795 9824
rect 12859 9760 12875 9824
rect 12939 9760 12947 9824
rect 12627 8736 12947 9760
rect 12627 8672 12635 8736
rect 12699 8672 12715 8736
rect 12779 8672 12795 8736
rect 12859 8672 12875 8736
rect 12939 8672 12947 8736
rect 12627 7648 12947 8672
rect 12627 7584 12635 7648
rect 12699 7584 12715 7648
rect 12779 7584 12795 7648
rect 12859 7584 12875 7648
rect 12939 7584 12947 7648
rect 12627 6560 12947 7584
rect 12627 6496 12635 6560
rect 12699 6496 12715 6560
rect 12779 6496 12795 6560
rect 12859 6496 12875 6560
rect 12939 6496 12947 6560
rect 12627 5472 12947 6496
rect 12627 5408 12635 5472
rect 12699 5408 12715 5472
rect 12779 5408 12795 5472
rect 12859 5408 12875 5472
rect 12939 5408 12947 5472
rect 12627 4384 12947 5408
rect 12627 4320 12635 4384
rect 12699 4320 12715 4384
rect 12779 4320 12795 4384
rect 12859 4320 12875 4384
rect 12939 4320 12947 4384
rect 12627 3296 12947 4320
rect 12627 3232 12635 3296
rect 12699 3232 12715 3296
rect 12779 3232 12795 3296
rect 12859 3232 12875 3296
rect 12939 3232 12947 3296
rect 12627 2208 12947 3232
rect 12627 2144 12635 2208
rect 12699 2144 12715 2208
rect 12779 2144 12795 2208
rect 12859 2144 12875 2208
rect 12939 2144 12947 2208
rect 12627 1120 12947 2144
rect 12627 1056 12635 1120
rect 12699 1056 12715 1120
rect 12779 1056 12795 1120
rect 12859 1056 12875 1120
rect 12939 1056 12947 1120
rect 12627 1040 12947 1056
use sky130_fd_sc_hd__buf_2  _115_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _116_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _117_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6256 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _118_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _119_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4048 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _120_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _122_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _123_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _124_
timestamp 1701704242
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _125_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6992 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _126_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1701704242
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1701704242
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1701704242
transform -1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _130_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _131_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132_
timestamp 1701704242
transform -1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _133_
timestamp 1701704242
transform 1 0 7636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 1701704242
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1701704242
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _136_
timestamp 1701704242
transform 1 0 7268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 1701704242
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1701704242
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _139_
timestamp 1701704242
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _140_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9752 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1701704242
transform -1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _142_
timestamp 1701704242
transform 1 0 7176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _143_
timestamp 1701704242
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _144_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _145_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _146_
timestamp 1701704242
transform 1 0 7268 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _147_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _148_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7728 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _149_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _150_
timestamp 1701704242
transform -1 0 5244 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _151_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 3680 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _152_
timestamp 1701704242
transform 1 0 3680 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _153_
timestamp 1701704242
transform 1 0 3956 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _154_
timestamp 1701704242
transform 1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _155_
timestamp 1701704242
transform 1 0 8832 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1701704242
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _157_
timestamp 1701704242
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _158_
timestamp 1701704242
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1701704242
transform -1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _160_
timestamp 1701704242
transform -1 0 8740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _161_
timestamp 1701704242
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _162_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9752 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _163_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10672 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _164_
timestamp 1701704242
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _165_
timestamp 1701704242
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1701704242
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1701704242
transform 1 0 5704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _168_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _169_
timestamp 1701704242
transform -1 0 3312 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1701704242
transform -1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _171_
timestamp 1701704242
transform 1 0 1932 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _172_
timestamp 1701704242
transform 1 0 3956 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _173_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _174_
timestamp 1701704242
transform 1 0 3956 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _175_
timestamp 1701704242
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _176_
timestamp 1701704242
transform 1 0 3036 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _177_
timestamp 1701704242
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _178_
timestamp 1701704242
transform 1 0 2852 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _179_
timestamp 1701704242
transform 1 0 1656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _180_
timestamp 1701704242
transform 1 0 2944 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _181_
timestamp 1701704242
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _182_
timestamp 1701704242
transform -1 0 3404 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _183_
timestamp 1701704242
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 1701704242
transform -1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _185_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 3680 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _186_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4324 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _187_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4232 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1701704242
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _189_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6624 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _190_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 7728 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1701704242
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _193_
timestamp 1701704242
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _194_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6164 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _195_
timestamp 1701704242
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 1701704242
transform 1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _197_
timestamp 1701704242
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _198_
timestamp 1701704242
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _199_
timestamp 1701704242
transform 1 0 5520 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _200_
timestamp 1701704242
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1701704242
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _202_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _203_
timestamp 1701704242
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _204_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 4784 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _205_
timestamp 1701704242
transform -1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1701704242
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1701704242
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _208_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5980 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _209_
timestamp 1701704242
transform 1 0 2944 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _210_
timestamp 1701704242
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _211_
timestamp 1701704242
transform 1 0 1380 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1701704242
transform 1 0 2024 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1701704242
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _214_
timestamp 1701704242
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _215_
timestamp 1701704242
transform 1 0 5336 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _216_
timestamp 1701704242
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _217_
timestamp 1701704242
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1701704242
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1701704242
transform 1 0 4324 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp 1701704242
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _221_
timestamp 1701704242
transform -1 0 5336 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _222_
timestamp 1701704242
transform 1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _223_
timestamp 1701704242
transform 1 0 3772 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 1701704242
transform 1 0 3128 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _225_
timestamp 1701704242
transform 1 0 6348 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 1701704242
transform 1 0 6992 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1701704242
transform -1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _228_
timestamp 1701704242
transform -1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _229_
timestamp 1701704242
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _230_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _231_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _232_
timestamp 1701704242
transform 1 0 2668 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _233_
timestamp 1701704242
transform 1 0 1380 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _234_
timestamp 1701704242
transform 1 0 1380 0 1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _235_
timestamp 1701704242
transform -1 0 3772 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _236_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3496 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1701704242
transform 1 0 4232 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _238_
timestamp 1701704242
transform 1 0 7268 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _239_
timestamp 1701704242
transform 1 0 5612 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _240_
timestamp 1701704242
transform 1 0 6348 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _241_
timestamp 1701704242
transform 1 0 6072 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _242_
timestamp 1701704242
transform 1 0 3772 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _243_
timestamp 1701704242
transform 1 0 1472 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1701704242
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1701704242
transform 1 0 1380 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1701704242
transform 1 0 2484 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1701704242
transform 1 0 4784 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1701704242
transform 1 0 2300 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _249_
timestamp 1701704242
transform 1 0 7268 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _250_
timestamp 1701704242
transform 1 0 7360 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _269_
timestamp 1701704242
transform -1 0 3680 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _270_
timestamp 1701704242
transform -1 0 4784 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout3
timestamp 1701704242
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout4
timestamp 1701704242
transform -1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout5
timestamp 1701704242
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout6
timestamp 1701704242
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 1701704242
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout8
timestamp 1701704242
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1701704242
transform -1 0 1748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout12
timestamp 1701704242
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_19 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_39 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4692 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_46 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5336 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1701704242
transform 1 0 6900 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1701704242
transform 1 0 11500 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_121
timestamp 1701704242
transform 1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_7
timestamp 1701704242
transform 1 0 1748 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_83
timestamp 1701704242
transform 1 0 8740 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_95
timestamp 1701704242
transform 1 0 9844 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1701704242
transform 1 0 11500 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_121
timestamp 1701704242
transform 1 0 12236 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_9
timestamp 1701704242
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_21
timestamp 1701704242
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1701704242
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_44
timestamp 1701704242
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_56
timestamp 1701704242
transform 1 0 6256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_64
timestamp 1701704242
transform 1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1701704242
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_109
timestamp 1701704242
transform 1 0 11132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_120
timestamp 1701704242
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_38
timestamp 1701704242
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_43
timestamp 1701704242
transform 1 0 5060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_106
timestamp 1701704242
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1701704242
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_120
timestamp 1701704242
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1701704242
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_58
timestamp 1701704242
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_70
timestamp 1701704242
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1701704242
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1701704242
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_120
timestamp 1701704242
transform 1 0 12144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1701704242
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_11
timestamp 1701704242
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_18
timestamp 1701704242
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_22
timestamp 1701704242
transform 1 0 3128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_33
timestamp 1701704242
transform 1 0 4140 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_41
timestamp 1701704242
transform 1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_46
timestamp 1701704242
transform 1 0 5336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_50
timestamp 1701704242
transform 1 0 5704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1701704242
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_69
timestamp 1701704242
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_80
timestamp 1701704242
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_88
timestamp 1701704242
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_94
timestamp 1701704242
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1701704242
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_19
timestamp 1701704242
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_46
timestamp 1701704242
transform 1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_71
timestamp 1701704242
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_80
timestamp 1701704242
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_100
timestamp 1701704242
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_112
timestamp 1701704242
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_121
timestamp 1701704242
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1701704242
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_17
timestamp 1701704242
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_29
timestamp 1701704242
transform 1 0 3772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_44
timestamp 1701704242
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_63
timestamp 1701704242
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_73
timestamp 1701704242
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_80
timestamp 1701704242
transform 1 0 8464 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_88
timestamp 1701704242
transform 1 0 9200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_94
timestamp 1701704242
transform 1 0 9752 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1701704242
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_117
timestamp 1701704242
transform 1 0 11868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_123
timestamp 1701704242
transform 1 0 12420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1701704242
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_21
timestamp 1701704242
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_40
timestamp 1701704242
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_44
timestamp 1701704242
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_61
timestamp 1701704242
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_65
timestamp 1701704242
transform 1 0 7084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_72
timestamp 1701704242
transform 1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_106
timestamp 1701704242
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1701704242
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_19
timestamp 1701704242
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1701704242
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 1701704242
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_82
timestamp 1701704242
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_94
timestamp 1701704242
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1701704242
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_123
timestamp 1701704242
transform 1 0 12420 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_22
timestamp 1701704242
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_46
timestamp 1701704242
transform 1 0 5336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_54
timestamp 1701704242
transform 1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_63
timestamp 1701704242
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1701704242
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_99
timestamp 1701704242
transform 1 0 10212 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_117
timestamp 1701704242
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_123
timestamp 1701704242
transform 1 0 12420 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1701704242
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_14
timestamp 1701704242
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_25
timestamp 1701704242
transform 1 0 3404 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_74
timestamp 1701704242
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_87
timestamp 1701704242
transform 1 0 9108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_93
timestamp 1701704242
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_97
timestamp 1701704242
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1701704242
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1701704242
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_20
timestamp 1701704242
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_49
timestamp 1701704242
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_64
timestamp 1701704242
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1701704242
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_106
timestamp 1701704242
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 1701704242
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_14
timestamp 1701704242
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_50
timestamp 1701704242
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_60
timestamp 1701704242
transform 1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_64
timestamp 1701704242
transform 1 0 6992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_68
timestamp 1701704242
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_83
timestamp 1701704242
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_91
timestamp 1701704242
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_99
timestamp 1701704242
transform 1 0 10212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1701704242
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1701704242
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_122
timestamp 1701704242
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_7
timestamp 1701704242
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_33
timestamp 1701704242
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_43
timestamp 1701704242
transform 1 0 5060 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_66
timestamp 1701704242
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_74
timestamp 1701704242
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_104
timestamp 1701704242
transform 1 0 10672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_115
timestamp 1701704242
transform 1 0 11684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_121
timestamp 1701704242
transform 1 0 12236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_3
timestamp 1701704242
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_14
timestamp 1701704242
transform 1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_18
timestamp 1701704242
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_26
timestamp 1701704242
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_38
timestamp 1701704242
transform 1 0 4600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_46
timestamp 1701704242
transform 1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_69
timestamp 1701704242
transform 1 0 7452 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_78
timestamp 1701704242
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_84
timestamp 1701704242
transform 1 0 8832 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_92
timestamp 1701704242
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_98
timestamp 1701704242
transform 1 0 10120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1701704242
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1701704242
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_121
timestamp 1701704242
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_42
timestamp 1701704242
transform 1 0 4968 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_55
timestamp 1701704242
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_59
timestamp 1701704242
transform 1 0 6532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_72
timestamp 1701704242
transform 1 0 7728 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1701704242
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 1701704242
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_95
timestamp 1701704242
transform 1 0 9844 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_101
timestamp 1701704242
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_114
timestamp 1701704242
transform 1 0 11592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_120
timestamp 1701704242
transform 1 0 12144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 1701704242
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_14
timestamp 1701704242
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_24
timestamp 1701704242
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_45
timestamp 1701704242
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_62
timestamp 1701704242
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_66
timestamp 1701704242
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_84
timestamp 1701704242
transform 1 0 8832 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1701704242
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_123
timestamp 1701704242
transform 1 0 12420 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_22
timestamp 1701704242
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_40
timestamp 1701704242
transform 1 0 4784 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_52
timestamp 1701704242
transform 1 0 5888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_58
timestamp 1701704242
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_74
timestamp 1701704242
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1701704242
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1701704242
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_105
timestamp 1701704242
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_117
timestamp 1701704242
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1701704242
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_11
timestamp 1701704242
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_29
timestamp 1701704242
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_60
timestamp 1701704242
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_72
timestamp 1701704242
transform 1 0 7728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_76
timestamp 1701704242
transform 1 0 8096 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_80
timestamp 1701704242
transform 1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_97
timestamp 1701704242
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1701704242
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1701704242
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 1701704242
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_21
timestamp 1701704242
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 1701704242
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_40
timestamp 1701704242
transform 1 0 4784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1701704242
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_64
timestamp 1701704242
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_78
timestamp 1701704242
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1701704242
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_94
timestamp 1701704242
transform 1 0 9752 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_113
timestamp 1701704242
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_121
timestamp 1701704242
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1701704242
transform 1 0 3772 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap9
timestamp 1701704242
transform -1 0 6440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_21
timestamp 1701704242
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 12788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_22
timestamp 1701704242
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 12788 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_23
timestamp 1701704242
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_24
timestamp 1701704242
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_25
timestamp 1701704242
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_26
timestamp 1701704242
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_27
timestamp 1701704242
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_28
timestamp 1701704242
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_29
timestamp 1701704242
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_30
timestamp 1701704242
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_31
timestamp 1701704242
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_32
timestamp 1701704242
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_33
timestamp 1701704242
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_34
timestamp 1701704242
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_35
timestamp 1701704242
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_36
timestamp 1701704242
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_37
timestamp 1701704242
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_38
timestamp 1701704242
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_39
timestamp 1701704242
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_40
timestamp 1701704242
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_41
timestamp 1701704242
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 1701704242
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_44
timestamp 1701704242
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_45
timestamp 1701704242
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp 1701704242
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp 1701704242
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp 1701704242
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp 1701704242
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp 1701704242
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp 1701704242
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 1701704242
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 1701704242
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 1701704242
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_55
timestamp 1701704242
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 1701704242
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1701704242
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_58
timestamp 1701704242
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_59
timestamp 1701704242
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_60
timestamp 1701704242
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_61
timestamp 1701704242
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_62
timestamp 1701704242
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_63
timestamp 1701704242
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_64
timestamp 1701704242
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_65
timestamp 1701704242
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_66
timestamp 1701704242
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_67
timestamp 1701704242
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_68
timestamp 1701704242
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_69
timestamp 1701704242
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_70
timestamp 1701704242
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_71
timestamp 1701704242
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_72
timestamp 1701704242
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_73
timestamp 1701704242
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_74
timestamp 1701704242
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_75
timestamp 1701704242
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_76
timestamp 1701704242
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_77
timestamp 1701704242
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_78
timestamp 1701704242
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_79
timestamp 1701704242
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_80
timestamp 1701704242
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_81
timestamp 1701704242
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_82
timestamp 1701704242
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_83
timestamp 1701704242
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_84
timestamp 1701704242
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_85
timestamp 1701704242
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_86
timestamp 1701704242
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_87
timestamp 1701704242
transform 1 0 11408 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[0\].cap
timestamp 1701704242
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[0\].cap_13 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[1\].cap
timestamp 1701704242
transform -1 0 8280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[1\].cap_20
timestamp 1701704242
transform 1 0 7176 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[2\].cap
timestamp 1701704242
transform -1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[2\].cap_21
timestamp 1701704242
transform 1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[3\].cap
timestamp 1701704242
transform -1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[3\].cap_22
timestamp 1701704242
transform 1 0 5428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[4\].cap_23
timestamp 1701704242
transform -1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[4\].cap
timestamp 1701704242
transform 1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[5\].cap_24
timestamp 1701704242
transform -1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[5\].cap
timestamp 1701704242
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[6\].cap_25
timestamp 1701704242
transform -1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[6\].cap
timestamp 1701704242
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[7\].cap
timestamp 1701704242
transform -1 0 6256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[7\].cap_26
timestamp 1701704242
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[8\].cap
timestamp 1701704242
transform -1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[8\].cap_27
timestamp 1701704242
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[9\].cap_28
timestamp 1701704242
transform -1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[9\].cap
timestamp 1701704242
transform 1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[10\].cap_14
timestamp 1701704242
transform -1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[10\].cap
timestamp 1701704242
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[11\].cap_15
timestamp 1701704242
transform -1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[11\].cap
timestamp 1701704242
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[12\].cap_16
timestamp 1701704242
transform -1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[12\].cap
timestamp 1701704242
transform 1 0 7452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[13\].cap
timestamp 1701704242
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[13\].cap_17
timestamp 1701704242
transform -1 0 8648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[14\].cap
timestamp 1701704242
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[14\].cap_18
timestamp 1701704242
transform -1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[15\].cap_19
timestamp 1701704242
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[15\].cap
timestamp 1701704242
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10396 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 10396 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform -1 0 10948 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform -1 0 11408 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform -1 0 10488 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 11408 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform -1 0 10304 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform -1 0 8464 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform 1 0 9292 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 8004 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 9384 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform 1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform 1 0 8004 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform 1 0 9752 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 11776 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform 1 0 9936 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 10764 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 9384 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 10672 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform -1 0 11224 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform -1 0 11224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1701704242
transform 1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1701704242
transform 1 0 11684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1701704242
transform 1 0 9660 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1701704242
transform 1 0 11776 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1701704242
transform -1 0 10304 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1701704242
transform 1 0 11224 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1701704242
transform -1 0 10764 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1701704242
transform 1 0 11868 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform 1 0 10396 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 12052 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform -1 0 12144 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 10304 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 11960 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform 1 0 10948 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform 1 0 11500 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1701704242
transform 1 0 11684 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1701704242
transform 1 0 10948 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1701704242
transform 1 0 11684 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1701704242
transform -1 0 12052 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1701704242
transform 1 0 9844 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1701704242
transform 1 0 11960 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1701704242
transform 1 0 11776 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1701704242
transform 1 0 12052 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1701704242
transform 1 0 10764 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1701704242
transform 1 0 12052 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1701704242
transform 1 0 10488 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1701704242
transform 1 0 11592 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1701704242
transform 1 0 10488 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1701704242
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1701704242
transform -1 0 12052 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1701704242
transform 1 0 11132 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1701704242
transform 1 0 12052 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1701704242
transform 1 0 11592 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1701704242
transform -1 0 12512 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1701704242
transform -1 0 11224 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1701704242
transform 1 0 11224 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1701704242
transform 1 0 11132 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1701704242
transform 1 0 10948 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1701704242
transform 1 0 11408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd_30
timestamp 1701704242
transform 1 0 8004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1701704242
transform 1 0 7544 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].vref_29
timestamp 1701704242
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 12052 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dcdc
timestamp 1701704242
transform 1 0 6532 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  temp1.inv1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2
timestamp 1701704242
transform -1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire10
timestamp 1701704242
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 552 400 672 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 1368 400 1488 0 FreeSans 480 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 0 2184 400 2304 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal3 s 0 3000 400 3120 0 FreeSans 480 0 0 0 io_in[3]
port 3 nsew signal input
flabel metal3 s 0 3816 400 3936 0 FreeSans 480 0 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 0 4632 400 4752 0 FreeSans 480 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal3 s 0 5448 400 5568 0 FreeSans 480 0 0 0 io_in[6]
port 6 nsew signal input
flabel metal3 s 0 6264 400 6384 0 FreeSans 480 0 0 0 io_in[7]
port 7 nsew signal input
flabel metal3 s 0 7080 400 7200 0 FreeSans 480 0 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal3 s 0 7896 400 8016 0 FreeSans 480 0 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal3 s 0 8712 400 8832 0 FreeSans 480 0 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal3 s 0 10344 400 10464 0 FreeSans 480 0 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal3 s 0 11160 400 11280 0 FreeSans 480 0 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal3 s 0 11976 400 12096 0 FreeSans 480 0 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal3 s 0 12792 400 12912 0 FreeSans 480 0 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 2404 1040 2724 12560 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 5325 1040 5645 12560 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 8246 1040 8566 12560 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 11167 1040 11487 12560 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 3864 1040 4184 12560 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 6785 1040 7105 12560 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 9706 1040 10026 12560 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 12627 1040 12947 12560 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 6946 12512 6946 12512 0 vccd1
rlabel via1 7025 11968 7025 11968 0 vssd1
rlabel metal2 1702 7004 1702 7004 0 _000_
rlabel via1 1697 7854 1697 7854 0 _001_
rlabel metal1 3169 8534 3169 8534 0 _002_
rlabel metal2 1702 9860 1702 9860 0 _003_
rlabel metal2 1702 10948 1702 10948 0 _004_
rlabel metal2 3818 11526 3818 11526 0 _005_
rlabel metal2 4370 10438 4370 10438 0 _006_
rlabel metal1 4687 8534 4687 8534 0 _007_
rlabel metal1 7636 10234 7636 10234 0 _008_
rlabel metal1 5832 8942 5832 8942 0 _009_
rlabel metal1 6440 6970 6440 6970 0 _010_
rlabel metal1 5964 4522 5964 4522 0 _011_
rlabel metal2 3450 6290 3450 6290 0 _012_
rlabel metal2 1978 5474 1978 5474 0 _013_
rlabel metal2 2254 4386 2254 4386 0 _014_
rlabel via1 1697 1326 1697 1326 0 _015_
rlabel metal1 2985 3026 2985 3026 0 _016_
rlabel metal1 5106 1530 5106 1530 0 _017_
rlabel metal2 3174 1734 3174 1734 0 _018_
rlabel metal1 7482 2006 7482 2006 0 _019_
rlabel metal1 7580 3026 7580 3026 0 _020_
rlabel metal1 3220 4250 3220 4250 0 _021_
rlabel metal1 4370 4658 4370 4658 0 _022_
rlabel metal1 4738 3502 4738 3502 0 _023_
rlabel metal1 6900 3026 6900 3026 0 _024_
rlabel metal1 9338 3094 9338 3094 0 _025_
rlabel via1 8602 2414 8602 2414 0 _026_
rlabel metal1 3266 10676 3266 10676 0 _027_
rlabel metal1 5934 10234 5934 10234 0 _028_
rlabel via1 2714 6901 2714 6901 0 _029_
rlabel metal1 2806 10642 2806 10642 0 _030_
rlabel metal2 2622 10914 2622 10914 0 _031_
rlabel metal1 2760 1734 2760 1734 0 _032_
rlabel metal1 1886 7412 1886 7412 0 _033_
rlabel metal1 2714 8296 2714 8296 0 _034_
rlabel metal2 3082 8500 3082 8500 0 _035_
rlabel metal1 1886 9520 1886 9520 0 _036_
rlabel metal1 1886 10676 1886 10676 0 _037_
rlabel metal1 3588 7242 3588 7242 0 _038_
rlabel metal2 4554 10506 4554 10506 0 _039_
rlabel metal1 2484 4114 2484 4114 0 _040_
rlabel metal1 5014 8976 5014 8976 0 _041_
rlabel metal1 7498 10064 7498 10064 0 _042_
rlabel metal1 6256 8330 6256 8330 0 _043_
rlabel metal1 6164 8602 6164 8602 0 _044_
rlabel metal1 6394 6698 6394 6698 0 _045_
rlabel metal1 6762 6766 6762 6766 0 _046_
rlabel metal2 5934 4352 5934 4352 0 _047_
rlabel metal1 6026 4692 6026 4692 0 _048_
rlabel metal1 5842 3706 5842 3706 0 _049_
rlabel metal1 4232 5746 4232 5746 0 _050_
rlabel metal1 3450 5712 3450 5712 0 _051_
rlabel metal2 4278 5406 4278 5406 0 _052_
rlabel metal1 2208 5202 2208 5202 0 _053_
rlabel metal1 5014 3638 5014 3638 0 _054_
rlabel metal1 2622 4080 2622 4080 0 _055_
rlabel metal2 2990 4284 2990 4284 0 _056_
rlabel metal1 1978 3128 1978 3128 0 _057_
rlabel metal1 2024 2414 2024 2414 0 _058_
rlabel metal1 5198 3162 5198 3162 0 _059_
rlabel metal1 5474 2414 5474 2414 0 _060_
rlabel metal1 3726 2414 3726 2414 0 _061_
rlabel metal1 4830 2346 4830 2346 0 _062_
rlabel metal1 4830 1258 4830 1258 0 _063_
rlabel metal2 4830 1802 4830 1802 0 _064_
rlabel metal1 6164 1870 6164 1870 0 _065_
rlabel metal1 3634 1360 3634 1360 0 _066_
rlabel metal1 6992 1326 6992 1326 0 _067_
rlabel metal1 7222 1530 7222 1530 0 _068_
rlabel metal1 7406 2414 7406 2414 0 _069_
rlabel metal1 4554 11084 4554 11084 0 _070_
rlabel metal1 6578 10540 6578 10540 0 _071_
rlabel metal1 6256 3162 6256 3162 0 _072_
rlabel metal1 4738 11186 4738 11186 0 _073_
rlabel metal1 4692 11730 4692 11730 0 _074_
rlabel metal1 7544 11186 7544 11186 0 _075_
rlabel metal1 7314 5780 7314 5780 0 _076_
rlabel metal1 7314 5168 7314 5168 0 _077_
rlabel metal1 7360 9010 7360 9010 0 _078_
rlabel metal1 8372 8466 8372 8466 0 _079_
rlabel metal1 9568 8806 9568 8806 0 _080_
rlabel metal1 8602 7344 8602 7344 0 _081_
rlabel metal2 7498 5440 7498 5440 0 _082_
rlabel metal1 9338 7752 9338 7752 0 _083_
rlabel metal1 7912 6766 7912 6766 0 _084_
rlabel metal1 9338 6664 9338 6664 0 _085_
rlabel metal1 7360 5270 7360 5270 0 _086_
rlabel metal1 8027 5338 8027 5338 0 _087_
rlabel metal1 8648 8942 8648 8942 0 _088_
rlabel metal1 9430 9010 9430 9010 0 _089_
rlabel metal1 5566 5746 5566 5746 0 _090_
rlabel metal1 7682 5780 7682 5780 0 _091_
rlabel metal1 6716 6290 6716 6290 0 _092_
rlabel metal1 8878 9010 8878 9010 0 _093_
rlabel metal1 7406 6222 7406 6222 0 _094_
rlabel metal1 9210 8942 9210 8942 0 _095_
rlabel metal1 4094 5644 4094 5644 0 _096_
rlabel metal1 5658 7854 5658 7854 0 ctr\[0\]
rlabel metal1 4600 2414 4600 2414 0 ctr\[10\]
rlabel metal1 4002 2074 4002 2074 0 ctr\[11\]
rlabel metal1 6624 1938 6624 1938 0 ctr\[12\]
rlabel metal1 8924 2822 8924 2822 0 ctr\[13\]
rlabel metal1 8602 10030 8602 10030 0 ctr\[1\]
rlabel metal1 8924 7854 8924 7854 0 ctr\[2\]
rlabel metal1 4600 7786 4600 7786 0 ctr\[3\]
rlabel metal2 4002 5814 4002 5814 0 ctr\[4\]
rlabel metal1 9154 9554 9154 9554 0 ctr\[5\]
rlabel metal1 6670 5644 6670 5644 0 ctr\[6\]
rlabel metal1 2944 4794 2944 4794 0 ctr\[7\]
rlabel metal1 1610 2958 1610 2958 0 ctr\[8\]
rlabel metal1 5612 5678 5612 5678 0 ctr\[9\]
rlabel metal1 4094 11866 4094 11866 0 in_measurement
rlabel metal3 2062 612 2062 612 0 io_in[0]
rlabel metal3 544 1428 544 1428 0 io_in[1]
rlabel metal2 1794 7055 1794 7055 0 io_out[0]
rlabel metal1 2346 8432 2346 8432 0 io_out[1]
rlabel metal1 1334 8976 1334 8976 0 io_out[2]
rlabel metal2 1794 9741 1794 9741 0 io_out[3]
rlabel metal1 2346 10608 2346 10608 0 io_out[4]
rlabel metal1 1840 11526 1840 11526 0 io_out[5]
rlabel metal3 820 12036 820 12036 0 io_out[6]
rlabel metal3 2338 12852 2338 12852 0 io_out[7]
rlabel metal1 1702 2006 1702 2006 0 net1
rlabel metal1 6118 5678 6118 5678 0 net10
rlabel metal1 5382 1938 5382 1938 0 net11
rlabel metal1 1472 10030 1472 10030 0 net12
rlabel metal1 10626 11798 10626 11798 0 net13
rlabel metal1 9200 12206 9200 12206 0 net14
rlabel metal1 6716 12206 6716 12206 0 net15
rlabel metal1 7728 12206 7728 12206 0 net16
rlabel metal1 8418 11798 8418 11798 0 net17
rlabel metal1 10902 11798 10902 11798 0 net18
rlabel metal1 11178 11798 11178 11798 0 net19
rlabel metal1 2254 2618 2254 2618 0 net2
rlabel metal1 8050 12240 8050 12240 0 net20
rlabel metal1 9798 11764 9798 11764 0 net21
rlabel metal1 5750 11764 5750 11764 0 net22
rlabel metal1 9062 11526 9062 11526 0 net23
rlabel metal1 10350 11798 10350 11798 0 net24
rlabel metal1 5612 11730 5612 11730 0 net25
rlabel metal1 6026 11764 6026 11764 0 net26
rlabel metal1 6394 11764 6394 11764 0 net27
rlabel metal1 9338 11730 9338 11730 0 net28
rlabel metal1 12052 7310 12052 7310 0 net29
rlabel metal1 11960 2482 11960 2482 0 net3
rlabel metal1 8004 9486 8004 9486 0 net30
rlabel metal1 11960 4658 11960 4658 0 net4
rlabel metal2 12098 9792 12098 9792 0 net5
rlabel metal1 12052 11186 12052 11186 0 net6
rlabel metal1 11684 2550 11684 2550 0 net7
rlabel metal1 11960 5338 11960 5338 0 net8
rlabel metal1 6473 10778 6473 10778 0 net9
rlabel metal1 10074 7922 10074 7922 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal1 9706 7820 9706 7820 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal1 10028 7514 10028 7514 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal1 10396 6222 10396 6222 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal1 10166 6800 10166 6800 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 10074 6460 10074 6460 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal1 9844 4590 9844 4590 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal1 8372 5202 8372 5202 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal1 9890 5202 9890 5202 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 10948 10574 10948 10574 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal1 10350 8976 10350 8976 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal2 10166 8670 10166 8670 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal1 10856 5202 10856 5202 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal1 10258 5712 10258 5712 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal2 10166 4828 10166 4828 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal1 7452 9146 7452 9146 0 temp1.dac.vdac_single.en_pupd
rlabel metal1 12466 11050 12466 11050 0 temp1.dac_vout_notouch_
rlabel metal1 10718 11696 10718 11696 0 temp1.dcdel_capnode_notouch_
rlabel metal1 5157 11730 5157 11730 0 temp1.dcdel_out_n
rlabel metal1 6992 11186 6992 11186 0 temp1.i_precharge_n
rlabel metal1 5543 11526 5543 11526 0 temp1.o_tempdelay
rlabel metal1 4784 10438 4784 10438 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 13930 13898
<< end >>
